package constants is 

type state is (RI ,RL ,Pool_Cal_ReadImg , Pool_Read_Img , conv_calc_ReadImg_ReadBias  , conv_ReadImg_ReadFilter , conv_ReadImg  , CONV , SAVE , IMGSTAT , SHLEFT ,SHUP ,CHECKS  , WRITE_IMG_WIDTH , FINISH); 

end constants;