
-- 
-- Definition of  Main
-- 
--      Sat May 11 17:20:03 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity nBitRegister_1 is
   port (
      D : IN std_logic_vector (0 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      EN : IN std_logic ;
      Q : OUT std_logic_vector (0 DOWNTO 0)) ;
end nBitRegister_1 ;

architecture Data_flow of nBitRegister_1 is
   signal Q_0_EXMPLR, NOT_CLK, nx50: std_logic ;

begin
   Q(0) <= Q_0_EXMPLR ;
   reg_Q_0 : dffr port map ( Q=>Q_0_EXMPLR, QB=>OPEN, D=>nx50, CLK=>NOT_CLK, 
      R=>RST);
   ix51 : mux21_ni port map ( Y=>nx50, A0=>Q_0_EXMPLR, A1=>D(0), S0=>EN);
   ix63 : inv01 port map ( Y=>NOT_CLK, A=>CLK);
end Data_flow ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity triStateBuffer_13 is
   port (
      D : IN std_logic_vector (12 DOWNTO 0) ;
      EN : IN std_logic ;
      F : OUT std_logic_vector (12 DOWNTO 0)) ;
end triStateBuffer_13 ;

architecture triBuffer of triStateBuffer_13 is
   signal nx185, nx188, nx191, nx194, nx197, nx200, nx203, nx206, nx209, 
      nx212, nx215, nx218, nx221, nx228, nx230: std_logic ;

begin
   tri_F_0 : tri01 port map ( Y=>F(0), A=>nx185, E=>nx228);
   ix186 : inv01 port map ( Y=>nx185, A=>D(0));
   tri_F_1 : tri01 port map ( Y=>F(1), A=>nx188, E=>nx228);
   ix189 : inv01 port map ( Y=>nx188, A=>D(1));
   tri_F_2 : tri01 port map ( Y=>F(2), A=>nx191, E=>nx228);
   ix192 : inv01 port map ( Y=>nx191, A=>D(2));
   tri_F_3 : tri01 port map ( Y=>F(3), A=>nx194, E=>nx228);
   ix195 : inv01 port map ( Y=>nx194, A=>D(3));
   tri_F_4 : tri01 port map ( Y=>F(4), A=>nx197, E=>nx228);
   ix198 : inv01 port map ( Y=>nx197, A=>D(4));
   tri_F_5 : tri01 port map ( Y=>F(5), A=>nx200, E=>nx228);
   ix201 : inv01 port map ( Y=>nx200, A=>D(5));
   tri_F_6 : tri01 port map ( Y=>F(6), A=>nx203, E=>nx228);
   ix204 : inv01 port map ( Y=>nx203, A=>D(6));
   tri_F_7 : tri01 port map ( Y=>F(7), A=>nx206, E=>nx230);
   ix207 : inv01 port map ( Y=>nx206, A=>D(7));
   tri_F_8 : tri01 port map ( Y=>F(8), A=>nx209, E=>nx230);
   ix210 : inv01 port map ( Y=>nx209, A=>D(8));
   tri_F_9 : tri01 port map ( Y=>F(9), A=>nx212, E=>nx230);
   ix213 : inv01 port map ( Y=>nx212, A=>D(9));
   tri_F_10 : tri01 port map ( Y=>F(10), A=>nx215, E=>nx230);
   ix216 : inv01 port map ( Y=>nx215, A=>D(10));
   tri_F_11 : tri01 port map ( Y=>F(11), A=>nx218, E=>nx230);
   ix219 : inv01 port map ( Y=>nx218, A=>D(11));
   tri_F_12 : tri01 port map ( Y=>F(12), A=>nx221, E=>nx230);
   ix222 : inv01 port map ( Y=>nx221, A=>D(12));
   ix227 : buf02 port map ( Y=>nx228, A=>EN);
   ix229 : buf02 port map ( Y=>nx230, A=>EN);
end triBuffer ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity nBitRegister_13 is
   port (
      D : IN std_logic_vector (12 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      EN : IN std_logic ;
      Q : OUT std_logic_vector (12 DOWNTO 0)) ;
end nBitRegister_13 ;

architecture Data_flow of nBitRegister_13 is
   signal Q_12_EXMPLR, Q_11_EXMPLR, Q_10_EXMPLR, Q_9_EXMPLR, Q_8_EXMPLR, 
      Q_7_EXMPLR, Q_6_EXMPLR, Q_5_EXMPLR, Q_4_EXMPLR, Q_3_EXMPLR, Q_2_EXMPLR, 
      Q_1_EXMPLR, Q_0_EXMPLR, nx194, nx204, nx214, nx224, nx234, nx244, 
      nx254, nx264, nx274, nx284, nx294, nx304, nx314, nx370, nx372, nx378, 
      nx380, nx382, nx384: std_logic ;

begin
   Q(12) <= Q_12_EXMPLR ;
   Q(11) <= Q_11_EXMPLR ;
   Q(10) <= Q_10_EXMPLR ;
   Q(9) <= Q_9_EXMPLR ;
   Q(8) <= Q_8_EXMPLR ;
   Q(7) <= Q_7_EXMPLR ;
   Q(6) <= Q_6_EXMPLR ;
   Q(5) <= Q_5_EXMPLR ;
   Q(4) <= Q_4_EXMPLR ;
   Q(3) <= Q_3_EXMPLR ;
   Q(2) <= Q_2_EXMPLR ;
   Q(1) <= Q_1_EXMPLR ;
   Q(0) <= Q_0_EXMPLR ;
   reg_Q_0 : dffr port map ( Q=>Q_0_EXMPLR, QB=>OPEN, D=>nx194, CLK=>nx370, 
      R=>nx378);
   ix195 : mux21_ni port map ( Y=>nx194, A0=>Q_0_EXMPLR, A1=>D(0), S0=>nx382
   );
   reg_Q_1 : dffr port map ( Q=>Q_1_EXMPLR, QB=>OPEN, D=>nx204, CLK=>nx370, 
      R=>nx378);
   ix205 : mux21_ni port map ( Y=>nx204, A0=>Q_1_EXMPLR, A1=>D(1), S0=>nx382
   );
   reg_Q_2 : dffr port map ( Q=>Q_2_EXMPLR, QB=>OPEN, D=>nx214, CLK=>nx370, 
      R=>nx378);
   ix215 : mux21_ni port map ( Y=>nx214, A0=>Q_2_EXMPLR, A1=>D(2), S0=>nx382
   );
   reg_Q_3 : dffr port map ( Q=>Q_3_EXMPLR, QB=>OPEN, D=>nx224, CLK=>nx370, 
      R=>nx378);
   ix225 : mux21_ni port map ( Y=>nx224, A0=>Q_3_EXMPLR, A1=>D(3), S0=>nx382
   );
   reg_Q_4 : dffr port map ( Q=>Q_4_EXMPLR, QB=>OPEN, D=>nx234, CLK=>nx370, 
      R=>nx378);
   ix235 : mux21_ni port map ( Y=>nx234, A0=>Q_4_EXMPLR, A1=>D(4), S0=>nx382
   );
   reg_Q_5 : dffr port map ( Q=>Q_5_EXMPLR, QB=>OPEN, D=>nx244, CLK=>nx370, 
      R=>nx378);
   ix245 : mux21_ni port map ( Y=>nx244, A0=>Q_5_EXMPLR, A1=>D(5), S0=>nx382
   );
   reg_Q_6 : dffr port map ( Q=>Q_6_EXMPLR, QB=>OPEN, D=>nx254, CLK=>nx370, 
      R=>nx378);
   ix255 : mux21_ni port map ( Y=>nx254, A0=>Q_6_EXMPLR, A1=>D(6), S0=>nx382
   );
   reg_Q_7 : dffr port map ( Q=>Q_7_EXMPLR, QB=>OPEN, D=>nx264, CLK=>nx372, 
      R=>nx380);
   ix265 : mux21_ni port map ( Y=>nx264, A0=>Q_7_EXMPLR, A1=>D(7), S0=>nx384
   );
   reg_Q_8 : dffr port map ( Q=>Q_8_EXMPLR, QB=>OPEN, D=>nx274, CLK=>nx372, 
      R=>nx380);
   ix275 : mux21_ni port map ( Y=>nx274, A0=>Q_8_EXMPLR, A1=>D(8), S0=>nx384
   );
   reg_Q_9 : dffr port map ( Q=>Q_9_EXMPLR, QB=>OPEN, D=>nx284, CLK=>nx372, 
      R=>nx380);
   ix285 : mux21_ni port map ( Y=>nx284, A0=>Q_9_EXMPLR, A1=>D(9), S0=>nx384
   );
   reg_Q_10 : dffr port map ( Q=>Q_10_EXMPLR, QB=>OPEN, D=>nx294, CLK=>nx372, 
      R=>nx380);
   ix295 : mux21_ni port map ( Y=>nx294, A0=>Q_10_EXMPLR, A1=>D(10), S0=>
      nx384);
   reg_Q_11 : dffr port map ( Q=>Q_11_EXMPLR, QB=>OPEN, D=>nx304, CLK=>nx372, 
      R=>nx380);
   ix305 : mux21_ni port map ( Y=>nx304, A0=>Q_11_EXMPLR, A1=>D(11), S0=>
      nx384);
   reg_Q_12 : dffr port map ( Q=>Q_12_EXMPLR, QB=>OPEN, D=>nx314, CLK=>nx372, 
      R=>nx380);
   ix315 : mux21_ni port map ( Y=>nx314, A0=>Q_12_EXMPLR, A1=>D(12), S0=>
      nx384);
   ix369 : inv02 port map ( Y=>nx370, A=>CLK);
   ix371 : inv02 port map ( Y=>nx372, A=>CLK);
   ix377 : buf02 port map ( Y=>nx378, A=>RST);
   ix379 : buf02 port map ( Y=>nx380, A=>RST);
   ix381 : buf02 port map ( Y=>nx382, A=>EN);
   ix383 : buf02 port map ( Y=>nx384, A=>EN);
end Data_flow ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;
use ieee.numeric_std.all;
entity RAM_25 is
   port (
      reset : IN std_logic ;
      CLK : IN std_logic ;
      W : IN std_logic ;
      R : IN std_logic ;
      address : IN std_logic_vector (12 DOWNTO 0) ;
      dataIn : IN std_logic_vector (15 DOWNTO 0) ;
      dataOut : OUT std_logic_vector (399 DOWNTO 0) ;
      MFC : OUT std_logic ;
      counterOut : OUT std_logic_vector (3 DOWNTO 0)) ;
end RAM_25 ;

architecture archRAM of RAM_25 is
   type ram_type is array( 0 to 5000) of std_logic_vector(15 downto 0);
   signal ram: ram_type;
   signal mfc_m:std_logic;
   signal CLKEvent: std_logic;
   signal cReset,cEnable:std_logic;
   signal cOutput:std_logic_vector(3 downto 0);
   component Counter is
       generic(n: integer := 16);
       port(
           enable:in std_logic;
           reset:in std_logic;
           clk:in std_logic;
           load:in std_logic;
           output:out std_logic_vector(n-1 downto 0);
           input:in std_logic_vector(n-1 downto 0));
   end component;

begin
   -- enable the register when w or r signal comes
   cEnable <= '1' when (((W =  '1') or (R = '1')) and (mfc_m = '0'))
   else '0';
   counterOut <= cOutput;
   c1: Counter 
   generic map(4)
   port map(cEnable,cReset,CLK,'0',cOutput,"0001");

   -- MFC appears one clock after 8th clocks
   MFC <= mfc_m;
   --CLKEvent<= '1' when (CLK'event and CLK = '1')  else '0';
   
   mfc_m <= '1' when (cOutput = "0010" and(CLK'event and CLK = '1'))
   else '0' when   (CLK'event and CLK = '1');

   -- reset the counter when comes to 8 or a signal read or write
   cReset <= '1' when ((reset = '1') or (cOutput = "0011")) -- or (W'event and W = '1') or (R'event and R = '1') )
    else '0';

   -- memory retrieve 28 pixel of data after 8 bits
   process(cOutput)
  variable k,j,adds:integer;
   begin
       k := -16;
       j := -1;
       if  (cOutput = "0011" and W = '1')then
           ram(to_integer(unsigned(address))) <= dataIn;
       elsif  (cOutput = "0011" and R = '1')then
           loop1: for i in 0 to 25-1 loop
               k := k + 16;
               j := j + 16;
            adds := i + to_integer(unsigned(address));
               dataOut(j downto k) <= ram(adds);
         end loop;

--- we need to output z when we dont have data
       end if ;
   end process;
end archRAM ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity triStateBuffer_448 is
   port (
      D : IN std_logic_vector (447 DOWNTO 0) ;
      EN : IN std_logic ;
      F : OUT std_logic_vector (447 DOWNTO 0)) ;
end triStateBuffer_448 ;

architecture triBuffer of triStateBuffer_448 is
   signal nx4535, nx4538, nx4541, nx4544, nx4547, nx4550, nx4553, nx4556, 
      nx4559, nx4562, nx4565, nx4568, nx4571, nx4574, nx4577, nx4580, nx4583, 
      nx4586, nx4589, nx4592, nx4595, nx4598, nx4601, nx4604, nx4607, nx4610, 
      nx4613, nx4616, nx4619, nx4622, nx4625, nx4628, nx4631, nx4634, nx4637, 
      nx4640, nx4643, nx4646, nx4649, nx4652, nx4655, nx4658, nx4661, nx4664, 
      nx4667, nx4670, nx4673, nx4676, nx4679, nx4682, nx4685, nx4688, nx4691, 
      nx4694, nx4697, nx4700, nx4703, nx4706, nx4709, nx4712, nx4715, nx4718, 
      nx4721, nx4724, nx4727, nx4730, nx4733, nx4736, nx4739, nx4742, nx4745, 
      nx4748, nx4751, nx4754, nx4757, nx4760, nx4763, nx4766, nx4769, nx4772, 
      nx4775, nx4778, nx4781, nx4784, nx4787, nx4790, nx4793, nx4796, nx4799, 
      nx4802, nx4805, nx4808, nx4811, nx4814, nx4817, nx4820, nx4823, nx4826, 
      nx4829, nx4832, nx4835, nx4838, nx4841, nx4844, nx4847, nx4850, nx4853, 
      nx4856, nx4859, nx4862, nx4865, nx4868, nx4871, nx4874, nx4877, nx4880, 
      nx4883, nx4886, nx4889, nx4892, nx4895, nx4898, nx4901, nx4904, nx4907, 
      nx4910, nx4913, nx4916, nx4919, nx4922, nx4925, nx4928, nx4931, nx4934, 
      nx4937, nx4940, nx4943, nx4946, nx4949, nx4952, nx4955, nx4958, nx4961, 
      nx4964, nx4967, nx4970, nx4973, nx4976, nx4979, nx4982, nx4985, nx4988, 
      nx4991, nx4994, nx4997, nx5000, nx5003, nx5006, nx5009, nx5012, nx5015, 
      nx5018, nx5021, nx5024, nx5027, nx5030, nx5033, nx5036, nx5039, nx5042, 
      nx5045, nx5048, nx5051, nx5054, nx5057, nx5060, nx5063, nx5066, nx5069, 
      nx5072, nx5075, nx5078, nx5081, nx5084, nx5087, nx5090, nx5093, nx5096, 
      nx5099, nx5102, nx5105, nx5108, nx5111, nx5114, nx5117, nx5120, nx5123, 
      nx5126, nx5129, nx5132, nx5135, nx5138, nx5141, nx5144, nx5147, nx5150, 
      nx5153, nx5156, nx5159, nx5162, nx5165, nx5168, nx5171, nx5174, nx5177, 
      nx5180, nx5183, nx5186, nx5189, nx5192, nx5195, nx5198, nx5201, nx5204, 
      nx5207, nx5210, nx5213, nx5216, nx5219, nx5222, nx5225, nx5228, nx5231, 
      nx5234, nx5237, nx5240, nx5243, nx5246, nx5249, nx5252, nx5255, nx5258, 
      nx5261, nx5264, nx5267, nx5270, nx5273, nx5276, nx5279, nx5282, nx5285, 
      nx5288, nx5291, nx5294, nx5297, nx5300, nx5303, nx5306, nx5309, nx5312, 
      nx5315, nx5318, nx5321, nx5324, nx5327, nx5330, nx5333, nx5336, nx5339, 
      nx5342, nx5345, nx5348, nx5351, nx5354, nx5357, nx5360, nx5363, nx5366, 
      nx5369, nx5372, nx5375, nx5378, nx5381, nx5384, nx5387, nx5390, nx5393, 
      nx5396, nx5399, nx5402, nx5405, nx5408, nx5411, nx5414, nx5417, nx5420, 
      nx5423, nx5426, nx5429, nx5432, nx5435, nx5438, nx5441, nx5444, nx5447, 
      nx5450, nx5453, nx5456, nx5459, nx5462, nx5465, nx5468, nx5471, nx5474, 
      nx5477, nx5480, nx5483, nx5486, nx5489, nx5492, nx5495, nx5498, nx5501, 
      nx5504, nx5507, nx5510, nx5513, nx5516, nx5519, nx5522, nx5525, nx5528, 
      nx5531, nx5534, nx5537, nx5540, nx5543, nx5546, nx5549, nx5552, nx5555, 
      nx5558, nx5561, nx5564, nx5567, nx5570, nx5573, nx5576, nx5579, nx5582, 
      nx5585, nx5588, nx5591, nx5594, nx5597, nx5600, nx5603, nx5606, nx5609, 
      nx5612, nx5615, nx5618, nx5621, nx5624, nx5627, nx5630, nx5633, nx5636, 
      nx5639, nx5642, nx5645, nx5648, nx5651, nx5654, nx5657, nx5660, nx5663, 
      nx5666, nx5669, nx5672, nx5675, nx5678, nx5681, nx5684, nx5687, nx5690, 
      nx5693, nx5696, nx5699, nx5702, nx5705, nx5708, nx5711, nx5714, nx5717, 
      nx5720, nx5723, nx5726, nx5729, nx5732, nx5735, nx5738, nx5741, nx5744, 
      nx5747, nx5750, nx5753, nx5756, nx5759, nx5762, nx5765, nx5768, nx5771, 
      nx5774, nx5777, nx5780, nx5783, nx5786, nx5789, nx5792, nx5795, nx5798, 
      nx5801, nx5804, nx5807, nx5810, nx5813, nx5816, nx5819, nx5822, nx5825, 
      nx5828, nx5831, nx5834, nx5837, nx5840, nx5843, nx5846, nx5849, nx5852, 
      nx5855, nx5858, nx5861, nx5864, nx5867, nx5870, nx5873, nx5876, nx5883, 
      nx5885, nx5887, nx5889, nx5891, nx5893, nx5895, nx5897, nx5899, nx5901, 
      nx5903, nx5905, nx5907, nx5909, nx5911, nx5913, nx5915, nx5917, nx5919, 
      nx5921, nx5923, nx5925, nx5927, nx5929, nx5931, nx5933, nx5935, nx5937, 
      nx5939, nx5941, nx5943, nx5945, nx5947, nx5949, nx5951, nx5953, nx5955, 
      nx5957, nx5959, nx5961, nx5963, nx5965, nx5967, nx5969, nx5971, nx5973, 
      nx5975, nx5977, nx5979, nx5981, nx5983, nx5985, nx5987, nx5989, nx5991, 
      nx5993, nx5995, nx5997, nx5999, nx6001, nx6003, nx6005, nx6007, nx6009, 
      nx6011, nx6013, nx6015, nx6017, nx6019, nx6021, nx6023, nx6025, nx6027, 
      nx6029, nx6035, nx6037: std_logic ;

begin
   tri_F_0 : tri01 port map ( Y=>F(0), A=>nx4535, E=>nx5885);
   ix4536 : inv01 port map ( Y=>nx4535, A=>D(0));
   tri_F_1 : tri01 port map ( Y=>F(1), A=>nx4538, E=>nx5885);
   ix4539 : inv01 port map ( Y=>nx4538, A=>D(1));
   tri_F_2 : tri01 port map ( Y=>F(2), A=>nx4541, E=>nx5885);
   ix4542 : inv01 port map ( Y=>nx4541, A=>D(2));
   tri_F_3 : tri01 port map ( Y=>F(3), A=>nx4544, E=>nx5885);
   ix4545 : inv01 port map ( Y=>nx4544, A=>D(3));
   tri_F_4 : tri01 port map ( Y=>F(4), A=>nx4547, E=>nx5885);
   ix4548 : inv01 port map ( Y=>nx4547, A=>D(4));
   tri_F_5 : tri01 port map ( Y=>F(5), A=>nx4550, E=>nx5885);
   ix4551 : inv01 port map ( Y=>nx4550, A=>D(5));
   tri_F_6 : tri01 port map ( Y=>F(6), A=>nx4553, E=>nx5885);
   ix4554 : inv01 port map ( Y=>nx4553, A=>D(6));
   tri_F_7 : tri01 port map ( Y=>F(7), A=>nx4556, E=>nx5887);
   ix4557 : inv01 port map ( Y=>nx4556, A=>D(7));
   tri_F_8 : tri01 port map ( Y=>F(8), A=>nx4559, E=>nx5887);
   ix4560 : inv01 port map ( Y=>nx4559, A=>D(8));
   tri_F_9 : tri01 port map ( Y=>F(9), A=>nx4562, E=>nx5887);
   ix4563 : inv01 port map ( Y=>nx4562, A=>D(9));
   tri_F_10 : tri01 port map ( Y=>F(10), A=>nx4565, E=>nx5887);
   ix4566 : inv01 port map ( Y=>nx4565, A=>D(10));
   tri_F_11 : tri01 port map ( Y=>F(11), A=>nx4568, E=>nx5887);
   ix4569 : inv01 port map ( Y=>nx4568, A=>D(11));
   tri_F_12 : tri01 port map ( Y=>F(12), A=>nx4571, E=>nx5887);
   ix4572 : inv01 port map ( Y=>nx4571, A=>D(12));
   tri_F_13 : tri01 port map ( Y=>F(13), A=>nx4574, E=>nx5887);
   ix4575 : inv01 port map ( Y=>nx4574, A=>D(13));
   tri_F_14 : tri01 port map ( Y=>F(14), A=>nx4577, E=>nx5889);
   ix4578 : inv01 port map ( Y=>nx4577, A=>D(14));
   tri_F_15 : tri01 port map ( Y=>F(15), A=>nx4580, E=>nx5889);
   ix4581 : inv01 port map ( Y=>nx4580, A=>D(15));
   tri_F_16 : tri01 port map ( Y=>F(16), A=>nx4583, E=>nx5889);
   ix4584 : inv01 port map ( Y=>nx4583, A=>D(16));
   tri_F_17 : tri01 port map ( Y=>F(17), A=>nx4586, E=>nx5889);
   ix4587 : inv01 port map ( Y=>nx4586, A=>D(17));
   tri_F_18 : tri01 port map ( Y=>F(18), A=>nx4589, E=>nx5889);
   ix4590 : inv01 port map ( Y=>nx4589, A=>D(18));
   tri_F_19 : tri01 port map ( Y=>F(19), A=>nx4592, E=>nx5889);
   ix4593 : inv01 port map ( Y=>nx4592, A=>D(19));
   tri_F_20 : tri01 port map ( Y=>F(20), A=>nx4595, E=>nx5889);
   ix4596 : inv01 port map ( Y=>nx4595, A=>D(20));
   tri_F_21 : tri01 port map ( Y=>F(21), A=>nx4598, E=>nx5891);
   ix4599 : inv01 port map ( Y=>nx4598, A=>D(21));
   tri_F_22 : tri01 port map ( Y=>F(22), A=>nx4601, E=>nx5891);
   ix4602 : inv01 port map ( Y=>nx4601, A=>D(22));
   tri_F_23 : tri01 port map ( Y=>F(23), A=>nx4604, E=>nx5891);
   ix4605 : inv01 port map ( Y=>nx4604, A=>D(23));
   tri_F_24 : tri01 port map ( Y=>F(24), A=>nx4607, E=>nx5891);
   ix4608 : inv01 port map ( Y=>nx4607, A=>D(24));
   tri_F_25 : tri01 port map ( Y=>F(25), A=>nx4610, E=>nx5891);
   ix4611 : inv01 port map ( Y=>nx4610, A=>D(25));
   tri_F_26 : tri01 port map ( Y=>F(26), A=>nx4613, E=>nx5891);
   ix4614 : inv01 port map ( Y=>nx4613, A=>D(26));
   tri_F_27 : tri01 port map ( Y=>F(27), A=>nx4616, E=>nx5891);
   ix4617 : inv01 port map ( Y=>nx4616, A=>D(27));
   tri_F_28 : tri01 port map ( Y=>F(28), A=>nx4619, E=>nx5893);
   ix4620 : inv01 port map ( Y=>nx4619, A=>D(28));
   tri_F_29 : tri01 port map ( Y=>F(29), A=>nx4622, E=>nx5893);
   ix4623 : inv01 port map ( Y=>nx4622, A=>D(29));
   tri_F_30 : tri01 port map ( Y=>F(30), A=>nx4625, E=>nx5893);
   ix4626 : inv01 port map ( Y=>nx4625, A=>D(30));
   tri_F_31 : tri01 port map ( Y=>F(31), A=>nx4628, E=>nx5893);
   ix4629 : inv01 port map ( Y=>nx4628, A=>D(31));
   tri_F_32 : tri01 port map ( Y=>F(32), A=>nx4631, E=>nx5893);
   ix4632 : inv01 port map ( Y=>nx4631, A=>D(32));
   tri_F_33 : tri01 port map ( Y=>F(33), A=>nx4634, E=>nx5893);
   ix4635 : inv01 port map ( Y=>nx4634, A=>D(33));
   tri_F_34 : tri01 port map ( Y=>F(34), A=>nx4637, E=>nx5893);
   ix4638 : inv01 port map ( Y=>nx4637, A=>D(34));
   tri_F_35 : tri01 port map ( Y=>F(35), A=>nx4640, E=>nx5895);
   ix4641 : inv01 port map ( Y=>nx4640, A=>D(35));
   tri_F_36 : tri01 port map ( Y=>F(36), A=>nx4643, E=>nx5895);
   ix4644 : inv01 port map ( Y=>nx4643, A=>D(36));
   tri_F_37 : tri01 port map ( Y=>F(37), A=>nx4646, E=>nx5895);
   ix4647 : inv01 port map ( Y=>nx4646, A=>D(37));
   tri_F_38 : tri01 port map ( Y=>F(38), A=>nx4649, E=>nx5895);
   ix4650 : inv01 port map ( Y=>nx4649, A=>D(38));
   tri_F_39 : tri01 port map ( Y=>F(39), A=>nx4652, E=>nx5895);
   ix4653 : inv01 port map ( Y=>nx4652, A=>D(39));
   tri_F_40 : tri01 port map ( Y=>F(40), A=>nx4655, E=>nx5895);
   ix4656 : inv01 port map ( Y=>nx4655, A=>D(40));
   tri_F_41 : tri01 port map ( Y=>F(41), A=>nx4658, E=>nx5895);
   ix4659 : inv01 port map ( Y=>nx4658, A=>D(41));
   tri_F_42 : tri01 port map ( Y=>F(42), A=>nx4661, E=>nx5897);
   ix4662 : inv01 port map ( Y=>nx4661, A=>D(42));
   tri_F_43 : tri01 port map ( Y=>F(43), A=>nx4664, E=>nx5897);
   ix4665 : inv01 port map ( Y=>nx4664, A=>D(43));
   tri_F_44 : tri01 port map ( Y=>F(44), A=>nx4667, E=>nx5897);
   ix4668 : inv01 port map ( Y=>nx4667, A=>D(44));
   tri_F_45 : tri01 port map ( Y=>F(45), A=>nx4670, E=>nx5897);
   ix4671 : inv01 port map ( Y=>nx4670, A=>D(45));
   tri_F_46 : tri01 port map ( Y=>F(46), A=>nx4673, E=>nx5897);
   ix4674 : inv01 port map ( Y=>nx4673, A=>D(46));
   tri_F_47 : tri01 port map ( Y=>F(47), A=>nx4676, E=>nx5897);
   ix4677 : inv01 port map ( Y=>nx4676, A=>D(47));
   tri_F_48 : tri01 port map ( Y=>F(48), A=>nx4679, E=>nx5897);
   ix4680 : inv01 port map ( Y=>nx4679, A=>D(48));
   tri_F_49 : tri01 port map ( Y=>F(49), A=>nx4682, E=>nx5899);
   ix4683 : inv01 port map ( Y=>nx4682, A=>D(49));
   tri_F_50 : tri01 port map ( Y=>F(50), A=>nx4685, E=>nx5899);
   ix4686 : inv01 port map ( Y=>nx4685, A=>D(50));
   tri_F_51 : tri01 port map ( Y=>F(51), A=>nx4688, E=>nx5899);
   ix4689 : inv01 port map ( Y=>nx4688, A=>D(51));
   tri_F_52 : tri01 port map ( Y=>F(52), A=>nx4691, E=>nx5899);
   ix4692 : inv01 port map ( Y=>nx4691, A=>D(52));
   tri_F_53 : tri01 port map ( Y=>F(53), A=>nx4694, E=>nx5899);
   ix4695 : inv01 port map ( Y=>nx4694, A=>D(53));
   tri_F_54 : tri01 port map ( Y=>F(54), A=>nx4697, E=>nx5899);
   ix4698 : inv01 port map ( Y=>nx4697, A=>D(54));
   tri_F_55 : tri01 port map ( Y=>F(55), A=>nx4700, E=>nx5899);
   ix4701 : inv01 port map ( Y=>nx4700, A=>D(55));
   tri_F_56 : tri01 port map ( Y=>F(56), A=>nx4703, E=>nx5901);
   ix4704 : inv01 port map ( Y=>nx4703, A=>D(56));
   tri_F_57 : tri01 port map ( Y=>F(57), A=>nx4706, E=>nx5901);
   ix4707 : inv01 port map ( Y=>nx4706, A=>D(57));
   tri_F_58 : tri01 port map ( Y=>F(58), A=>nx4709, E=>nx5901);
   ix4710 : inv01 port map ( Y=>nx4709, A=>D(58));
   tri_F_59 : tri01 port map ( Y=>F(59), A=>nx4712, E=>nx5901);
   ix4713 : inv01 port map ( Y=>nx4712, A=>D(59));
   tri_F_60 : tri01 port map ( Y=>F(60), A=>nx4715, E=>nx5901);
   ix4716 : inv01 port map ( Y=>nx4715, A=>D(60));
   tri_F_61 : tri01 port map ( Y=>F(61), A=>nx4718, E=>nx5901);
   ix4719 : inv01 port map ( Y=>nx4718, A=>D(61));
   tri_F_62 : tri01 port map ( Y=>F(62), A=>nx4721, E=>nx5901);
   ix4722 : inv01 port map ( Y=>nx4721, A=>D(62));
   tri_F_63 : tri01 port map ( Y=>F(63), A=>nx4724, E=>nx5903);
   ix4725 : inv01 port map ( Y=>nx4724, A=>D(63));
   tri_F_64 : tri01 port map ( Y=>F(64), A=>nx4727, E=>nx5903);
   ix4728 : inv01 port map ( Y=>nx4727, A=>D(64));
   tri_F_65 : tri01 port map ( Y=>F(65), A=>nx4730, E=>nx5903);
   ix4731 : inv01 port map ( Y=>nx4730, A=>D(65));
   tri_F_66 : tri01 port map ( Y=>F(66), A=>nx4733, E=>nx5903);
   ix4734 : inv01 port map ( Y=>nx4733, A=>D(66));
   tri_F_67 : tri01 port map ( Y=>F(67), A=>nx4736, E=>nx5903);
   ix4737 : inv01 port map ( Y=>nx4736, A=>D(67));
   tri_F_68 : tri01 port map ( Y=>F(68), A=>nx4739, E=>nx5903);
   ix4740 : inv01 port map ( Y=>nx4739, A=>D(68));
   tri_F_69 : tri01 port map ( Y=>F(69), A=>nx4742, E=>nx5903);
   ix4743 : inv01 port map ( Y=>nx4742, A=>D(69));
   tri_F_70 : tri01 port map ( Y=>F(70), A=>nx4745, E=>nx5905);
   ix4746 : inv01 port map ( Y=>nx4745, A=>D(70));
   tri_F_71 : tri01 port map ( Y=>F(71), A=>nx4748, E=>nx5905);
   ix4749 : inv01 port map ( Y=>nx4748, A=>D(71));
   tri_F_72 : tri01 port map ( Y=>F(72), A=>nx4751, E=>nx5905);
   ix4752 : inv01 port map ( Y=>nx4751, A=>D(72));
   tri_F_73 : tri01 port map ( Y=>F(73), A=>nx4754, E=>nx5905);
   ix4755 : inv01 port map ( Y=>nx4754, A=>D(73));
   tri_F_74 : tri01 port map ( Y=>F(74), A=>nx4757, E=>nx5905);
   ix4758 : inv01 port map ( Y=>nx4757, A=>D(74));
   tri_F_75 : tri01 port map ( Y=>F(75), A=>nx4760, E=>nx5905);
   ix4761 : inv01 port map ( Y=>nx4760, A=>D(75));
   tri_F_76 : tri01 port map ( Y=>F(76), A=>nx4763, E=>nx5905);
   ix4764 : inv01 port map ( Y=>nx4763, A=>D(76));
   tri_F_77 : tri01 port map ( Y=>F(77), A=>nx4766, E=>nx5907);
   ix4767 : inv01 port map ( Y=>nx4766, A=>D(77));
   tri_F_78 : tri01 port map ( Y=>F(78), A=>nx4769, E=>nx5907);
   ix4770 : inv01 port map ( Y=>nx4769, A=>D(78));
   tri_F_79 : tri01 port map ( Y=>F(79), A=>nx4772, E=>nx5907);
   ix4773 : inv01 port map ( Y=>nx4772, A=>D(79));
   tri_F_80 : tri01 port map ( Y=>F(80), A=>nx4775, E=>nx5907);
   ix4776 : inv01 port map ( Y=>nx4775, A=>D(80));
   tri_F_81 : tri01 port map ( Y=>F(81), A=>nx4778, E=>nx5907);
   ix4779 : inv01 port map ( Y=>nx4778, A=>D(81));
   tri_F_82 : tri01 port map ( Y=>F(82), A=>nx4781, E=>nx5907);
   ix4782 : inv01 port map ( Y=>nx4781, A=>D(82));
   tri_F_83 : tri01 port map ( Y=>F(83), A=>nx4784, E=>nx5907);
   ix4785 : inv01 port map ( Y=>nx4784, A=>D(83));
   tri_F_84 : tri01 port map ( Y=>F(84), A=>nx4787, E=>nx5909);
   ix4788 : inv01 port map ( Y=>nx4787, A=>D(84));
   tri_F_85 : tri01 port map ( Y=>F(85), A=>nx4790, E=>nx5909);
   ix4791 : inv01 port map ( Y=>nx4790, A=>D(85));
   tri_F_86 : tri01 port map ( Y=>F(86), A=>nx4793, E=>nx5909);
   ix4794 : inv01 port map ( Y=>nx4793, A=>D(86));
   tri_F_87 : tri01 port map ( Y=>F(87), A=>nx4796, E=>nx5909);
   ix4797 : inv01 port map ( Y=>nx4796, A=>D(87));
   tri_F_88 : tri01 port map ( Y=>F(88), A=>nx4799, E=>nx5909);
   ix4800 : inv01 port map ( Y=>nx4799, A=>D(88));
   tri_F_89 : tri01 port map ( Y=>F(89), A=>nx4802, E=>nx5909);
   ix4803 : inv01 port map ( Y=>nx4802, A=>D(89));
   tri_F_90 : tri01 port map ( Y=>F(90), A=>nx4805, E=>nx5909);
   ix4806 : inv01 port map ( Y=>nx4805, A=>D(90));
   tri_F_91 : tri01 port map ( Y=>F(91), A=>nx4808, E=>nx5911);
   ix4809 : inv01 port map ( Y=>nx4808, A=>D(91));
   tri_F_92 : tri01 port map ( Y=>F(92), A=>nx4811, E=>nx5911);
   ix4812 : inv01 port map ( Y=>nx4811, A=>D(92));
   tri_F_93 : tri01 port map ( Y=>F(93), A=>nx4814, E=>nx5911);
   ix4815 : inv01 port map ( Y=>nx4814, A=>D(93));
   tri_F_94 : tri01 port map ( Y=>F(94), A=>nx4817, E=>nx5911);
   ix4818 : inv01 port map ( Y=>nx4817, A=>D(94));
   tri_F_95 : tri01 port map ( Y=>F(95), A=>nx4820, E=>nx5911);
   ix4821 : inv01 port map ( Y=>nx4820, A=>D(95));
   tri_F_96 : tri01 port map ( Y=>F(96), A=>nx4823, E=>nx5911);
   ix4824 : inv01 port map ( Y=>nx4823, A=>D(96));
   tri_F_97 : tri01 port map ( Y=>F(97), A=>nx4826, E=>nx5911);
   ix4827 : inv01 port map ( Y=>nx4826, A=>D(97));
   tri_F_98 : tri01 port map ( Y=>F(98), A=>nx4829, E=>nx5913);
   ix4830 : inv01 port map ( Y=>nx4829, A=>D(98));
   tri_F_99 : tri01 port map ( Y=>F(99), A=>nx4832, E=>nx5913);
   ix4833 : inv01 port map ( Y=>nx4832, A=>D(99));
   tri_F_100 : tri01 port map ( Y=>F(100), A=>nx4835, E=>nx5913);
   ix4836 : inv01 port map ( Y=>nx4835, A=>D(100));
   tri_F_101 : tri01 port map ( Y=>F(101), A=>nx4838, E=>nx5913);
   ix4839 : inv01 port map ( Y=>nx4838, A=>D(101));
   tri_F_102 : tri01 port map ( Y=>F(102), A=>nx4841, E=>nx5913);
   ix4842 : inv01 port map ( Y=>nx4841, A=>D(102));
   tri_F_103 : tri01 port map ( Y=>F(103), A=>nx4844, E=>nx5913);
   ix4845 : inv01 port map ( Y=>nx4844, A=>D(103));
   tri_F_104 : tri01 port map ( Y=>F(104), A=>nx4847, E=>nx5913);
   ix4848 : inv01 port map ( Y=>nx4847, A=>D(104));
   tri_F_105 : tri01 port map ( Y=>F(105), A=>nx4850, E=>nx5915);
   ix4851 : inv01 port map ( Y=>nx4850, A=>D(105));
   tri_F_106 : tri01 port map ( Y=>F(106), A=>nx4853, E=>nx5915);
   ix4854 : inv01 port map ( Y=>nx4853, A=>D(106));
   tri_F_107 : tri01 port map ( Y=>F(107), A=>nx4856, E=>nx5915);
   ix4857 : inv01 port map ( Y=>nx4856, A=>D(107));
   tri_F_108 : tri01 port map ( Y=>F(108), A=>nx4859, E=>nx5915);
   ix4860 : inv01 port map ( Y=>nx4859, A=>D(108));
   tri_F_109 : tri01 port map ( Y=>F(109), A=>nx4862, E=>nx5915);
   ix4863 : inv01 port map ( Y=>nx4862, A=>D(109));
   tri_F_110 : tri01 port map ( Y=>F(110), A=>nx4865, E=>nx5915);
   ix4866 : inv01 port map ( Y=>nx4865, A=>D(110));
   tri_F_111 : tri01 port map ( Y=>F(111), A=>nx4868, E=>nx5915);
   ix4869 : inv01 port map ( Y=>nx4868, A=>D(111));
   tri_F_112 : tri01 port map ( Y=>F(112), A=>nx4871, E=>nx5917);
   ix4872 : inv01 port map ( Y=>nx4871, A=>D(112));
   tri_F_113 : tri01 port map ( Y=>F(113), A=>nx4874, E=>nx5917);
   ix4875 : inv01 port map ( Y=>nx4874, A=>D(113));
   tri_F_114 : tri01 port map ( Y=>F(114), A=>nx4877, E=>nx5917);
   ix4878 : inv01 port map ( Y=>nx4877, A=>D(114));
   tri_F_115 : tri01 port map ( Y=>F(115), A=>nx4880, E=>nx5917);
   ix4881 : inv01 port map ( Y=>nx4880, A=>D(115));
   tri_F_116 : tri01 port map ( Y=>F(116), A=>nx4883, E=>nx5917);
   ix4884 : inv01 port map ( Y=>nx4883, A=>D(116));
   tri_F_117 : tri01 port map ( Y=>F(117), A=>nx4886, E=>nx5917);
   ix4887 : inv01 port map ( Y=>nx4886, A=>D(117));
   tri_F_118 : tri01 port map ( Y=>F(118), A=>nx4889, E=>nx5917);
   ix4890 : inv01 port map ( Y=>nx4889, A=>D(118));
   tri_F_119 : tri01 port map ( Y=>F(119), A=>nx4892, E=>nx5919);
   ix4893 : inv01 port map ( Y=>nx4892, A=>D(119));
   tri_F_120 : tri01 port map ( Y=>F(120), A=>nx4895, E=>nx5919);
   ix4896 : inv01 port map ( Y=>nx4895, A=>D(120));
   tri_F_121 : tri01 port map ( Y=>F(121), A=>nx4898, E=>nx5919);
   ix4899 : inv01 port map ( Y=>nx4898, A=>D(121));
   tri_F_122 : tri01 port map ( Y=>F(122), A=>nx4901, E=>nx5919);
   ix4902 : inv01 port map ( Y=>nx4901, A=>D(122));
   tri_F_123 : tri01 port map ( Y=>F(123), A=>nx4904, E=>nx5919);
   ix4905 : inv01 port map ( Y=>nx4904, A=>D(123));
   tri_F_124 : tri01 port map ( Y=>F(124), A=>nx4907, E=>nx5919);
   ix4908 : inv01 port map ( Y=>nx4907, A=>D(124));
   tri_F_125 : tri01 port map ( Y=>F(125), A=>nx4910, E=>nx5919);
   ix4911 : inv01 port map ( Y=>nx4910, A=>D(125));
   tri_F_126 : tri01 port map ( Y=>F(126), A=>nx4913, E=>nx5921);
   ix4914 : inv01 port map ( Y=>nx4913, A=>D(126));
   tri_F_127 : tri01 port map ( Y=>F(127), A=>nx4916, E=>nx5921);
   ix4917 : inv01 port map ( Y=>nx4916, A=>D(127));
   tri_F_128 : tri01 port map ( Y=>F(128), A=>nx4919, E=>nx5921);
   ix4920 : inv01 port map ( Y=>nx4919, A=>D(128));
   tri_F_129 : tri01 port map ( Y=>F(129), A=>nx4922, E=>nx5921);
   ix4923 : inv01 port map ( Y=>nx4922, A=>D(129));
   tri_F_130 : tri01 port map ( Y=>F(130), A=>nx4925, E=>nx5921);
   ix4926 : inv01 port map ( Y=>nx4925, A=>D(130));
   tri_F_131 : tri01 port map ( Y=>F(131), A=>nx4928, E=>nx5921);
   ix4929 : inv01 port map ( Y=>nx4928, A=>D(131));
   tri_F_132 : tri01 port map ( Y=>F(132), A=>nx4931, E=>nx5921);
   ix4932 : inv01 port map ( Y=>nx4931, A=>D(132));
   tri_F_133 : tri01 port map ( Y=>F(133), A=>nx4934, E=>nx5923);
   ix4935 : inv01 port map ( Y=>nx4934, A=>D(133));
   tri_F_134 : tri01 port map ( Y=>F(134), A=>nx4937, E=>nx5923);
   ix4938 : inv01 port map ( Y=>nx4937, A=>D(134));
   tri_F_135 : tri01 port map ( Y=>F(135), A=>nx4940, E=>nx5923);
   ix4941 : inv01 port map ( Y=>nx4940, A=>D(135));
   tri_F_136 : tri01 port map ( Y=>F(136), A=>nx4943, E=>nx5923);
   ix4944 : inv01 port map ( Y=>nx4943, A=>D(136));
   tri_F_137 : tri01 port map ( Y=>F(137), A=>nx4946, E=>nx5923);
   ix4947 : inv01 port map ( Y=>nx4946, A=>D(137));
   tri_F_138 : tri01 port map ( Y=>F(138), A=>nx4949, E=>nx5923);
   ix4950 : inv01 port map ( Y=>nx4949, A=>D(138));
   tri_F_139 : tri01 port map ( Y=>F(139), A=>nx4952, E=>nx5923);
   ix4953 : inv01 port map ( Y=>nx4952, A=>D(139));
   tri_F_140 : tri01 port map ( Y=>F(140), A=>nx4955, E=>nx5925);
   ix4956 : inv01 port map ( Y=>nx4955, A=>D(140));
   tri_F_141 : tri01 port map ( Y=>F(141), A=>nx4958, E=>nx5925);
   ix4959 : inv01 port map ( Y=>nx4958, A=>D(141));
   tri_F_142 : tri01 port map ( Y=>F(142), A=>nx4961, E=>nx5925);
   ix4962 : inv01 port map ( Y=>nx4961, A=>D(142));
   tri_F_143 : tri01 port map ( Y=>F(143), A=>nx4964, E=>nx5925);
   ix4965 : inv01 port map ( Y=>nx4964, A=>D(143));
   tri_F_144 : tri01 port map ( Y=>F(144), A=>nx4967, E=>nx5925);
   ix4968 : inv01 port map ( Y=>nx4967, A=>D(144));
   tri_F_145 : tri01 port map ( Y=>F(145), A=>nx4970, E=>nx5925);
   ix4971 : inv01 port map ( Y=>nx4970, A=>D(145));
   tri_F_146 : tri01 port map ( Y=>F(146), A=>nx4973, E=>nx5925);
   ix4974 : inv01 port map ( Y=>nx4973, A=>D(146));
   tri_F_147 : tri01 port map ( Y=>F(147), A=>nx4976, E=>nx5927);
   ix4977 : inv01 port map ( Y=>nx4976, A=>D(147));
   tri_F_148 : tri01 port map ( Y=>F(148), A=>nx4979, E=>nx5927);
   ix4980 : inv01 port map ( Y=>nx4979, A=>D(148));
   tri_F_149 : tri01 port map ( Y=>F(149), A=>nx4982, E=>nx5927);
   ix4983 : inv01 port map ( Y=>nx4982, A=>D(149));
   tri_F_150 : tri01 port map ( Y=>F(150), A=>nx4985, E=>nx5927);
   ix4986 : inv01 port map ( Y=>nx4985, A=>D(150));
   tri_F_151 : tri01 port map ( Y=>F(151), A=>nx4988, E=>nx5927);
   ix4989 : inv01 port map ( Y=>nx4988, A=>D(151));
   tri_F_152 : tri01 port map ( Y=>F(152), A=>nx4991, E=>nx5927);
   ix4992 : inv01 port map ( Y=>nx4991, A=>D(152));
   tri_F_153 : tri01 port map ( Y=>F(153), A=>nx4994, E=>nx5927);
   ix4995 : inv01 port map ( Y=>nx4994, A=>D(153));
   tri_F_154 : tri01 port map ( Y=>F(154), A=>nx4997, E=>nx5929);
   ix4998 : inv01 port map ( Y=>nx4997, A=>D(154));
   tri_F_155 : tri01 port map ( Y=>F(155), A=>nx5000, E=>nx5929);
   ix5001 : inv01 port map ( Y=>nx5000, A=>D(155));
   tri_F_156 : tri01 port map ( Y=>F(156), A=>nx5003, E=>nx5929);
   ix5004 : inv01 port map ( Y=>nx5003, A=>D(156));
   tri_F_157 : tri01 port map ( Y=>F(157), A=>nx5006, E=>nx5929);
   ix5007 : inv01 port map ( Y=>nx5006, A=>D(157));
   tri_F_158 : tri01 port map ( Y=>F(158), A=>nx5009, E=>nx5929);
   ix5010 : inv01 port map ( Y=>nx5009, A=>D(158));
   tri_F_159 : tri01 port map ( Y=>F(159), A=>nx5012, E=>nx5929);
   ix5013 : inv01 port map ( Y=>nx5012, A=>D(159));
   tri_F_160 : tri01 port map ( Y=>F(160), A=>nx5015, E=>nx5929);
   ix5016 : inv01 port map ( Y=>nx5015, A=>D(160));
   tri_F_161 : tri01 port map ( Y=>F(161), A=>nx5018, E=>nx5931);
   ix5019 : inv01 port map ( Y=>nx5018, A=>D(161));
   tri_F_162 : tri01 port map ( Y=>F(162), A=>nx5021, E=>nx5931);
   ix5022 : inv01 port map ( Y=>nx5021, A=>D(162));
   tri_F_163 : tri01 port map ( Y=>F(163), A=>nx5024, E=>nx5931);
   ix5025 : inv01 port map ( Y=>nx5024, A=>D(163));
   tri_F_164 : tri01 port map ( Y=>F(164), A=>nx5027, E=>nx5931);
   ix5028 : inv01 port map ( Y=>nx5027, A=>D(164));
   tri_F_165 : tri01 port map ( Y=>F(165), A=>nx5030, E=>nx5931);
   ix5031 : inv01 port map ( Y=>nx5030, A=>D(165));
   tri_F_166 : tri01 port map ( Y=>F(166), A=>nx5033, E=>nx5931);
   ix5034 : inv01 port map ( Y=>nx5033, A=>D(166));
   tri_F_167 : tri01 port map ( Y=>F(167), A=>nx5036, E=>nx5931);
   ix5037 : inv01 port map ( Y=>nx5036, A=>D(167));
   tri_F_168 : tri01 port map ( Y=>F(168), A=>nx5039, E=>nx5933);
   ix5040 : inv01 port map ( Y=>nx5039, A=>D(168));
   tri_F_169 : tri01 port map ( Y=>F(169), A=>nx5042, E=>nx5933);
   ix5043 : inv01 port map ( Y=>nx5042, A=>D(169));
   tri_F_170 : tri01 port map ( Y=>F(170), A=>nx5045, E=>nx5933);
   ix5046 : inv01 port map ( Y=>nx5045, A=>D(170));
   tri_F_171 : tri01 port map ( Y=>F(171), A=>nx5048, E=>nx5933);
   ix5049 : inv01 port map ( Y=>nx5048, A=>D(171));
   tri_F_172 : tri01 port map ( Y=>F(172), A=>nx5051, E=>nx5933);
   ix5052 : inv01 port map ( Y=>nx5051, A=>D(172));
   tri_F_173 : tri01 port map ( Y=>F(173), A=>nx5054, E=>nx5933);
   ix5055 : inv01 port map ( Y=>nx5054, A=>D(173));
   tri_F_174 : tri01 port map ( Y=>F(174), A=>nx5057, E=>nx5933);
   ix5058 : inv01 port map ( Y=>nx5057, A=>D(174));
   tri_F_175 : tri01 port map ( Y=>F(175), A=>nx5060, E=>nx5935);
   ix5061 : inv01 port map ( Y=>nx5060, A=>D(175));
   tri_F_176 : tri01 port map ( Y=>F(176), A=>nx5063, E=>nx5935);
   ix5064 : inv01 port map ( Y=>nx5063, A=>D(176));
   tri_F_177 : tri01 port map ( Y=>F(177), A=>nx5066, E=>nx5935);
   ix5067 : inv01 port map ( Y=>nx5066, A=>D(177));
   tri_F_178 : tri01 port map ( Y=>F(178), A=>nx5069, E=>nx5935);
   ix5070 : inv01 port map ( Y=>nx5069, A=>D(178));
   tri_F_179 : tri01 port map ( Y=>F(179), A=>nx5072, E=>nx5935);
   ix5073 : inv01 port map ( Y=>nx5072, A=>D(179));
   tri_F_180 : tri01 port map ( Y=>F(180), A=>nx5075, E=>nx5935);
   ix5076 : inv01 port map ( Y=>nx5075, A=>D(180));
   tri_F_181 : tri01 port map ( Y=>F(181), A=>nx5078, E=>nx5935);
   ix5079 : inv01 port map ( Y=>nx5078, A=>D(181));
   tri_F_182 : tri01 port map ( Y=>F(182), A=>nx5081, E=>nx5937);
   ix5082 : inv01 port map ( Y=>nx5081, A=>D(182));
   tri_F_183 : tri01 port map ( Y=>F(183), A=>nx5084, E=>nx5937);
   ix5085 : inv01 port map ( Y=>nx5084, A=>D(183));
   tri_F_184 : tri01 port map ( Y=>F(184), A=>nx5087, E=>nx5937);
   ix5088 : inv01 port map ( Y=>nx5087, A=>D(184));
   tri_F_185 : tri01 port map ( Y=>F(185), A=>nx5090, E=>nx5937);
   ix5091 : inv01 port map ( Y=>nx5090, A=>D(185));
   tri_F_186 : tri01 port map ( Y=>F(186), A=>nx5093, E=>nx5937);
   ix5094 : inv01 port map ( Y=>nx5093, A=>D(186));
   tri_F_187 : tri01 port map ( Y=>F(187), A=>nx5096, E=>nx5937);
   ix5097 : inv01 port map ( Y=>nx5096, A=>D(187));
   tri_F_188 : tri01 port map ( Y=>F(188), A=>nx5099, E=>nx5937);
   ix5100 : inv01 port map ( Y=>nx5099, A=>D(188));
   tri_F_189 : tri01 port map ( Y=>F(189), A=>nx5102, E=>nx5939);
   ix5103 : inv01 port map ( Y=>nx5102, A=>D(189));
   tri_F_190 : tri01 port map ( Y=>F(190), A=>nx5105, E=>nx5939);
   ix5106 : inv01 port map ( Y=>nx5105, A=>D(190));
   tri_F_191 : tri01 port map ( Y=>F(191), A=>nx5108, E=>nx5939);
   ix5109 : inv01 port map ( Y=>nx5108, A=>D(191));
   tri_F_192 : tri01 port map ( Y=>F(192), A=>nx5111, E=>nx5939);
   ix5112 : inv01 port map ( Y=>nx5111, A=>D(192));
   tri_F_193 : tri01 port map ( Y=>F(193), A=>nx5114, E=>nx5939);
   ix5115 : inv01 port map ( Y=>nx5114, A=>D(193));
   tri_F_194 : tri01 port map ( Y=>F(194), A=>nx5117, E=>nx5939);
   ix5118 : inv01 port map ( Y=>nx5117, A=>D(194));
   tri_F_195 : tri01 port map ( Y=>F(195), A=>nx5120, E=>nx5939);
   ix5121 : inv01 port map ( Y=>nx5120, A=>D(195));
   tri_F_196 : tri01 port map ( Y=>F(196), A=>nx5123, E=>nx5941);
   ix5124 : inv01 port map ( Y=>nx5123, A=>D(196));
   tri_F_197 : tri01 port map ( Y=>F(197), A=>nx5126, E=>nx5941);
   ix5127 : inv01 port map ( Y=>nx5126, A=>D(197));
   tri_F_198 : tri01 port map ( Y=>F(198), A=>nx5129, E=>nx5941);
   ix5130 : inv01 port map ( Y=>nx5129, A=>D(198));
   tri_F_199 : tri01 port map ( Y=>F(199), A=>nx5132, E=>nx5941);
   ix5133 : inv01 port map ( Y=>nx5132, A=>D(199));
   tri_F_200 : tri01 port map ( Y=>F(200), A=>nx5135, E=>nx5941);
   ix5136 : inv01 port map ( Y=>nx5135, A=>D(200));
   tri_F_201 : tri01 port map ( Y=>F(201), A=>nx5138, E=>nx5941);
   ix5139 : inv01 port map ( Y=>nx5138, A=>D(201));
   tri_F_202 : tri01 port map ( Y=>F(202), A=>nx5141, E=>nx5941);
   ix5142 : inv01 port map ( Y=>nx5141, A=>D(202));
   tri_F_203 : tri01 port map ( Y=>F(203), A=>nx5144, E=>nx5943);
   ix5145 : inv01 port map ( Y=>nx5144, A=>D(203));
   tri_F_204 : tri01 port map ( Y=>F(204), A=>nx5147, E=>nx5943);
   ix5148 : inv01 port map ( Y=>nx5147, A=>D(204));
   tri_F_205 : tri01 port map ( Y=>F(205), A=>nx5150, E=>nx5943);
   ix5151 : inv01 port map ( Y=>nx5150, A=>D(205));
   tri_F_206 : tri01 port map ( Y=>F(206), A=>nx5153, E=>nx5943);
   ix5154 : inv01 port map ( Y=>nx5153, A=>D(206));
   tri_F_207 : tri01 port map ( Y=>F(207), A=>nx5156, E=>nx5943);
   ix5157 : inv01 port map ( Y=>nx5156, A=>D(207));
   tri_F_208 : tri01 port map ( Y=>F(208), A=>nx5159, E=>nx5943);
   ix5160 : inv01 port map ( Y=>nx5159, A=>D(208));
   tri_F_209 : tri01 port map ( Y=>F(209), A=>nx5162, E=>nx5943);
   ix5163 : inv01 port map ( Y=>nx5162, A=>D(209));
   tri_F_210 : tri01 port map ( Y=>F(210), A=>nx5165, E=>nx5945);
   ix5166 : inv01 port map ( Y=>nx5165, A=>D(210));
   tri_F_211 : tri01 port map ( Y=>F(211), A=>nx5168, E=>nx5945);
   ix5169 : inv01 port map ( Y=>nx5168, A=>D(211));
   tri_F_212 : tri01 port map ( Y=>F(212), A=>nx5171, E=>nx5945);
   ix5172 : inv01 port map ( Y=>nx5171, A=>D(212));
   tri_F_213 : tri01 port map ( Y=>F(213), A=>nx5174, E=>nx5945);
   ix5175 : inv01 port map ( Y=>nx5174, A=>D(213));
   tri_F_214 : tri01 port map ( Y=>F(214), A=>nx5177, E=>nx5945);
   ix5178 : inv01 port map ( Y=>nx5177, A=>D(214));
   tri_F_215 : tri01 port map ( Y=>F(215), A=>nx5180, E=>nx5945);
   ix5181 : inv01 port map ( Y=>nx5180, A=>D(215));
   tri_F_216 : tri01 port map ( Y=>F(216), A=>nx5183, E=>nx5945);
   ix5184 : inv01 port map ( Y=>nx5183, A=>D(216));
   tri_F_217 : tri01 port map ( Y=>F(217), A=>nx5186, E=>nx5947);
   ix5187 : inv01 port map ( Y=>nx5186, A=>D(217));
   tri_F_218 : tri01 port map ( Y=>F(218), A=>nx5189, E=>nx5947);
   ix5190 : inv01 port map ( Y=>nx5189, A=>D(218));
   tri_F_219 : tri01 port map ( Y=>F(219), A=>nx5192, E=>nx5947);
   ix5193 : inv01 port map ( Y=>nx5192, A=>D(219));
   tri_F_220 : tri01 port map ( Y=>F(220), A=>nx5195, E=>nx5947);
   ix5196 : inv01 port map ( Y=>nx5195, A=>D(220));
   tri_F_221 : tri01 port map ( Y=>F(221), A=>nx5198, E=>nx5947);
   ix5199 : inv01 port map ( Y=>nx5198, A=>D(221));
   tri_F_222 : tri01 port map ( Y=>F(222), A=>nx5201, E=>nx5947);
   ix5202 : inv01 port map ( Y=>nx5201, A=>D(222));
   tri_F_223 : tri01 port map ( Y=>F(223), A=>nx5204, E=>nx5947);
   ix5205 : inv01 port map ( Y=>nx5204, A=>D(223));
   tri_F_224 : tri01 port map ( Y=>F(224), A=>nx5207, E=>nx5949);
   ix5208 : inv01 port map ( Y=>nx5207, A=>D(224));
   tri_F_225 : tri01 port map ( Y=>F(225), A=>nx5210, E=>nx5949);
   ix5211 : inv01 port map ( Y=>nx5210, A=>D(225));
   tri_F_226 : tri01 port map ( Y=>F(226), A=>nx5213, E=>nx5949);
   ix5214 : inv01 port map ( Y=>nx5213, A=>D(226));
   tri_F_227 : tri01 port map ( Y=>F(227), A=>nx5216, E=>nx5949);
   ix5217 : inv01 port map ( Y=>nx5216, A=>D(227));
   tri_F_228 : tri01 port map ( Y=>F(228), A=>nx5219, E=>nx5949);
   ix5220 : inv01 port map ( Y=>nx5219, A=>D(228));
   tri_F_229 : tri01 port map ( Y=>F(229), A=>nx5222, E=>nx5949);
   ix5223 : inv01 port map ( Y=>nx5222, A=>D(229));
   tri_F_230 : tri01 port map ( Y=>F(230), A=>nx5225, E=>nx5949);
   ix5226 : inv01 port map ( Y=>nx5225, A=>D(230));
   tri_F_231 : tri01 port map ( Y=>F(231), A=>nx5228, E=>nx5951);
   ix5229 : inv01 port map ( Y=>nx5228, A=>D(231));
   tri_F_232 : tri01 port map ( Y=>F(232), A=>nx5231, E=>nx5951);
   ix5232 : inv01 port map ( Y=>nx5231, A=>D(232));
   tri_F_233 : tri01 port map ( Y=>F(233), A=>nx5234, E=>nx5951);
   ix5235 : inv01 port map ( Y=>nx5234, A=>D(233));
   tri_F_234 : tri01 port map ( Y=>F(234), A=>nx5237, E=>nx5951);
   ix5238 : inv01 port map ( Y=>nx5237, A=>D(234));
   tri_F_235 : tri01 port map ( Y=>F(235), A=>nx5240, E=>nx5951);
   ix5241 : inv01 port map ( Y=>nx5240, A=>D(235));
   tri_F_236 : tri01 port map ( Y=>F(236), A=>nx5243, E=>nx5951);
   ix5244 : inv01 port map ( Y=>nx5243, A=>D(236));
   tri_F_237 : tri01 port map ( Y=>F(237), A=>nx5246, E=>nx5951);
   ix5247 : inv01 port map ( Y=>nx5246, A=>D(237));
   tri_F_238 : tri01 port map ( Y=>F(238), A=>nx5249, E=>nx5953);
   ix5250 : inv01 port map ( Y=>nx5249, A=>D(238));
   tri_F_239 : tri01 port map ( Y=>F(239), A=>nx5252, E=>nx5953);
   ix5253 : inv01 port map ( Y=>nx5252, A=>D(239));
   tri_F_240 : tri01 port map ( Y=>F(240), A=>nx5255, E=>nx5953);
   ix5256 : inv01 port map ( Y=>nx5255, A=>D(240));
   tri_F_241 : tri01 port map ( Y=>F(241), A=>nx5258, E=>nx5953);
   ix5259 : inv01 port map ( Y=>nx5258, A=>D(241));
   tri_F_242 : tri01 port map ( Y=>F(242), A=>nx5261, E=>nx5953);
   ix5262 : inv01 port map ( Y=>nx5261, A=>D(242));
   tri_F_243 : tri01 port map ( Y=>F(243), A=>nx5264, E=>nx5953);
   ix5265 : inv01 port map ( Y=>nx5264, A=>D(243));
   tri_F_244 : tri01 port map ( Y=>F(244), A=>nx5267, E=>nx5953);
   ix5268 : inv01 port map ( Y=>nx5267, A=>D(244));
   tri_F_245 : tri01 port map ( Y=>F(245), A=>nx5270, E=>nx5955);
   ix5271 : inv01 port map ( Y=>nx5270, A=>D(245));
   tri_F_246 : tri01 port map ( Y=>F(246), A=>nx5273, E=>nx5955);
   ix5274 : inv01 port map ( Y=>nx5273, A=>D(246));
   tri_F_247 : tri01 port map ( Y=>F(247), A=>nx5276, E=>nx5955);
   ix5277 : inv01 port map ( Y=>nx5276, A=>D(247));
   tri_F_248 : tri01 port map ( Y=>F(248), A=>nx5279, E=>nx5955);
   ix5280 : inv01 port map ( Y=>nx5279, A=>D(248));
   tri_F_249 : tri01 port map ( Y=>F(249), A=>nx5282, E=>nx5955);
   ix5283 : inv01 port map ( Y=>nx5282, A=>D(249));
   tri_F_250 : tri01 port map ( Y=>F(250), A=>nx5285, E=>nx5955);
   ix5286 : inv01 port map ( Y=>nx5285, A=>D(250));
   tri_F_251 : tri01 port map ( Y=>F(251), A=>nx5288, E=>nx5955);
   ix5289 : inv01 port map ( Y=>nx5288, A=>D(251));
   tri_F_252 : tri01 port map ( Y=>F(252), A=>nx5291, E=>nx5957);
   ix5292 : inv01 port map ( Y=>nx5291, A=>D(252));
   tri_F_253 : tri01 port map ( Y=>F(253), A=>nx5294, E=>nx5957);
   ix5295 : inv01 port map ( Y=>nx5294, A=>D(253));
   tri_F_254 : tri01 port map ( Y=>F(254), A=>nx5297, E=>nx5957);
   ix5298 : inv01 port map ( Y=>nx5297, A=>D(254));
   tri_F_255 : tri01 port map ( Y=>F(255), A=>nx5300, E=>nx5957);
   ix5301 : inv01 port map ( Y=>nx5300, A=>D(255));
   tri_F_256 : tri01 port map ( Y=>F(256), A=>nx5303, E=>nx5957);
   ix5304 : inv01 port map ( Y=>nx5303, A=>D(256));
   tri_F_257 : tri01 port map ( Y=>F(257), A=>nx5306, E=>nx5957);
   ix5307 : inv01 port map ( Y=>nx5306, A=>D(257));
   tri_F_258 : tri01 port map ( Y=>F(258), A=>nx5309, E=>nx5957);
   ix5310 : inv01 port map ( Y=>nx5309, A=>D(258));
   tri_F_259 : tri01 port map ( Y=>F(259), A=>nx5312, E=>nx5959);
   ix5313 : inv01 port map ( Y=>nx5312, A=>D(259));
   tri_F_260 : tri01 port map ( Y=>F(260), A=>nx5315, E=>nx5959);
   ix5316 : inv01 port map ( Y=>nx5315, A=>D(260));
   tri_F_261 : tri01 port map ( Y=>F(261), A=>nx5318, E=>nx5959);
   ix5319 : inv01 port map ( Y=>nx5318, A=>D(261));
   tri_F_262 : tri01 port map ( Y=>F(262), A=>nx5321, E=>nx5959);
   ix5322 : inv01 port map ( Y=>nx5321, A=>D(262));
   tri_F_263 : tri01 port map ( Y=>F(263), A=>nx5324, E=>nx5959);
   ix5325 : inv01 port map ( Y=>nx5324, A=>D(263));
   tri_F_264 : tri01 port map ( Y=>F(264), A=>nx5327, E=>nx5959);
   ix5328 : inv01 port map ( Y=>nx5327, A=>D(264));
   tri_F_265 : tri01 port map ( Y=>F(265), A=>nx5330, E=>nx5959);
   ix5331 : inv01 port map ( Y=>nx5330, A=>D(265));
   tri_F_266 : tri01 port map ( Y=>F(266), A=>nx5333, E=>nx5961);
   ix5334 : inv01 port map ( Y=>nx5333, A=>D(266));
   tri_F_267 : tri01 port map ( Y=>F(267), A=>nx5336, E=>nx5961);
   ix5337 : inv01 port map ( Y=>nx5336, A=>D(267));
   tri_F_268 : tri01 port map ( Y=>F(268), A=>nx5339, E=>nx5961);
   ix5340 : inv01 port map ( Y=>nx5339, A=>D(268));
   tri_F_269 : tri01 port map ( Y=>F(269), A=>nx5342, E=>nx5961);
   ix5343 : inv01 port map ( Y=>nx5342, A=>D(269));
   tri_F_270 : tri01 port map ( Y=>F(270), A=>nx5345, E=>nx5961);
   ix5346 : inv01 port map ( Y=>nx5345, A=>D(270));
   tri_F_271 : tri01 port map ( Y=>F(271), A=>nx5348, E=>nx5961);
   ix5349 : inv01 port map ( Y=>nx5348, A=>D(271));
   tri_F_272 : tri01 port map ( Y=>F(272), A=>nx5351, E=>nx5961);
   ix5352 : inv01 port map ( Y=>nx5351, A=>D(272));
   tri_F_273 : tri01 port map ( Y=>F(273), A=>nx5354, E=>nx5963);
   ix5355 : inv01 port map ( Y=>nx5354, A=>D(273));
   tri_F_274 : tri01 port map ( Y=>F(274), A=>nx5357, E=>nx5963);
   ix5358 : inv01 port map ( Y=>nx5357, A=>D(274));
   tri_F_275 : tri01 port map ( Y=>F(275), A=>nx5360, E=>nx5963);
   ix5361 : inv01 port map ( Y=>nx5360, A=>D(275));
   tri_F_276 : tri01 port map ( Y=>F(276), A=>nx5363, E=>nx5963);
   ix5364 : inv01 port map ( Y=>nx5363, A=>D(276));
   tri_F_277 : tri01 port map ( Y=>F(277), A=>nx5366, E=>nx5963);
   ix5367 : inv01 port map ( Y=>nx5366, A=>D(277));
   tri_F_278 : tri01 port map ( Y=>F(278), A=>nx5369, E=>nx5963);
   ix5370 : inv01 port map ( Y=>nx5369, A=>D(278));
   tri_F_279 : tri01 port map ( Y=>F(279), A=>nx5372, E=>nx5963);
   ix5373 : inv01 port map ( Y=>nx5372, A=>D(279));
   tri_F_280 : tri01 port map ( Y=>F(280), A=>nx5375, E=>nx5965);
   ix5376 : inv01 port map ( Y=>nx5375, A=>D(280));
   tri_F_281 : tri01 port map ( Y=>F(281), A=>nx5378, E=>nx5965);
   ix5379 : inv01 port map ( Y=>nx5378, A=>D(281));
   tri_F_282 : tri01 port map ( Y=>F(282), A=>nx5381, E=>nx5965);
   ix5382 : inv01 port map ( Y=>nx5381, A=>D(282));
   tri_F_283 : tri01 port map ( Y=>F(283), A=>nx5384, E=>nx5965);
   ix5385 : inv01 port map ( Y=>nx5384, A=>D(283));
   tri_F_284 : tri01 port map ( Y=>F(284), A=>nx5387, E=>nx5965);
   ix5388 : inv01 port map ( Y=>nx5387, A=>D(284));
   tri_F_285 : tri01 port map ( Y=>F(285), A=>nx5390, E=>nx5965);
   ix5391 : inv01 port map ( Y=>nx5390, A=>D(285));
   tri_F_286 : tri01 port map ( Y=>F(286), A=>nx5393, E=>nx5965);
   ix5394 : inv01 port map ( Y=>nx5393, A=>D(286));
   tri_F_287 : tri01 port map ( Y=>F(287), A=>nx5396, E=>nx5967);
   ix5397 : inv01 port map ( Y=>nx5396, A=>D(287));
   tri_F_288 : tri01 port map ( Y=>F(288), A=>nx5399, E=>nx5967);
   ix5400 : inv01 port map ( Y=>nx5399, A=>D(288));
   tri_F_289 : tri01 port map ( Y=>F(289), A=>nx5402, E=>nx5967);
   ix5403 : inv01 port map ( Y=>nx5402, A=>D(289));
   tri_F_290 : tri01 port map ( Y=>F(290), A=>nx5405, E=>nx5967);
   ix5406 : inv01 port map ( Y=>nx5405, A=>D(290));
   tri_F_291 : tri01 port map ( Y=>F(291), A=>nx5408, E=>nx5967);
   ix5409 : inv01 port map ( Y=>nx5408, A=>D(291));
   tri_F_292 : tri01 port map ( Y=>F(292), A=>nx5411, E=>nx5967);
   ix5412 : inv01 port map ( Y=>nx5411, A=>D(292));
   tri_F_293 : tri01 port map ( Y=>F(293), A=>nx5414, E=>nx5967);
   ix5415 : inv01 port map ( Y=>nx5414, A=>D(293));
   tri_F_294 : tri01 port map ( Y=>F(294), A=>nx5417, E=>nx5969);
   ix5418 : inv01 port map ( Y=>nx5417, A=>D(294));
   tri_F_295 : tri01 port map ( Y=>F(295), A=>nx5420, E=>nx5969);
   ix5421 : inv01 port map ( Y=>nx5420, A=>D(295));
   tri_F_296 : tri01 port map ( Y=>F(296), A=>nx5423, E=>nx5969);
   ix5424 : inv01 port map ( Y=>nx5423, A=>D(296));
   tri_F_297 : tri01 port map ( Y=>F(297), A=>nx5426, E=>nx5969);
   ix5427 : inv01 port map ( Y=>nx5426, A=>D(297));
   tri_F_298 : tri01 port map ( Y=>F(298), A=>nx5429, E=>nx5969);
   ix5430 : inv01 port map ( Y=>nx5429, A=>D(298));
   tri_F_299 : tri01 port map ( Y=>F(299), A=>nx5432, E=>nx5969);
   ix5433 : inv01 port map ( Y=>nx5432, A=>D(299));
   tri_F_300 : tri01 port map ( Y=>F(300), A=>nx5435, E=>nx5969);
   ix5436 : inv01 port map ( Y=>nx5435, A=>D(300));
   tri_F_301 : tri01 port map ( Y=>F(301), A=>nx5438, E=>nx5971);
   ix5439 : inv01 port map ( Y=>nx5438, A=>D(301));
   tri_F_302 : tri01 port map ( Y=>F(302), A=>nx5441, E=>nx5971);
   ix5442 : inv01 port map ( Y=>nx5441, A=>D(302));
   tri_F_303 : tri01 port map ( Y=>F(303), A=>nx5444, E=>nx5971);
   ix5445 : inv01 port map ( Y=>nx5444, A=>D(303));
   tri_F_304 : tri01 port map ( Y=>F(304), A=>nx5447, E=>nx5971);
   ix5448 : inv01 port map ( Y=>nx5447, A=>D(304));
   tri_F_305 : tri01 port map ( Y=>F(305), A=>nx5450, E=>nx5971);
   ix5451 : inv01 port map ( Y=>nx5450, A=>D(305));
   tri_F_306 : tri01 port map ( Y=>F(306), A=>nx5453, E=>nx5971);
   ix5454 : inv01 port map ( Y=>nx5453, A=>D(306));
   tri_F_307 : tri01 port map ( Y=>F(307), A=>nx5456, E=>nx5971);
   ix5457 : inv01 port map ( Y=>nx5456, A=>D(307));
   tri_F_308 : tri01 port map ( Y=>F(308), A=>nx5459, E=>nx5973);
   ix5460 : inv01 port map ( Y=>nx5459, A=>D(308));
   tri_F_309 : tri01 port map ( Y=>F(309), A=>nx5462, E=>nx5973);
   ix5463 : inv01 port map ( Y=>nx5462, A=>D(309));
   tri_F_310 : tri01 port map ( Y=>F(310), A=>nx5465, E=>nx5973);
   ix5466 : inv01 port map ( Y=>nx5465, A=>D(310));
   tri_F_311 : tri01 port map ( Y=>F(311), A=>nx5468, E=>nx5973);
   ix5469 : inv01 port map ( Y=>nx5468, A=>D(311));
   tri_F_312 : tri01 port map ( Y=>F(312), A=>nx5471, E=>nx5973);
   ix5472 : inv01 port map ( Y=>nx5471, A=>D(312));
   tri_F_313 : tri01 port map ( Y=>F(313), A=>nx5474, E=>nx5973);
   ix5475 : inv01 port map ( Y=>nx5474, A=>D(313));
   tri_F_314 : tri01 port map ( Y=>F(314), A=>nx5477, E=>nx5973);
   ix5478 : inv01 port map ( Y=>nx5477, A=>D(314));
   tri_F_315 : tri01 port map ( Y=>F(315), A=>nx5480, E=>nx5975);
   ix5481 : inv01 port map ( Y=>nx5480, A=>D(315));
   tri_F_316 : tri01 port map ( Y=>F(316), A=>nx5483, E=>nx5975);
   ix5484 : inv01 port map ( Y=>nx5483, A=>D(316));
   tri_F_317 : tri01 port map ( Y=>F(317), A=>nx5486, E=>nx5975);
   ix5487 : inv01 port map ( Y=>nx5486, A=>D(317));
   tri_F_318 : tri01 port map ( Y=>F(318), A=>nx5489, E=>nx5975);
   ix5490 : inv01 port map ( Y=>nx5489, A=>D(318));
   tri_F_319 : tri01 port map ( Y=>F(319), A=>nx5492, E=>nx5975);
   ix5493 : inv01 port map ( Y=>nx5492, A=>D(319));
   tri_F_320 : tri01 port map ( Y=>F(320), A=>nx5495, E=>nx5975);
   ix5496 : inv01 port map ( Y=>nx5495, A=>D(320));
   tri_F_321 : tri01 port map ( Y=>F(321), A=>nx5498, E=>nx5975);
   ix5499 : inv01 port map ( Y=>nx5498, A=>D(321));
   tri_F_322 : tri01 port map ( Y=>F(322), A=>nx5501, E=>nx5977);
   ix5502 : inv01 port map ( Y=>nx5501, A=>D(322));
   tri_F_323 : tri01 port map ( Y=>F(323), A=>nx5504, E=>nx5977);
   ix5505 : inv01 port map ( Y=>nx5504, A=>D(323));
   tri_F_324 : tri01 port map ( Y=>F(324), A=>nx5507, E=>nx5977);
   ix5508 : inv01 port map ( Y=>nx5507, A=>D(324));
   tri_F_325 : tri01 port map ( Y=>F(325), A=>nx5510, E=>nx5977);
   ix5511 : inv01 port map ( Y=>nx5510, A=>D(325));
   tri_F_326 : tri01 port map ( Y=>F(326), A=>nx5513, E=>nx5977);
   ix5514 : inv01 port map ( Y=>nx5513, A=>D(326));
   tri_F_327 : tri01 port map ( Y=>F(327), A=>nx5516, E=>nx5977);
   ix5517 : inv01 port map ( Y=>nx5516, A=>D(327));
   tri_F_328 : tri01 port map ( Y=>F(328), A=>nx5519, E=>nx5977);
   ix5520 : inv01 port map ( Y=>nx5519, A=>D(328));
   tri_F_329 : tri01 port map ( Y=>F(329), A=>nx5522, E=>nx5979);
   ix5523 : inv01 port map ( Y=>nx5522, A=>D(329));
   tri_F_330 : tri01 port map ( Y=>F(330), A=>nx5525, E=>nx5979);
   ix5526 : inv01 port map ( Y=>nx5525, A=>D(330));
   tri_F_331 : tri01 port map ( Y=>F(331), A=>nx5528, E=>nx5979);
   ix5529 : inv01 port map ( Y=>nx5528, A=>D(331));
   tri_F_332 : tri01 port map ( Y=>F(332), A=>nx5531, E=>nx5979);
   ix5532 : inv01 port map ( Y=>nx5531, A=>D(332));
   tri_F_333 : tri01 port map ( Y=>F(333), A=>nx5534, E=>nx5979);
   ix5535 : inv01 port map ( Y=>nx5534, A=>D(333));
   tri_F_334 : tri01 port map ( Y=>F(334), A=>nx5537, E=>nx5979);
   ix5538 : inv01 port map ( Y=>nx5537, A=>D(334));
   tri_F_335 : tri01 port map ( Y=>F(335), A=>nx5540, E=>nx5979);
   ix5541 : inv01 port map ( Y=>nx5540, A=>D(335));
   tri_F_336 : tri01 port map ( Y=>F(336), A=>nx5543, E=>nx5981);
   ix5544 : inv01 port map ( Y=>nx5543, A=>D(336));
   tri_F_337 : tri01 port map ( Y=>F(337), A=>nx5546, E=>nx5981);
   ix5547 : inv01 port map ( Y=>nx5546, A=>D(337));
   tri_F_338 : tri01 port map ( Y=>F(338), A=>nx5549, E=>nx5981);
   ix5550 : inv01 port map ( Y=>nx5549, A=>D(338));
   tri_F_339 : tri01 port map ( Y=>F(339), A=>nx5552, E=>nx5981);
   ix5553 : inv01 port map ( Y=>nx5552, A=>D(339));
   tri_F_340 : tri01 port map ( Y=>F(340), A=>nx5555, E=>nx5981);
   ix5556 : inv01 port map ( Y=>nx5555, A=>D(340));
   tri_F_341 : tri01 port map ( Y=>F(341), A=>nx5558, E=>nx5981);
   ix5559 : inv01 port map ( Y=>nx5558, A=>D(341));
   tri_F_342 : tri01 port map ( Y=>F(342), A=>nx5561, E=>nx5981);
   ix5562 : inv01 port map ( Y=>nx5561, A=>D(342));
   tri_F_343 : tri01 port map ( Y=>F(343), A=>nx5564, E=>nx5983);
   ix5565 : inv01 port map ( Y=>nx5564, A=>D(343));
   tri_F_344 : tri01 port map ( Y=>F(344), A=>nx5567, E=>nx5983);
   ix5568 : inv01 port map ( Y=>nx5567, A=>D(344));
   tri_F_345 : tri01 port map ( Y=>F(345), A=>nx5570, E=>nx5983);
   ix5571 : inv01 port map ( Y=>nx5570, A=>D(345));
   tri_F_346 : tri01 port map ( Y=>F(346), A=>nx5573, E=>nx5983);
   ix5574 : inv01 port map ( Y=>nx5573, A=>D(346));
   tri_F_347 : tri01 port map ( Y=>F(347), A=>nx5576, E=>nx5983);
   ix5577 : inv01 port map ( Y=>nx5576, A=>D(347));
   tri_F_348 : tri01 port map ( Y=>F(348), A=>nx5579, E=>nx5983);
   ix5580 : inv01 port map ( Y=>nx5579, A=>D(348));
   tri_F_349 : tri01 port map ( Y=>F(349), A=>nx5582, E=>nx5983);
   ix5583 : inv01 port map ( Y=>nx5582, A=>D(349));
   tri_F_350 : tri01 port map ( Y=>F(350), A=>nx5585, E=>nx5985);
   ix5586 : inv01 port map ( Y=>nx5585, A=>D(350));
   tri_F_351 : tri01 port map ( Y=>F(351), A=>nx5588, E=>nx5985);
   ix5589 : inv01 port map ( Y=>nx5588, A=>D(351));
   tri_F_352 : tri01 port map ( Y=>F(352), A=>nx5591, E=>nx5985);
   ix5592 : inv01 port map ( Y=>nx5591, A=>D(352));
   tri_F_353 : tri01 port map ( Y=>F(353), A=>nx5594, E=>nx5985);
   ix5595 : inv01 port map ( Y=>nx5594, A=>D(353));
   tri_F_354 : tri01 port map ( Y=>F(354), A=>nx5597, E=>nx5985);
   ix5598 : inv01 port map ( Y=>nx5597, A=>D(354));
   tri_F_355 : tri01 port map ( Y=>F(355), A=>nx5600, E=>nx5985);
   ix5601 : inv01 port map ( Y=>nx5600, A=>D(355));
   tri_F_356 : tri01 port map ( Y=>F(356), A=>nx5603, E=>nx5985);
   ix5604 : inv01 port map ( Y=>nx5603, A=>D(356));
   tri_F_357 : tri01 port map ( Y=>F(357), A=>nx5606, E=>nx5987);
   ix5607 : inv01 port map ( Y=>nx5606, A=>D(357));
   tri_F_358 : tri01 port map ( Y=>F(358), A=>nx5609, E=>nx5987);
   ix5610 : inv01 port map ( Y=>nx5609, A=>D(358));
   tri_F_359 : tri01 port map ( Y=>F(359), A=>nx5612, E=>nx5987);
   ix5613 : inv01 port map ( Y=>nx5612, A=>D(359));
   tri_F_360 : tri01 port map ( Y=>F(360), A=>nx5615, E=>nx5987);
   ix5616 : inv01 port map ( Y=>nx5615, A=>D(360));
   tri_F_361 : tri01 port map ( Y=>F(361), A=>nx5618, E=>nx5987);
   ix5619 : inv01 port map ( Y=>nx5618, A=>D(361));
   tri_F_362 : tri01 port map ( Y=>F(362), A=>nx5621, E=>nx5987);
   ix5622 : inv01 port map ( Y=>nx5621, A=>D(362));
   tri_F_363 : tri01 port map ( Y=>F(363), A=>nx5624, E=>nx5987);
   ix5625 : inv01 port map ( Y=>nx5624, A=>D(363));
   tri_F_364 : tri01 port map ( Y=>F(364), A=>nx5627, E=>nx5989);
   ix5628 : inv01 port map ( Y=>nx5627, A=>D(364));
   tri_F_365 : tri01 port map ( Y=>F(365), A=>nx5630, E=>nx5989);
   ix5631 : inv01 port map ( Y=>nx5630, A=>D(365));
   tri_F_366 : tri01 port map ( Y=>F(366), A=>nx5633, E=>nx5989);
   ix5634 : inv01 port map ( Y=>nx5633, A=>D(366));
   tri_F_367 : tri01 port map ( Y=>F(367), A=>nx5636, E=>nx5989);
   ix5637 : inv01 port map ( Y=>nx5636, A=>D(367));
   tri_F_368 : tri01 port map ( Y=>F(368), A=>nx5639, E=>nx5989);
   ix5640 : inv01 port map ( Y=>nx5639, A=>D(368));
   tri_F_369 : tri01 port map ( Y=>F(369), A=>nx5642, E=>nx5989);
   ix5643 : inv01 port map ( Y=>nx5642, A=>D(369));
   tri_F_370 : tri01 port map ( Y=>F(370), A=>nx5645, E=>nx5989);
   ix5646 : inv01 port map ( Y=>nx5645, A=>D(370));
   tri_F_371 : tri01 port map ( Y=>F(371), A=>nx5648, E=>nx5991);
   ix5649 : inv01 port map ( Y=>nx5648, A=>D(371));
   tri_F_372 : tri01 port map ( Y=>F(372), A=>nx5651, E=>nx5991);
   ix5652 : inv01 port map ( Y=>nx5651, A=>D(372));
   tri_F_373 : tri01 port map ( Y=>F(373), A=>nx5654, E=>nx5991);
   ix5655 : inv01 port map ( Y=>nx5654, A=>D(373));
   tri_F_374 : tri01 port map ( Y=>F(374), A=>nx5657, E=>nx5991);
   ix5658 : inv01 port map ( Y=>nx5657, A=>D(374));
   tri_F_375 : tri01 port map ( Y=>F(375), A=>nx5660, E=>nx5991);
   ix5661 : inv01 port map ( Y=>nx5660, A=>D(375));
   tri_F_376 : tri01 port map ( Y=>F(376), A=>nx5663, E=>nx5991);
   ix5664 : inv01 port map ( Y=>nx5663, A=>D(376));
   tri_F_377 : tri01 port map ( Y=>F(377), A=>nx5666, E=>nx5991);
   ix5667 : inv01 port map ( Y=>nx5666, A=>D(377));
   tri_F_378 : tri01 port map ( Y=>F(378), A=>nx5669, E=>nx5993);
   ix5670 : inv01 port map ( Y=>nx5669, A=>D(378));
   tri_F_379 : tri01 port map ( Y=>F(379), A=>nx5672, E=>nx5993);
   ix5673 : inv01 port map ( Y=>nx5672, A=>D(379));
   tri_F_380 : tri01 port map ( Y=>F(380), A=>nx5675, E=>nx5993);
   ix5676 : inv01 port map ( Y=>nx5675, A=>D(380));
   tri_F_381 : tri01 port map ( Y=>F(381), A=>nx5678, E=>nx5993);
   ix5679 : inv01 port map ( Y=>nx5678, A=>D(381));
   tri_F_382 : tri01 port map ( Y=>F(382), A=>nx5681, E=>nx5993);
   ix5682 : inv01 port map ( Y=>nx5681, A=>D(382));
   tri_F_383 : tri01 port map ( Y=>F(383), A=>nx5684, E=>nx5993);
   ix5685 : inv01 port map ( Y=>nx5684, A=>D(383));
   tri_F_384 : tri01 port map ( Y=>F(384), A=>nx5687, E=>nx5993);
   ix5688 : inv01 port map ( Y=>nx5687, A=>D(384));
   tri_F_385 : tri01 port map ( Y=>F(385), A=>nx5690, E=>nx5995);
   ix5691 : inv01 port map ( Y=>nx5690, A=>D(385));
   tri_F_386 : tri01 port map ( Y=>F(386), A=>nx5693, E=>nx5995);
   ix5694 : inv01 port map ( Y=>nx5693, A=>D(386));
   tri_F_387 : tri01 port map ( Y=>F(387), A=>nx5696, E=>nx5995);
   ix5697 : inv01 port map ( Y=>nx5696, A=>D(387));
   tri_F_388 : tri01 port map ( Y=>F(388), A=>nx5699, E=>nx5995);
   ix5700 : inv01 port map ( Y=>nx5699, A=>D(388));
   tri_F_389 : tri01 port map ( Y=>F(389), A=>nx5702, E=>nx5995);
   ix5703 : inv01 port map ( Y=>nx5702, A=>D(389));
   tri_F_390 : tri01 port map ( Y=>F(390), A=>nx5705, E=>nx5995);
   ix5706 : inv01 port map ( Y=>nx5705, A=>D(390));
   tri_F_391 : tri01 port map ( Y=>F(391), A=>nx5708, E=>nx5995);
   ix5709 : inv01 port map ( Y=>nx5708, A=>D(391));
   tri_F_392 : tri01 port map ( Y=>F(392), A=>nx5711, E=>nx5997);
   ix5712 : inv01 port map ( Y=>nx5711, A=>D(392));
   tri_F_393 : tri01 port map ( Y=>F(393), A=>nx5714, E=>nx5997);
   ix5715 : inv01 port map ( Y=>nx5714, A=>D(393));
   tri_F_394 : tri01 port map ( Y=>F(394), A=>nx5717, E=>nx5997);
   ix5718 : inv01 port map ( Y=>nx5717, A=>D(394));
   tri_F_395 : tri01 port map ( Y=>F(395), A=>nx5720, E=>nx5997);
   ix5721 : inv01 port map ( Y=>nx5720, A=>D(395));
   tri_F_396 : tri01 port map ( Y=>F(396), A=>nx5723, E=>nx5997);
   ix5724 : inv01 port map ( Y=>nx5723, A=>D(396));
   tri_F_397 : tri01 port map ( Y=>F(397), A=>nx5726, E=>nx5997);
   ix5727 : inv01 port map ( Y=>nx5726, A=>D(397));
   tri_F_398 : tri01 port map ( Y=>F(398), A=>nx5729, E=>nx5997);
   ix5730 : inv01 port map ( Y=>nx5729, A=>D(398));
   tri_F_399 : tri01 port map ( Y=>F(399), A=>nx5732, E=>nx5999);
   ix5733 : inv01 port map ( Y=>nx5732, A=>D(399));
   tri_F_400 : tri01 port map ( Y=>F(400), A=>nx5735, E=>nx5999);
   ix5736 : inv01 port map ( Y=>nx5735, A=>D(400));
   tri_F_401 : tri01 port map ( Y=>F(401), A=>nx5738, E=>nx5999);
   ix5739 : inv01 port map ( Y=>nx5738, A=>D(401));
   tri_F_402 : tri01 port map ( Y=>F(402), A=>nx5741, E=>nx5999);
   ix5742 : inv01 port map ( Y=>nx5741, A=>D(402));
   tri_F_403 : tri01 port map ( Y=>F(403), A=>nx5744, E=>nx5999);
   ix5745 : inv01 port map ( Y=>nx5744, A=>D(403));
   tri_F_404 : tri01 port map ( Y=>F(404), A=>nx5747, E=>nx5999);
   ix5748 : inv01 port map ( Y=>nx5747, A=>D(404));
   tri_F_405 : tri01 port map ( Y=>F(405), A=>nx5750, E=>nx5999);
   ix5751 : inv01 port map ( Y=>nx5750, A=>D(405));
   tri_F_406 : tri01 port map ( Y=>F(406), A=>nx5753, E=>nx6001);
   ix5754 : inv01 port map ( Y=>nx5753, A=>D(406));
   tri_F_407 : tri01 port map ( Y=>F(407), A=>nx5756, E=>nx6001);
   ix5757 : inv01 port map ( Y=>nx5756, A=>D(407));
   tri_F_408 : tri01 port map ( Y=>F(408), A=>nx5759, E=>nx6001);
   ix5760 : inv01 port map ( Y=>nx5759, A=>D(408));
   tri_F_409 : tri01 port map ( Y=>F(409), A=>nx5762, E=>nx6001);
   ix5763 : inv01 port map ( Y=>nx5762, A=>D(409));
   tri_F_410 : tri01 port map ( Y=>F(410), A=>nx5765, E=>nx6001);
   ix5766 : inv01 port map ( Y=>nx5765, A=>D(410));
   tri_F_411 : tri01 port map ( Y=>F(411), A=>nx5768, E=>nx6001);
   ix5769 : inv01 port map ( Y=>nx5768, A=>D(411));
   tri_F_412 : tri01 port map ( Y=>F(412), A=>nx5771, E=>nx6001);
   ix5772 : inv01 port map ( Y=>nx5771, A=>D(412));
   tri_F_413 : tri01 port map ( Y=>F(413), A=>nx5774, E=>nx6003);
   ix5775 : inv01 port map ( Y=>nx5774, A=>D(413));
   tri_F_414 : tri01 port map ( Y=>F(414), A=>nx5777, E=>nx6003);
   ix5778 : inv01 port map ( Y=>nx5777, A=>D(414));
   tri_F_415 : tri01 port map ( Y=>F(415), A=>nx5780, E=>nx6003);
   ix5781 : inv01 port map ( Y=>nx5780, A=>D(415));
   tri_F_416 : tri01 port map ( Y=>F(416), A=>nx5783, E=>nx6003);
   ix5784 : inv01 port map ( Y=>nx5783, A=>D(416));
   tri_F_417 : tri01 port map ( Y=>F(417), A=>nx5786, E=>nx6003);
   ix5787 : inv01 port map ( Y=>nx5786, A=>D(417));
   tri_F_418 : tri01 port map ( Y=>F(418), A=>nx5789, E=>nx6003);
   ix5790 : inv01 port map ( Y=>nx5789, A=>D(418));
   tri_F_419 : tri01 port map ( Y=>F(419), A=>nx5792, E=>nx6003);
   ix5793 : inv01 port map ( Y=>nx5792, A=>D(419));
   tri_F_420 : tri01 port map ( Y=>F(420), A=>nx5795, E=>nx6005);
   ix5796 : inv01 port map ( Y=>nx5795, A=>D(420));
   tri_F_421 : tri01 port map ( Y=>F(421), A=>nx5798, E=>nx6005);
   ix5799 : inv01 port map ( Y=>nx5798, A=>D(421));
   tri_F_422 : tri01 port map ( Y=>F(422), A=>nx5801, E=>nx6005);
   ix5802 : inv01 port map ( Y=>nx5801, A=>D(422));
   tri_F_423 : tri01 port map ( Y=>F(423), A=>nx5804, E=>nx6005);
   ix5805 : inv01 port map ( Y=>nx5804, A=>D(423));
   tri_F_424 : tri01 port map ( Y=>F(424), A=>nx5807, E=>nx6005);
   ix5808 : inv01 port map ( Y=>nx5807, A=>D(424));
   tri_F_425 : tri01 port map ( Y=>F(425), A=>nx5810, E=>nx6005);
   ix5811 : inv01 port map ( Y=>nx5810, A=>D(425));
   tri_F_426 : tri01 port map ( Y=>F(426), A=>nx5813, E=>nx6005);
   ix5814 : inv01 port map ( Y=>nx5813, A=>D(426));
   tri_F_427 : tri01 port map ( Y=>F(427), A=>nx5816, E=>nx6007);
   ix5817 : inv01 port map ( Y=>nx5816, A=>D(427));
   tri_F_428 : tri01 port map ( Y=>F(428), A=>nx5819, E=>nx6007);
   ix5820 : inv01 port map ( Y=>nx5819, A=>D(428));
   tri_F_429 : tri01 port map ( Y=>F(429), A=>nx5822, E=>nx6007);
   ix5823 : inv01 port map ( Y=>nx5822, A=>D(429));
   tri_F_430 : tri01 port map ( Y=>F(430), A=>nx5825, E=>nx6007);
   ix5826 : inv01 port map ( Y=>nx5825, A=>D(430));
   tri_F_431 : tri01 port map ( Y=>F(431), A=>nx5828, E=>nx6007);
   ix5829 : inv01 port map ( Y=>nx5828, A=>D(431));
   tri_F_432 : tri01 port map ( Y=>F(432), A=>nx5831, E=>nx6007);
   ix5832 : inv01 port map ( Y=>nx5831, A=>D(432));
   tri_F_433 : tri01 port map ( Y=>F(433), A=>nx5834, E=>nx6007);
   ix5835 : inv01 port map ( Y=>nx5834, A=>D(433));
   tri_F_434 : tri01 port map ( Y=>F(434), A=>nx5837, E=>nx6009);
   ix5838 : inv01 port map ( Y=>nx5837, A=>D(434));
   tri_F_435 : tri01 port map ( Y=>F(435), A=>nx5840, E=>nx6009);
   ix5841 : inv01 port map ( Y=>nx5840, A=>D(435));
   tri_F_436 : tri01 port map ( Y=>F(436), A=>nx5843, E=>nx6009);
   ix5844 : inv01 port map ( Y=>nx5843, A=>D(436));
   tri_F_437 : tri01 port map ( Y=>F(437), A=>nx5846, E=>nx6009);
   ix5847 : inv01 port map ( Y=>nx5846, A=>D(437));
   tri_F_438 : tri01 port map ( Y=>F(438), A=>nx5849, E=>nx6009);
   ix5850 : inv01 port map ( Y=>nx5849, A=>D(438));
   tri_F_439 : tri01 port map ( Y=>F(439), A=>nx5852, E=>nx6009);
   ix5853 : inv01 port map ( Y=>nx5852, A=>D(439));
   tri_F_440 : tri01 port map ( Y=>F(440), A=>nx5855, E=>nx6009);
   ix5856 : inv01 port map ( Y=>nx5855, A=>D(440));
   tri_F_441 : tri01 port map ( Y=>F(441), A=>nx5858, E=>nx6011);
   ix5859 : inv01 port map ( Y=>nx5858, A=>D(441));
   tri_F_442 : tri01 port map ( Y=>F(442), A=>nx5861, E=>nx6011);
   ix5862 : inv01 port map ( Y=>nx5861, A=>D(442));
   tri_F_443 : tri01 port map ( Y=>F(443), A=>nx5864, E=>nx6011);
   ix5865 : inv01 port map ( Y=>nx5864, A=>D(443));
   tri_F_444 : tri01 port map ( Y=>F(444), A=>nx5867, E=>nx6011);
   ix5868 : inv01 port map ( Y=>nx5867, A=>D(444));
   tri_F_445 : tri01 port map ( Y=>F(445), A=>nx5870, E=>nx6011);
   ix5871 : inv01 port map ( Y=>nx5870, A=>D(445));
   tri_F_446 : tri01 port map ( Y=>F(446), A=>nx5873, E=>nx6011);
   ix5874 : inv01 port map ( Y=>nx5873, A=>D(446));
   tri_F_447 : tri01 port map ( Y=>F(447), A=>nx5876, E=>nx6011);
   ix5877 : inv01 port map ( Y=>nx5876, A=>D(447));
   ix5882 : inv01 port map ( Y=>nx5883, A=>EN);
   ix5884 : inv01 port map ( Y=>nx5885, A=>nx6013);
   ix5886 : inv01 port map ( Y=>nx5887, A=>nx6013);
   ix5888 : inv01 port map ( Y=>nx5889, A=>nx6013);
   ix5890 : inv01 port map ( Y=>nx5891, A=>nx6013);
   ix5892 : inv01 port map ( Y=>nx5893, A=>nx6013);
   ix5894 : inv01 port map ( Y=>nx5895, A=>nx6013);
   ix5896 : inv01 port map ( Y=>nx5897, A=>nx6013);
   ix5898 : inv01 port map ( Y=>nx5899, A=>nx6015);
   ix5900 : inv01 port map ( Y=>nx5901, A=>nx6015);
   ix5902 : inv01 port map ( Y=>nx5903, A=>nx6015);
   ix5904 : inv01 port map ( Y=>nx5905, A=>nx6015);
   ix5906 : inv01 port map ( Y=>nx5907, A=>nx6015);
   ix5908 : inv01 port map ( Y=>nx5909, A=>nx6015);
   ix5910 : inv01 port map ( Y=>nx5911, A=>nx6015);
   ix5912 : inv01 port map ( Y=>nx5913, A=>nx6017);
   ix5914 : inv01 port map ( Y=>nx5915, A=>nx6017);
   ix5916 : inv01 port map ( Y=>nx5917, A=>nx6017);
   ix5918 : inv01 port map ( Y=>nx5919, A=>nx6017);
   ix5920 : inv01 port map ( Y=>nx5921, A=>nx6017);
   ix5922 : inv01 port map ( Y=>nx5923, A=>nx6017);
   ix5924 : inv01 port map ( Y=>nx5925, A=>nx6017);
   ix5926 : inv01 port map ( Y=>nx5927, A=>nx6019);
   ix5928 : inv01 port map ( Y=>nx5929, A=>nx6019);
   ix5930 : inv01 port map ( Y=>nx5931, A=>nx6019);
   ix5932 : inv01 port map ( Y=>nx5933, A=>nx6019);
   ix5934 : inv01 port map ( Y=>nx5935, A=>nx6019);
   ix5936 : inv01 port map ( Y=>nx5937, A=>nx6019);
   ix5938 : inv01 port map ( Y=>nx5939, A=>nx6019);
   ix5940 : inv01 port map ( Y=>nx5941, A=>nx6021);
   ix5942 : inv01 port map ( Y=>nx5943, A=>nx6021);
   ix5944 : inv01 port map ( Y=>nx5945, A=>nx6021);
   ix5946 : inv01 port map ( Y=>nx5947, A=>nx6021);
   ix5948 : inv01 port map ( Y=>nx5949, A=>nx6021);
   ix5950 : inv01 port map ( Y=>nx5951, A=>nx6021);
   ix5952 : inv01 port map ( Y=>nx5953, A=>nx6021);
   ix5954 : inv01 port map ( Y=>nx5955, A=>nx6023);
   ix5956 : inv01 port map ( Y=>nx5957, A=>nx6023);
   ix5958 : inv01 port map ( Y=>nx5959, A=>nx6023);
   ix5960 : inv01 port map ( Y=>nx5961, A=>nx6023);
   ix5962 : inv01 port map ( Y=>nx5963, A=>nx6023);
   ix5964 : inv01 port map ( Y=>nx5965, A=>nx6023);
   ix5966 : inv01 port map ( Y=>nx5967, A=>nx6023);
   ix5968 : inv01 port map ( Y=>nx5969, A=>nx6025);
   ix5970 : inv01 port map ( Y=>nx5971, A=>nx6025);
   ix5972 : inv01 port map ( Y=>nx5973, A=>nx6025);
   ix5974 : inv01 port map ( Y=>nx5975, A=>nx6025);
   ix5976 : inv01 port map ( Y=>nx5977, A=>nx6025);
   ix5978 : inv01 port map ( Y=>nx5979, A=>nx6025);
   ix5980 : inv01 port map ( Y=>nx5981, A=>nx6025);
   ix5982 : inv01 port map ( Y=>nx5983, A=>nx6027);
   ix5984 : inv01 port map ( Y=>nx5985, A=>nx6027);
   ix5986 : inv01 port map ( Y=>nx5987, A=>nx6027);
   ix5988 : inv01 port map ( Y=>nx5989, A=>nx6027);
   ix5990 : inv01 port map ( Y=>nx5991, A=>nx6027);
   ix5992 : inv01 port map ( Y=>nx5993, A=>nx6027);
   ix5994 : inv01 port map ( Y=>nx5995, A=>nx6027);
   ix5996 : inv01 port map ( Y=>nx5997, A=>nx6029);
   ix5998 : inv01 port map ( Y=>nx5999, A=>nx6029);
   ix6000 : inv01 port map ( Y=>nx6001, A=>nx6029);
   ix6002 : inv01 port map ( Y=>nx6003, A=>nx6029);
   ix6004 : inv01 port map ( Y=>nx6005, A=>nx6029);
   ix6006 : inv01 port map ( Y=>nx6007, A=>nx6029);
   ix6008 : inv01 port map ( Y=>nx6009, A=>nx6029);
   ix6010 : inv01 port map ( Y=>nx6011, A=>nx5883);
   ix6012 : inv01 port map ( Y=>nx6013, A=>nx6035);
   ix6014 : inv01 port map ( Y=>nx6015, A=>nx6035);
   ix6016 : inv01 port map ( Y=>nx6017, A=>nx6035);
   ix6018 : inv01 port map ( Y=>nx6019, A=>nx6035);
   ix6020 : inv01 port map ( Y=>nx6021, A=>nx6035);
   ix6022 : inv01 port map ( Y=>nx6023, A=>nx6035);
   ix6024 : inv01 port map ( Y=>nx6025, A=>nx6035);
   ix6026 : inv01 port map ( Y=>nx6027, A=>nx6037);
   ix6028 : inv01 port map ( Y=>nx6029, A=>nx6037);
   ix6034 : inv01 port map ( Y=>nx6035, A=>nx5883);
   ix6036 : inv01 port map ( Y=>nx6037, A=>nx5883);
end triBuffer ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity triStateBuffer_16 is
   port (
      D : IN std_logic_vector (15 DOWNTO 0) ;
      EN : IN std_logic ;
      F : OUT std_logic_vector (15 DOWNTO 0)) ;
end triStateBuffer_16 ;

architecture triBuffer of triStateBuffer_16 is
   signal nx215, nx218, nx221, nx224, nx227, nx230, nx233, nx236, nx239, 
      nx242, nx245, nx248, nx251, nx254, nx257, nx260, nx267, nx269, nx271, 
      nx273: std_logic ;

begin
   tri_F_0 : tri01 port map ( Y=>F(0), A=>nx215, E=>nx269);
   ix216 : inv01 port map ( Y=>nx215, A=>D(0));
   tri_F_1 : tri01 port map ( Y=>F(1), A=>nx218, E=>nx269);
   ix219 : inv01 port map ( Y=>nx218, A=>D(1));
   tri_F_2 : tri01 port map ( Y=>F(2), A=>nx221, E=>nx269);
   ix222 : inv01 port map ( Y=>nx221, A=>D(2));
   tri_F_3 : tri01 port map ( Y=>F(3), A=>nx224, E=>nx269);
   ix225 : inv01 port map ( Y=>nx224, A=>D(3));
   tri_F_4 : tri01 port map ( Y=>F(4), A=>nx227, E=>nx269);
   ix228 : inv01 port map ( Y=>nx227, A=>D(4));
   tri_F_5 : tri01 port map ( Y=>F(5), A=>nx230, E=>nx269);
   ix231 : inv01 port map ( Y=>nx230, A=>D(5));
   tri_F_6 : tri01 port map ( Y=>F(6), A=>nx233, E=>nx269);
   ix234 : inv01 port map ( Y=>nx233, A=>D(6));
   tri_F_7 : tri01 port map ( Y=>F(7), A=>nx236, E=>nx271);
   ix237 : inv01 port map ( Y=>nx236, A=>D(7));
   tri_F_8 : tri01 port map ( Y=>F(8), A=>nx239, E=>nx271);
   ix240 : inv01 port map ( Y=>nx239, A=>D(8));
   tri_F_9 : tri01 port map ( Y=>F(9), A=>nx242, E=>nx271);
   ix243 : inv01 port map ( Y=>nx242, A=>D(9));
   tri_F_10 : tri01 port map ( Y=>F(10), A=>nx245, E=>nx271);
   ix246 : inv01 port map ( Y=>nx245, A=>D(10));
   tri_F_11 : tri01 port map ( Y=>F(11), A=>nx248, E=>nx271);
   ix249 : inv01 port map ( Y=>nx248, A=>D(11));
   tri_F_12 : tri01 port map ( Y=>F(12), A=>nx251, E=>nx271);
   ix252 : inv01 port map ( Y=>nx251, A=>D(12));
   tri_F_13 : tri01 port map ( Y=>F(13), A=>nx254, E=>nx271);
   ix255 : inv01 port map ( Y=>nx254, A=>D(13));
   tri_F_14 : tri01 port map ( Y=>F(14), A=>nx257, E=>nx273);
   ix258 : inv01 port map ( Y=>nx257, A=>D(14));
   tri_F_15 : tri01 port map ( Y=>F(15), A=>nx260, E=>nx273);
   ix261 : inv01 port map ( Y=>nx260, A=>D(15));
   ix266 : inv01 port map ( Y=>nx267, A=>EN);
   ix268 : inv01 port map ( Y=>nx269, A=>nx267);
   ix270 : inv01 port map ( Y=>nx271, A=>nx267);
   ix272 : inv01 port map ( Y=>nx273, A=>nx267);
end triBuffer ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;
use ieee.numeric_std.all;

entity RAM_28 is
   port (
      reset : IN std_logic ;
      CLK : IN std_logic ;
      W : IN std_logic ;
      R : IN std_logic ;
      address : IN std_logic_vector (12 DOWNTO 0) ;
      dataIn : IN std_logic_vector (15 DOWNTO 0) ;
      dataOut : OUT std_logic_vector (447 DOWNTO 0) ;
      MFC : OUT std_logic ;
      counterOut : OUT std_logic_vector (3 DOWNTO 0)) ;
end RAM_28 ;

architecture archRAM of RAM_28 is
   type ram_type is array( 0 to 5000) of std_logic_vector(15 downto 0);
   signal ram: ram_type;
   signal mfc_m:std_logic;
   signal CLKEvent: std_logic;
   signal cReset,cEnable:std_logic;
   signal cOutput:std_logic_vector(3 downto 0);
   component Counter is
       generic(n: integer := 16);
       port(
           enable:in std_logic;
           reset:in std_logic;
           clk:in std_logic;
           load:in std_logic;
           output:out std_logic_vector(n-1 downto 0);
           input:in std_logic_vector(n-1 downto 0));
   end component;

begin
   -- enable the register when w or r signal comes
   cEnable <= '1' when (((W =  '1') or (R = '1')) and (mfc_m = '0'))
   else '0';
   counterOut <= cOutput;
   c1: Counter 
   generic map(4)
   port map(cEnable,cReset,CLK,'0',cOutput,"0001");

   -- MFC appears one clock after 8th clocks
   MFC <= mfc_m;
   --CLKEvent<= '1' when (CLK'event and CLK = '1')  else '0';
   
   mfc_m <= '1' when (cOutput = "0010" and(CLK'event and CLK = '1'))
   else '0' when   (CLK'event and CLK = '1');

   -- reset the counter when comes to 8 or a signal read or write
   cReset <= '1' when ((reset = '1') or (cOutput = "0011")) -- or (W'event and W = '1') or (R'event and R = '1') )
    else '0';

   -- memory retrieve 28 pixel of data after 8 bits
   process(cOutput)
  variable k,j,adds:integer;
   begin
       k := -16;
       j := -1;
       if  (cOutput = "0011" and W = '1')then
           ram(to_integer(unsigned(address))) <= dataIn;
       elsif  (cOutput = "0011" and R = '1')then
           loop1: for i in 0 to 27 loop
               k := k + 16;
               j := j + 16;
            adds := i + to_integer(unsigned(address));
               dataOut(j downto k) <= ram(adds);
         end loop;

--- we need to output z when we dont have data
       end if ;
   end process;
   end archRAM ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;
use ieee.numeric_std.all;

entity memoryDMA is
   port (
      resetEN : IN std_logic ;
      AddressIn : IN std_logic_vector (12 DOWNTO 0) ;
      dataIn : IN std_logic_vector (15 DOWNTO 0) ;
      switcherEN : IN std_logic ;
      ramSelector : IN std_logic ;
      readEn : IN std_logic ;
      writeEn : IN std_logic ;
      CLK : IN std_logic ;
      Normal : IN std_logic ;
      MFC : OUT std_logic ;
      counterOut : OUT std_logic_vector (3 DOWNTO 0) ;
      dataOut : OUT std_logic_vector (447 DOWNTO 0)) ;
end memoryDMA ;

architecture DMAmemory of memoryDMA is
   component triStateBuffer_448
      port (
         D : IN std_logic_vector (447 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (447 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component RAM_28
      port (
         reset : IN std_logic ;
         CLK : IN std_logic ;
         W : IN std_logic ;
         R : IN std_logic ;
         address : IN std_logic_vector (12 DOWNTO 0) ;
         dataIn : IN std_logic_vector (15 DOWNTO 0) ;
         dataOut : OUT std_logic_vector (447 DOWNTO 0) ;
         MFC : OUT std_logic ;
         counterOut : OUT std_logic_vector (3 DOWNTO 0)) ;
   end component ;
   signal dataOut_447_EXMPLR, dataOut_446_EXMPLR, dataOut_445_EXMPLR, 
      dataOut_444_EXMPLR, dataOut_443_EXMPLR, dataOut_442_EXMPLR, 
      dataOut_441_EXMPLR, dataOut_440_EXMPLR, dataOut_439_EXMPLR, 
      dataOut_438_EXMPLR, dataOut_437_EXMPLR, dataOut_436_EXMPLR, 
      dataOut_435_EXMPLR, dataOut_434_EXMPLR, dataOut_433_EXMPLR, 
      dataOut_432_EXMPLR, dataOut_431_EXMPLR, dataOut_430_EXMPLR, 
      dataOut_429_EXMPLR, dataOut_428_EXMPLR, dataOut_427_EXMPLR, 
      dataOut_426_EXMPLR, dataOut_425_EXMPLR, dataOut_424_EXMPLR, 
      dataOut_423_EXMPLR, dataOut_422_EXMPLR, dataOut_421_EXMPLR, 
      dataOut_420_EXMPLR, dataOut_419_EXMPLR, dataOut_418_EXMPLR, 
      dataOut_417_EXMPLR, dataOut_416_EXMPLR, dataOut_415_EXMPLR, 
      dataOut_414_EXMPLR, dataOut_413_EXMPLR, dataOut_412_EXMPLR, 
      dataOut_411_EXMPLR, dataOut_410_EXMPLR, dataOut_409_EXMPLR, 
      dataOut_408_EXMPLR, dataOut_407_EXMPLR, dataOut_406_EXMPLR, 
      dataOut_405_EXMPLR, dataOut_404_EXMPLR, dataOut_403_EXMPLR, 
      dataOut_402_EXMPLR, dataOut_401_EXMPLR, dataOut_400_EXMPLR, 
      dataOut_399_EXMPLR, dataOut_398_EXMPLR, dataOut_397_EXMPLR, 
      dataOut_396_EXMPLR, dataOut_395_EXMPLR, dataOut_394_EXMPLR, 
      dataOut_393_EXMPLR, dataOut_392_EXMPLR, dataOut_391_EXMPLR, 
      dataOut_390_EXMPLR, dataOut_389_EXMPLR, dataOut_388_EXMPLR, 
      dataOut_387_EXMPLR, dataOut_386_EXMPLR, dataOut_385_EXMPLR, 
      dataOut_384_EXMPLR, dataOut_383_EXMPLR, dataOut_382_EXMPLR, 
      dataOut_381_EXMPLR, dataOut_380_EXMPLR, dataOut_379_EXMPLR, 
      dataOut_378_EXMPLR, dataOut_377_EXMPLR, dataOut_376_EXMPLR, 
      dataOut_375_EXMPLR, dataOut_374_EXMPLR, dataOut_373_EXMPLR, 
      dataOut_372_EXMPLR, dataOut_371_EXMPLR, dataOut_370_EXMPLR, 
      dataOut_369_EXMPLR, dataOut_368_EXMPLR, dataOut_367_EXMPLR, 
      dataOut_366_EXMPLR, dataOut_365_EXMPLR, dataOut_364_EXMPLR, 
      dataOut_363_EXMPLR, dataOut_362_EXMPLR, dataOut_361_EXMPLR, 
      dataOut_360_EXMPLR, dataOut_359_EXMPLR, dataOut_358_EXMPLR, 
      dataOut_357_EXMPLR, dataOut_356_EXMPLR, dataOut_355_EXMPLR, 
      dataOut_354_EXMPLR, dataOut_353_EXMPLR, dataOut_352_EXMPLR, 
      dataOut_351_EXMPLR, dataOut_350_EXMPLR, dataOut_349_EXMPLR, 
      dataOut_348_EXMPLR, dataOut_347_EXMPLR, dataOut_346_EXMPLR, 
      dataOut_345_EXMPLR, dataOut_344_EXMPLR, dataOut_343_EXMPLR, 
      dataOut_342_EXMPLR, dataOut_341_EXMPLR, dataOut_340_EXMPLR, 
      dataOut_339_EXMPLR, dataOut_338_EXMPLR, dataOut_337_EXMPLR, 
      dataOut_336_EXMPLR, dataOut_335_EXMPLR, dataOut_334_EXMPLR, 
      dataOut_333_EXMPLR, dataOut_332_EXMPLR, dataOut_331_EXMPLR, 
      dataOut_330_EXMPLR, dataOut_329_EXMPLR, dataOut_328_EXMPLR, 
      dataOut_327_EXMPLR, dataOut_326_EXMPLR, dataOut_325_EXMPLR, 
      dataOut_324_EXMPLR, dataOut_323_EXMPLR, dataOut_322_EXMPLR, 
      dataOut_321_EXMPLR, dataOut_320_EXMPLR, dataOut_319_EXMPLR, 
      dataOut_318_EXMPLR, dataOut_317_EXMPLR, dataOut_316_EXMPLR, 
      dataOut_315_EXMPLR, dataOut_314_EXMPLR, dataOut_313_EXMPLR, 
      dataOut_312_EXMPLR, dataOut_311_EXMPLR, dataOut_310_EXMPLR, 
      dataOut_309_EXMPLR, dataOut_308_EXMPLR, dataOut_307_EXMPLR, 
      dataOut_306_EXMPLR, dataOut_305_EXMPLR, dataOut_304_EXMPLR, 
      dataOut_303_EXMPLR, dataOut_302_EXMPLR, dataOut_301_EXMPLR, 
      dataOut_300_EXMPLR, dataOut_299_EXMPLR, dataOut_298_EXMPLR, 
      dataOut_297_EXMPLR, dataOut_296_EXMPLR, dataOut_295_EXMPLR, 
      dataOut_294_EXMPLR, dataOut_293_EXMPLR, dataOut_292_EXMPLR, 
      dataOut_291_EXMPLR, dataOut_290_EXMPLR, dataOut_289_EXMPLR, 
      dataOut_288_EXMPLR, dataOut_287_EXMPLR, dataOut_286_EXMPLR, 
      dataOut_285_EXMPLR, dataOut_284_EXMPLR, dataOut_283_EXMPLR, 
      dataOut_282_EXMPLR, dataOut_281_EXMPLR, dataOut_280_EXMPLR, 
      dataOut_279_EXMPLR, dataOut_278_EXMPLR, dataOut_277_EXMPLR, 
      dataOut_276_EXMPLR, dataOut_275_EXMPLR, dataOut_274_EXMPLR, 
      dataOut_273_EXMPLR, dataOut_272_EXMPLR, dataOut_271_EXMPLR, 
      dataOut_270_EXMPLR, dataOut_269_EXMPLR, dataOut_268_EXMPLR, 
      dataOut_267_EXMPLR, dataOut_266_EXMPLR, dataOut_265_EXMPLR, 
      dataOut_264_EXMPLR, dataOut_263_EXMPLR, dataOut_262_EXMPLR, 
      dataOut_261_EXMPLR, dataOut_260_EXMPLR, dataOut_259_EXMPLR, 
      dataOut_258_EXMPLR, dataOut_257_EXMPLR, dataOut_256_EXMPLR, 
      dataOut_255_EXMPLR, dataOut_254_EXMPLR, dataOut_253_EXMPLR, 
      dataOut_252_EXMPLR, dataOut_251_EXMPLR, dataOut_250_EXMPLR, 
      dataOut_249_EXMPLR, dataOut_248_EXMPLR, dataOut_247_EXMPLR, 
      dataOut_246_EXMPLR, dataOut_245_EXMPLR, dataOut_244_EXMPLR, 
      dataOut_243_EXMPLR, dataOut_242_EXMPLR, dataOut_241_EXMPLR, 
      dataOut_240_EXMPLR, dataOut_239_EXMPLR, dataOut_238_EXMPLR, 
      dataOut_237_EXMPLR, dataOut_236_EXMPLR, dataOut_235_EXMPLR, 
      dataOut_234_EXMPLR, dataOut_233_EXMPLR, dataOut_232_EXMPLR, 
      dataOut_231_EXMPLR, dataOut_230_EXMPLR, dataOut_229_EXMPLR, 
      dataOut_228_EXMPLR, dataOut_227_EXMPLR, dataOut_226_EXMPLR, 
      dataOut_225_EXMPLR, dataOut_224_EXMPLR, dataOut_223_EXMPLR, 
      dataOut_222_EXMPLR, dataOut_221_EXMPLR, dataOut_220_EXMPLR, 
      dataOut_219_EXMPLR, dataOut_218_EXMPLR, dataOut_217_EXMPLR, 
      dataOut_216_EXMPLR, dataOut_215_EXMPLR, dataOut_214_EXMPLR, 
      dataOut_213_EXMPLR, dataOut_212_EXMPLR, dataOut_211_EXMPLR, 
      dataOut_210_EXMPLR, dataOut_209_EXMPLR, dataOut_208_EXMPLR, 
      dataOut_207_EXMPLR, dataOut_206_EXMPLR, dataOut_205_EXMPLR, 
      dataOut_204_EXMPLR, dataOut_203_EXMPLR, dataOut_202_EXMPLR, 
      dataOut_201_EXMPLR, dataOut_200_EXMPLR, dataOut_199_EXMPLR, 
      dataOut_198_EXMPLR, dataOut_197_EXMPLR, dataOut_196_EXMPLR, 
      dataOut_195_EXMPLR, dataOut_194_EXMPLR, dataOut_193_EXMPLR, 
      dataOut_192_EXMPLR, dataOut_191_EXMPLR, dataOut_190_EXMPLR, 
      dataOut_189_EXMPLR, dataOut_188_EXMPLR, dataOut_187_EXMPLR, 
      dataOut_186_EXMPLR, dataOut_185_EXMPLR, dataOut_184_EXMPLR, 
      dataOut_183_EXMPLR, dataOut_182_EXMPLR, dataOut_181_EXMPLR, 
      dataOut_180_EXMPLR, dataOut_179_EXMPLR, dataOut_178_EXMPLR, 
      dataOut_177_EXMPLR, dataOut_176_EXMPLR, dataOut_175_EXMPLR, 
      dataOut_174_EXMPLR, dataOut_173_EXMPLR, dataOut_172_EXMPLR, 
      dataOut_171_EXMPLR, dataOut_170_EXMPLR, dataOut_169_EXMPLR, 
      dataOut_168_EXMPLR, dataOut_167_EXMPLR, dataOut_166_EXMPLR, 
      dataOut_165_EXMPLR, dataOut_164_EXMPLR, dataOut_163_EXMPLR, 
      dataOut_162_EXMPLR, dataOut_161_EXMPLR, dataOut_160_EXMPLR, 
      dataOut_159_EXMPLR, dataOut_158_EXMPLR, dataOut_157_EXMPLR, 
      dataOut_156_EXMPLR, dataOut_155_EXMPLR, dataOut_154_EXMPLR, 
      dataOut_153_EXMPLR, dataOut_152_EXMPLR, dataOut_151_EXMPLR, 
      dataOut_150_EXMPLR, dataOut_149_EXMPLR, dataOut_148_EXMPLR, 
      dataOut_147_EXMPLR, dataOut_146_EXMPLR, dataOut_145_EXMPLR, 
      dataOut_144_EXMPLR, dataOut_143_EXMPLR, dataOut_142_EXMPLR, 
      dataOut_141_EXMPLR, dataOut_140_EXMPLR, dataOut_139_EXMPLR, 
      dataOut_138_EXMPLR, dataOut_137_EXMPLR, dataOut_136_EXMPLR, 
      dataOut_135_EXMPLR, dataOut_134_EXMPLR, dataOut_133_EXMPLR, 
      dataOut_132_EXMPLR, dataOut_131_EXMPLR, dataOut_130_EXMPLR, 
      dataOut_129_EXMPLR, dataOut_128_EXMPLR, dataOut_127_EXMPLR, 
      dataOut_126_EXMPLR, dataOut_125_EXMPLR, dataOut_124_EXMPLR, 
      dataOut_123_EXMPLR, dataOut_122_EXMPLR, dataOut_121_EXMPLR, 
      dataOut_120_EXMPLR, dataOut_119_EXMPLR, dataOut_118_EXMPLR, 
      dataOut_117_EXMPLR, dataOut_116_EXMPLR, dataOut_115_EXMPLR, 
      dataOut_114_EXMPLR, dataOut_113_EXMPLR, dataOut_112_EXMPLR, 
      dataOut_111_EXMPLR, dataOut_110_EXMPLR, dataOut_109_EXMPLR, 
      dataOut_108_EXMPLR, dataOut_107_EXMPLR, dataOut_106_EXMPLR, 
      dataOut_105_EXMPLR, dataOut_104_EXMPLR, dataOut_103_EXMPLR, 
      dataOut_102_EXMPLR, dataOut_101_EXMPLR, dataOut_100_EXMPLR, 
      dataOut_99_EXMPLR, dataOut_98_EXMPLR, dataOut_97_EXMPLR, 
      dataOut_96_EXMPLR, dataOut_95_EXMPLR, dataOut_94_EXMPLR, 
      dataOut_93_EXMPLR, dataOut_92_EXMPLR, dataOut_91_EXMPLR, 
      dataOut_90_EXMPLR, dataOut_89_EXMPLR, dataOut_88_EXMPLR, 
      dataOut_87_EXMPLR, dataOut_86_EXMPLR, dataOut_85_EXMPLR, 
      dataOut_84_EXMPLR, dataOut_83_EXMPLR, dataOut_82_EXMPLR, 
      dataOut_81_EXMPLR, dataOut_80_EXMPLR, dataOut_79_EXMPLR, 
      dataOut_78_EXMPLR, dataOut_77_EXMPLR, dataOut_76_EXMPLR, 
      dataOut_75_EXMPLR, dataOut_74_EXMPLR, dataOut_73_EXMPLR, 
      dataOut_72_EXMPLR, dataOut_71_EXMPLR, dataOut_70_EXMPLR, 
      dataOut_69_EXMPLR, dataOut_68_EXMPLR, dataOut_67_EXMPLR, 
      dataOut_66_EXMPLR, dataOut_65_EXMPLR, dataOut_64_EXMPLR, 
      dataOut_63_EXMPLR, dataOut_62_EXMPLR, dataOut_61_EXMPLR, 
      dataOut_60_EXMPLR, dataOut_59_EXMPLR, dataOut_58_EXMPLR, 
      dataOut_57_EXMPLR, dataOut_56_EXMPLR, dataOut_55_EXMPLR, 
      dataOut_54_EXMPLR, dataOut_53_EXMPLR, dataOut_52_EXMPLR, 
      dataOut_51_EXMPLR, dataOut_50_EXMPLR, dataOut_49_EXMPLR, 
      dataOut_48_EXMPLR, dataOut_47_EXMPLR, dataOut_46_EXMPLR, 
      dataOut_45_EXMPLR, dataOut_44_EXMPLR, dataOut_43_EXMPLR, 
      dataOut_42_EXMPLR, dataOut_41_EXMPLR, dataOut_40_EXMPLR, 
      dataOut_39_EXMPLR, dataOut_38_EXMPLR, dataOut_37_EXMPLR, 
      dataOut_36_EXMPLR, dataOut_35_EXMPLR, dataOut_34_EXMPLR, 
      dataOut_33_EXMPLR, dataOut_32_EXMPLR, dataOut_31_EXMPLR, 
      dataOut_30_EXMPLR, dataOut_29_EXMPLR, dataOut_28_EXMPLR, 
      dataOut_27_EXMPLR, dataOut_26_EXMPLR, dataOut_25_EXMPLR, 
      dataOut_24_EXMPLR, dataOut_23_EXMPLR, dataOut_22_EXMPLR, 
      dataOut_21_EXMPLR, dataOut_20_EXMPLR, dataOut_19_EXMPLR, 
      dataOut_18_EXMPLR, dataOut_17_EXMPLR, dataOut_16_EXMPLR, 
      dataOut_15_EXMPLR, dataOut_14_EXMPLR, dataOut_13_EXMPLR, 
      dataOut_12_EXMPLR, dataOut_11_EXMPLR, dataOut_10_EXMPLR, 
      dataOut_9_EXMPLR, dataOut_8_EXMPLR, dataOut_7_EXMPLR, dataOut_6_EXMPLR, 
      dataOut_5_EXMPLR, dataOut_4_EXMPLR, dataOut_3_EXMPLR, dataOut_2_EXMPLR, 
      dataOut_1_EXMPLR, dataOut_0_EXMPLR, dataFromRam1_447, dataFromRam2_447, 
      dataToRam1_15, dataToRam1_14, dataToRam1_13, dataToRam1_12, 
      dataToRam1_11, dataToRam1_10, dataToRam1_9, dataToRam1_8, dataToRam1_7, 
      dataToRam1_6, dataToRam1_5, dataToRam1_4, dataToRam1_3, dataToRam1_2, 
      dataToRam1_1, dataToRam1_0, dataToRam2_15, dataToRam2_14, 
      dataToRam2_13, dataToRam2_12, dataToRam2_11, dataToRam2_10, 
      dataToRam2_9, dataToRam2_8, dataToRam2_7, dataToRam2_6, dataToRam2_5, 
      dataToRam2_4, dataToRam2_3, dataToRam2_2, dataToRam2_1, dataToRam2_0, 
      mfcOfRam1, mfcOfRam2, DInput, ram2Read, ram1Read, ram2Write, ram1Write, 
      GND, test, nx5632, nx5653, nx5655, nx5657, nx5659, nx5661, nx5663, 
      nx5665, nx5667, nx5669, nx5671, nx5673, nx5675, nx5677, nx5679, nx5681, 
      nx5683, nx5685, nx5687, nx5689, nx5691, nx5693, nx5695, nx5697, nx5699, 
      nx5701, nx5703, nx5705, nx5707, nx5709, nx5711, nx5713, nx5715, nx5717, 
      nx5719, nx5721, nx5723, nx5725, nx5727, nx5729, nx5731, nx5733, nx5735, 
      nx5737, nx5739, nx5741, nx5743, nx5745, nx5747, nx5749, nx5751, nx5753, 
      nx5755, nx5757, nx5759, nx5761, nx5763, nx5765, nx5767, nx5769, nx5771, 
      nx5773, nx5775, nx5777, nx5779, nx5781, nx5783, nx5785, nx5787, nx5789, 
      nx5791, nx5793, nx5795, nx5797, nx5799, nx5801, nx5803, nx5805, nx5807, 
      nx5809, nx5811, nx5813, nx5815, nx5817, nx5819, nx5821, nx5823, nx5825, 
      nx5827, nx5829, nx5831, nx5833, nx5835, nx5837, nx5839, nx5841, nx5843, 
      nx5845, nx5847, nx5849, nx5851, nx5853, nx5855, nx5857, nx5859, nx5861, 
      nx5863, nx5865, nx5867, nx5869, nx5871, nx5873, nx5875, nx5877, nx5879, 
      nx5881, nx5883, nx5885, nx5887, nx5889, nx5891, nx5893, nx5895, nx5897, 
      nx5899, nx5901, nx5903, nx5905, nx5907, nx5909, nx5911, nx5913, nx5915, 
      nx5917, nx5919, nx5921, nx5923, nx5925, nx5927, nx5929, nx5931, nx5933, 
      nx5935, nx5937, nx5939, nx5941, nx5943, nx5945, nx5947, nx5953, nx5955, 
      nx5957, nx5959: std_logic ;
   
   signal DANGLING : std_logic_vector (901 downto 0 );

begin
   dataOut(447) <= dataOut_447_EXMPLR ;
   dataOut(446) <= dataOut_446_EXMPLR ;
   dataOut(445) <= dataOut_445_EXMPLR ;
   dataOut(444) <= dataOut_444_EXMPLR ;
   dataOut(443) <= dataOut_443_EXMPLR ;
   dataOut(442) <= dataOut_442_EXMPLR ;
   dataOut(441) <= dataOut_441_EXMPLR ;
   dataOut(440) <= dataOut_440_EXMPLR ;
   dataOut(439) <= dataOut_439_EXMPLR ;
   dataOut(438) <= dataOut_438_EXMPLR ;
   dataOut(437) <= dataOut_437_EXMPLR ;
   dataOut(436) <= dataOut_436_EXMPLR ;
   dataOut(435) <= dataOut_435_EXMPLR ;
   dataOut(434) <= dataOut_434_EXMPLR ;
   dataOut(433) <= dataOut_433_EXMPLR ;
   dataOut(432) <= dataOut_432_EXMPLR ;
   dataOut(431) <= dataOut_431_EXMPLR ;
   dataOut(430) <= dataOut_430_EXMPLR ;
   dataOut(429) <= dataOut_429_EXMPLR ;
   dataOut(428) <= dataOut_428_EXMPLR ;
   dataOut(427) <= dataOut_427_EXMPLR ;
   dataOut(426) <= dataOut_426_EXMPLR ;
   dataOut(425) <= dataOut_425_EXMPLR ;
   dataOut(424) <= dataOut_424_EXMPLR ;
   dataOut(423) <= dataOut_423_EXMPLR ;
   dataOut(422) <= dataOut_422_EXMPLR ;
   dataOut(421) <= dataOut_421_EXMPLR ;
   dataOut(420) <= dataOut_420_EXMPLR ;
   dataOut(419) <= dataOut_419_EXMPLR ;
   dataOut(418) <= dataOut_418_EXMPLR ;
   dataOut(417) <= dataOut_417_EXMPLR ;
   dataOut(416) <= dataOut_416_EXMPLR ;
   dataOut(415) <= dataOut_415_EXMPLR ;
   dataOut(414) <= dataOut_414_EXMPLR ;
   dataOut(413) <= dataOut_413_EXMPLR ;
   dataOut(412) <= dataOut_412_EXMPLR ;
   dataOut(411) <= dataOut_411_EXMPLR ;
   dataOut(410) <= dataOut_410_EXMPLR ;
   dataOut(409) <= dataOut_409_EXMPLR ;
   dataOut(408) <= dataOut_408_EXMPLR ;
   dataOut(407) <= dataOut_407_EXMPLR ;
   dataOut(406) <= dataOut_406_EXMPLR ;
   dataOut(405) <= dataOut_405_EXMPLR ;
   dataOut(404) <= dataOut_404_EXMPLR ;
   dataOut(403) <= dataOut_403_EXMPLR ;
   dataOut(402) <= dataOut_402_EXMPLR ;
   dataOut(401) <= dataOut_401_EXMPLR ;
   dataOut(400) <= dataOut_400_EXMPLR ;
   dataOut(399) <= dataOut_399_EXMPLR ;
   dataOut(398) <= dataOut_398_EXMPLR ;
   dataOut(397) <= dataOut_397_EXMPLR ;
   dataOut(396) <= dataOut_396_EXMPLR ;
   dataOut(395) <= dataOut_395_EXMPLR ;
   dataOut(394) <= dataOut_394_EXMPLR ;
   dataOut(393) <= dataOut_393_EXMPLR ;
   dataOut(392) <= dataOut_392_EXMPLR ;
   dataOut(391) <= dataOut_391_EXMPLR ;
   dataOut(390) <= dataOut_390_EXMPLR ;
   dataOut(389) <= dataOut_389_EXMPLR ;
   dataOut(388) <= dataOut_388_EXMPLR ;
   dataOut(387) <= dataOut_387_EXMPLR ;
   dataOut(386) <= dataOut_386_EXMPLR ;
   dataOut(385) <= dataOut_385_EXMPLR ;
   dataOut(384) <= dataOut_384_EXMPLR ;
   dataOut(383) <= dataOut_383_EXMPLR ;
   dataOut(382) <= dataOut_382_EXMPLR ;
   dataOut(381) <= dataOut_381_EXMPLR ;
   dataOut(380) <= dataOut_380_EXMPLR ;
   dataOut(379) <= dataOut_379_EXMPLR ;
   dataOut(378) <= dataOut_378_EXMPLR ;
   dataOut(377) <= dataOut_377_EXMPLR ;
   dataOut(376) <= dataOut_376_EXMPLR ;
   dataOut(375) <= dataOut_375_EXMPLR ;
   dataOut(374) <= dataOut_374_EXMPLR ;
   dataOut(373) <= dataOut_373_EXMPLR ;
   dataOut(372) <= dataOut_372_EXMPLR ;
   dataOut(371) <= dataOut_371_EXMPLR ;
   dataOut(370) <= dataOut_370_EXMPLR ;
   dataOut(369) <= dataOut_369_EXMPLR ;
   dataOut(368) <= dataOut_368_EXMPLR ;
   dataOut(367) <= dataOut_367_EXMPLR ;
   dataOut(366) <= dataOut_366_EXMPLR ;
   dataOut(365) <= dataOut_365_EXMPLR ;
   dataOut(364) <= dataOut_364_EXMPLR ;
   dataOut(363) <= dataOut_363_EXMPLR ;
   dataOut(362) <= dataOut_362_EXMPLR ;
   dataOut(361) <= dataOut_361_EXMPLR ;
   dataOut(360) <= dataOut_360_EXMPLR ;
   dataOut(359) <= dataOut_359_EXMPLR ;
   dataOut(358) <= dataOut_358_EXMPLR ;
   dataOut(357) <= dataOut_357_EXMPLR ;
   dataOut(356) <= dataOut_356_EXMPLR ;
   dataOut(355) <= dataOut_355_EXMPLR ;
   dataOut(354) <= dataOut_354_EXMPLR ;
   dataOut(353) <= dataOut_353_EXMPLR ;
   dataOut(352) <= dataOut_352_EXMPLR ;
   dataOut(351) <= dataOut_351_EXMPLR ;
   dataOut(350) <= dataOut_350_EXMPLR ;
   dataOut(349) <= dataOut_349_EXMPLR ;
   dataOut(348) <= dataOut_348_EXMPLR ;
   dataOut(347) <= dataOut_347_EXMPLR ;
   dataOut(346) <= dataOut_346_EXMPLR ;
   dataOut(345) <= dataOut_345_EXMPLR ;
   dataOut(344) <= dataOut_344_EXMPLR ;
   dataOut(343) <= dataOut_343_EXMPLR ;
   dataOut(342) <= dataOut_342_EXMPLR ;
   dataOut(341) <= dataOut_341_EXMPLR ;
   dataOut(340) <= dataOut_340_EXMPLR ;
   dataOut(339) <= dataOut_339_EXMPLR ;
   dataOut(338) <= dataOut_338_EXMPLR ;
   dataOut(337) <= dataOut_337_EXMPLR ;
   dataOut(336) <= dataOut_336_EXMPLR ;
   dataOut(335) <= dataOut_335_EXMPLR ;
   dataOut(334) <= dataOut_334_EXMPLR ;
   dataOut(333) <= dataOut_333_EXMPLR ;
   dataOut(332) <= dataOut_332_EXMPLR ;
   dataOut(331) <= dataOut_331_EXMPLR ;
   dataOut(330) <= dataOut_330_EXMPLR ;
   dataOut(329) <= dataOut_329_EXMPLR ;
   dataOut(328) <= dataOut_328_EXMPLR ;
   dataOut(327) <= dataOut_327_EXMPLR ;
   dataOut(326) <= dataOut_326_EXMPLR ;
   dataOut(325) <= dataOut_325_EXMPLR ;
   dataOut(324) <= dataOut_324_EXMPLR ;
   dataOut(323) <= dataOut_323_EXMPLR ;
   dataOut(322) <= dataOut_322_EXMPLR ;
   dataOut(321) <= dataOut_321_EXMPLR ;
   dataOut(320) <= dataOut_320_EXMPLR ;
   dataOut(319) <= dataOut_319_EXMPLR ;
   dataOut(318) <= dataOut_318_EXMPLR ;
   dataOut(317) <= dataOut_317_EXMPLR ;
   dataOut(316) <= dataOut_316_EXMPLR ;
   dataOut(315) <= dataOut_315_EXMPLR ;
   dataOut(314) <= dataOut_314_EXMPLR ;
   dataOut(313) <= dataOut_313_EXMPLR ;
   dataOut(312) <= dataOut_312_EXMPLR ;
   dataOut(311) <= dataOut_311_EXMPLR ;
   dataOut(310) <= dataOut_310_EXMPLR ;
   dataOut(309) <= dataOut_309_EXMPLR ;
   dataOut(308) <= dataOut_308_EXMPLR ;
   dataOut(307) <= dataOut_307_EXMPLR ;
   dataOut(306) <= dataOut_306_EXMPLR ;
   dataOut(305) <= dataOut_305_EXMPLR ;
   dataOut(304) <= dataOut_304_EXMPLR ;
   dataOut(303) <= dataOut_303_EXMPLR ;
   dataOut(302) <= dataOut_302_EXMPLR ;
   dataOut(301) <= dataOut_301_EXMPLR ;
   dataOut(300) <= dataOut_300_EXMPLR ;
   dataOut(299) <= dataOut_299_EXMPLR ;
   dataOut(298) <= dataOut_298_EXMPLR ;
   dataOut(297) <= dataOut_297_EXMPLR ;
   dataOut(296) <= dataOut_296_EXMPLR ;
   dataOut(295) <= dataOut_295_EXMPLR ;
   dataOut(294) <= dataOut_294_EXMPLR ;
   dataOut(293) <= dataOut_293_EXMPLR ;
   dataOut(292) <= dataOut_292_EXMPLR ;
   dataOut(291) <= dataOut_291_EXMPLR ;
   dataOut(290) <= dataOut_290_EXMPLR ;
   dataOut(289) <= dataOut_289_EXMPLR ;
   dataOut(288) <= dataOut_288_EXMPLR ;
   dataOut(287) <= dataOut_287_EXMPLR ;
   dataOut(286) <= dataOut_286_EXMPLR ;
   dataOut(285) <= dataOut_285_EXMPLR ;
   dataOut(284) <= dataOut_284_EXMPLR ;
   dataOut(283) <= dataOut_283_EXMPLR ;
   dataOut(282) <= dataOut_282_EXMPLR ;
   dataOut(281) <= dataOut_281_EXMPLR ;
   dataOut(280) <= dataOut_280_EXMPLR ;
   dataOut(279) <= dataOut_279_EXMPLR ;
   dataOut(278) <= dataOut_278_EXMPLR ;
   dataOut(277) <= dataOut_277_EXMPLR ;
   dataOut(276) <= dataOut_276_EXMPLR ;
   dataOut(275) <= dataOut_275_EXMPLR ;
   dataOut(274) <= dataOut_274_EXMPLR ;
   dataOut(273) <= dataOut_273_EXMPLR ;
   dataOut(272) <= dataOut_272_EXMPLR ;
   dataOut(271) <= dataOut_271_EXMPLR ;
   dataOut(270) <= dataOut_270_EXMPLR ;
   dataOut(269) <= dataOut_269_EXMPLR ;
   dataOut(268) <= dataOut_268_EXMPLR ;
   dataOut(267) <= dataOut_267_EXMPLR ;
   dataOut(266) <= dataOut_266_EXMPLR ;
   dataOut(265) <= dataOut_265_EXMPLR ;
   dataOut(264) <= dataOut_264_EXMPLR ;
   dataOut(263) <= dataOut_263_EXMPLR ;
   dataOut(262) <= dataOut_262_EXMPLR ;
   dataOut(261) <= dataOut_261_EXMPLR ;
   dataOut(260) <= dataOut_260_EXMPLR ;
   dataOut(259) <= dataOut_259_EXMPLR ;
   dataOut(258) <= dataOut_258_EXMPLR ;
   dataOut(257) <= dataOut_257_EXMPLR ;
   dataOut(256) <= dataOut_256_EXMPLR ;
   dataOut(255) <= dataOut_255_EXMPLR ;
   dataOut(254) <= dataOut_254_EXMPLR ;
   dataOut(253) <= dataOut_253_EXMPLR ;
   dataOut(252) <= dataOut_252_EXMPLR ;
   dataOut(251) <= dataOut_251_EXMPLR ;
   dataOut(250) <= dataOut_250_EXMPLR ;
   dataOut(249) <= dataOut_249_EXMPLR ;
   dataOut(248) <= dataOut_248_EXMPLR ;
   dataOut(247) <= dataOut_247_EXMPLR ;
   dataOut(246) <= dataOut_246_EXMPLR ;
   dataOut(245) <= dataOut_245_EXMPLR ;
   dataOut(244) <= dataOut_244_EXMPLR ;
   dataOut(243) <= dataOut_243_EXMPLR ;
   dataOut(242) <= dataOut_242_EXMPLR ;
   dataOut(241) <= dataOut_241_EXMPLR ;
   dataOut(240) <= dataOut_240_EXMPLR ;
   dataOut(239) <= dataOut_239_EXMPLR ;
   dataOut(238) <= dataOut_238_EXMPLR ;
   dataOut(237) <= dataOut_237_EXMPLR ;
   dataOut(236) <= dataOut_236_EXMPLR ;
   dataOut(235) <= dataOut_235_EXMPLR ;
   dataOut(234) <= dataOut_234_EXMPLR ;
   dataOut(233) <= dataOut_233_EXMPLR ;
   dataOut(232) <= dataOut_232_EXMPLR ;
   dataOut(231) <= dataOut_231_EXMPLR ;
   dataOut(230) <= dataOut_230_EXMPLR ;
   dataOut(229) <= dataOut_229_EXMPLR ;
   dataOut(228) <= dataOut_228_EXMPLR ;
   dataOut(227) <= dataOut_227_EXMPLR ;
   dataOut(226) <= dataOut_226_EXMPLR ;
   dataOut(225) <= dataOut_225_EXMPLR ;
   dataOut(224) <= dataOut_224_EXMPLR ;
   dataOut(223) <= dataOut_223_EXMPLR ;
   dataOut(222) <= dataOut_222_EXMPLR ;
   dataOut(221) <= dataOut_221_EXMPLR ;
   dataOut(220) <= dataOut_220_EXMPLR ;
   dataOut(219) <= dataOut_219_EXMPLR ;
   dataOut(218) <= dataOut_218_EXMPLR ;
   dataOut(217) <= dataOut_217_EXMPLR ;
   dataOut(216) <= dataOut_216_EXMPLR ;
   dataOut(215) <= dataOut_215_EXMPLR ;
   dataOut(214) <= dataOut_214_EXMPLR ;
   dataOut(213) <= dataOut_213_EXMPLR ;
   dataOut(212) <= dataOut_212_EXMPLR ;
   dataOut(211) <= dataOut_211_EXMPLR ;
   dataOut(210) <= dataOut_210_EXMPLR ;
   dataOut(209) <= dataOut_209_EXMPLR ;
   dataOut(208) <= dataOut_208_EXMPLR ;
   dataOut(207) <= dataOut_207_EXMPLR ;
   dataOut(206) <= dataOut_206_EXMPLR ;
   dataOut(205) <= dataOut_205_EXMPLR ;
   dataOut(204) <= dataOut_204_EXMPLR ;
   dataOut(203) <= dataOut_203_EXMPLR ;
   dataOut(202) <= dataOut_202_EXMPLR ;
   dataOut(201) <= dataOut_201_EXMPLR ;
   dataOut(200) <= dataOut_200_EXMPLR ;
   dataOut(199) <= dataOut_199_EXMPLR ;
   dataOut(198) <= dataOut_198_EXMPLR ;
   dataOut(197) <= dataOut_197_EXMPLR ;
   dataOut(196) <= dataOut_196_EXMPLR ;
   dataOut(195) <= dataOut_195_EXMPLR ;
   dataOut(194) <= dataOut_194_EXMPLR ;
   dataOut(193) <= dataOut_193_EXMPLR ;
   dataOut(192) <= dataOut_192_EXMPLR ;
   dataOut(191) <= dataOut_191_EXMPLR ;
   dataOut(190) <= dataOut_190_EXMPLR ;
   dataOut(189) <= dataOut_189_EXMPLR ;
   dataOut(188) <= dataOut_188_EXMPLR ;
   dataOut(187) <= dataOut_187_EXMPLR ;
   dataOut(186) <= dataOut_186_EXMPLR ;
   dataOut(185) <= dataOut_185_EXMPLR ;
   dataOut(184) <= dataOut_184_EXMPLR ;
   dataOut(183) <= dataOut_183_EXMPLR ;
   dataOut(182) <= dataOut_182_EXMPLR ;
   dataOut(181) <= dataOut_181_EXMPLR ;
   dataOut(180) <= dataOut_180_EXMPLR ;
   dataOut(179) <= dataOut_179_EXMPLR ;
   dataOut(178) <= dataOut_178_EXMPLR ;
   dataOut(177) <= dataOut_177_EXMPLR ;
   dataOut(176) <= dataOut_176_EXMPLR ;
   dataOut(175) <= dataOut_175_EXMPLR ;
   dataOut(174) <= dataOut_174_EXMPLR ;
   dataOut(173) <= dataOut_173_EXMPLR ;
   dataOut(172) <= dataOut_172_EXMPLR ;
   dataOut(171) <= dataOut_171_EXMPLR ;
   dataOut(170) <= dataOut_170_EXMPLR ;
   dataOut(169) <= dataOut_169_EXMPLR ;
   dataOut(168) <= dataOut_168_EXMPLR ;
   dataOut(167) <= dataOut_167_EXMPLR ;
   dataOut(166) <= dataOut_166_EXMPLR ;
   dataOut(165) <= dataOut_165_EXMPLR ;
   dataOut(164) <= dataOut_164_EXMPLR ;
   dataOut(163) <= dataOut_163_EXMPLR ;
   dataOut(162) <= dataOut_162_EXMPLR ;
   dataOut(161) <= dataOut_161_EXMPLR ;
   dataOut(160) <= dataOut_160_EXMPLR ;
   dataOut(159) <= dataOut_159_EXMPLR ;
   dataOut(158) <= dataOut_158_EXMPLR ;
   dataOut(157) <= dataOut_157_EXMPLR ;
   dataOut(156) <= dataOut_156_EXMPLR ;
   dataOut(155) <= dataOut_155_EXMPLR ;
   dataOut(154) <= dataOut_154_EXMPLR ;
   dataOut(153) <= dataOut_153_EXMPLR ;
   dataOut(152) <= dataOut_152_EXMPLR ;
   dataOut(151) <= dataOut_151_EXMPLR ;
   dataOut(150) <= dataOut_150_EXMPLR ;
   dataOut(149) <= dataOut_149_EXMPLR ;
   dataOut(148) <= dataOut_148_EXMPLR ;
   dataOut(147) <= dataOut_147_EXMPLR ;
   dataOut(146) <= dataOut_146_EXMPLR ;
   dataOut(145) <= dataOut_145_EXMPLR ;
   dataOut(144) <= dataOut_144_EXMPLR ;
   dataOut(143) <= dataOut_143_EXMPLR ;
   dataOut(142) <= dataOut_142_EXMPLR ;
   dataOut(141) <= dataOut_141_EXMPLR ;
   dataOut(140) <= dataOut_140_EXMPLR ;
   dataOut(139) <= dataOut_139_EXMPLR ;
   dataOut(138) <= dataOut_138_EXMPLR ;
   dataOut(137) <= dataOut_137_EXMPLR ;
   dataOut(136) <= dataOut_136_EXMPLR ;
   dataOut(135) <= dataOut_135_EXMPLR ;
   dataOut(134) <= dataOut_134_EXMPLR ;
   dataOut(133) <= dataOut_133_EXMPLR ;
   dataOut(132) <= dataOut_132_EXMPLR ;
   dataOut(131) <= dataOut_131_EXMPLR ;
   dataOut(130) <= dataOut_130_EXMPLR ;
   dataOut(129) <= dataOut_129_EXMPLR ;
   dataOut(128) <= dataOut_128_EXMPLR ;
   dataOut(127) <= dataOut_127_EXMPLR ;
   dataOut(126) <= dataOut_126_EXMPLR ;
   dataOut(125) <= dataOut_125_EXMPLR ;
   dataOut(124) <= dataOut_124_EXMPLR ;
   dataOut(123) <= dataOut_123_EXMPLR ;
   dataOut(122) <= dataOut_122_EXMPLR ;
   dataOut(121) <= dataOut_121_EXMPLR ;
   dataOut(120) <= dataOut_120_EXMPLR ;
   dataOut(119) <= dataOut_119_EXMPLR ;
   dataOut(118) <= dataOut_118_EXMPLR ;
   dataOut(117) <= dataOut_117_EXMPLR ;
   dataOut(116) <= dataOut_116_EXMPLR ;
   dataOut(115) <= dataOut_115_EXMPLR ;
   dataOut(114) <= dataOut_114_EXMPLR ;
   dataOut(113) <= dataOut_113_EXMPLR ;
   dataOut(112) <= dataOut_112_EXMPLR ;
   dataOut(111) <= dataOut_111_EXMPLR ;
   dataOut(110) <= dataOut_110_EXMPLR ;
   dataOut(109) <= dataOut_109_EXMPLR ;
   dataOut(108) <= dataOut_108_EXMPLR ;
   dataOut(107) <= dataOut_107_EXMPLR ;
   dataOut(106) <= dataOut_106_EXMPLR ;
   dataOut(105) <= dataOut_105_EXMPLR ;
   dataOut(104) <= dataOut_104_EXMPLR ;
   dataOut(103) <= dataOut_103_EXMPLR ;
   dataOut(102) <= dataOut_102_EXMPLR ;
   dataOut(101) <= dataOut_101_EXMPLR ;
   dataOut(100) <= dataOut_100_EXMPLR ;
   dataOut(99) <= dataOut_99_EXMPLR ;
   dataOut(98) <= dataOut_98_EXMPLR ;
   dataOut(97) <= dataOut_97_EXMPLR ;
   dataOut(96) <= dataOut_96_EXMPLR ;
   dataOut(95) <= dataOut_95_EXMPLR ;
   dataOut(94) <= dataOut_94_EXMPLR ;
   dataOut(93) <= dataOut_93_EXMPLR ;
   dataOut(92) <= dataOut_92_EXMPLR ;
   dataOut(91) <= dataOut_91_EXMPLR ;
   dataOut(90) <= dataOut_90_EXMPLR ;
   dataOut(89) <= dataOut_89_EXMPLR ;
   dataOut(88) <= dataOut_88_EXMPLR ;
   dataOut(87) <= dataOut_87_EXMPLR ;
   dataOut(86) <= dataOut_86_EXMPLR ;
   dataOut(85) <= dataOut_85_EXMPLR ;
   dataOut(84) <= dataOut_84_EXMPLR ;
   dataOut(83) <= dataOut_83_EXMPLR ;
   dataOut(82) <= dataOut_82_EXMPLR ;
   dataOut(81) <= dataOut_81_EXMPLR ;
   dataOut(80) <= dataOut_80_EXMPLR ;
   dataOut(79) <= dataOut_79_EXMPLR ;
   dataOut(78) <= dataOut_78_EXMPLR ;
   dataOut(77) <= dataOut_77_EXMPLR ;
   dataOut(76) <= dataOut_76_EXMPLR ;
   dataOut(75) <= dataOut_75_EXMPLR ;
   dataOut(74) <= dataOut_74_EXMPLR ;
   dataOut(73) <= dataOut_73_EXMPLR ;
   dataOut(72) <= dataOut_72_EXMPLR ;
   dataOut(71) <= dataOut_71_EXMPLR ;
   dataOut(70) <= dataOut_70_EXMPLR ;
   dataOut(69) <= dataOut_69_EXMPLR ;
   dataOut(68) <= dataOut_68_EXMPLR ;
   dataOut(67) <= dataOut_67_EXMPLR ;
   dataOut(66) <= dataOut_66_EXMPLR ;
   dataOut(65) <= dataOut_65_EXMPLR ;
   dataOut(64) <= dataOut_64_EXMPLR ;
   dataOut(63) <= dataOut_63_EXMPLR ;
   dataOut(62) <= dataOut_62_EXMPLR ;
   dataOut(61) <= dataOut_61_EXMPLR ;
   dataOut(60) <= dataOut_60_EXMPLR ;
   dataOut(59) <= dataOut_59_EXMPLR ;
   dataOut(58) <= dataOut_58_EXMPLR ;
   dataOut(57) <= dataOut_57_EXMPLR ;
   dataOut(56) <= dataOut_56_EXMPLR ;
   dataOut(55) <= dataOut_55_EXMPLR ;
   dataOut(54) <= dataOut_54_EXMPLR ;
   dataOut(53) <= dataOut_53_EXMPLR ;
   dataOut(52) <= dataOut_52_EXMPLR ;
   dataOut(51) <= dataOut_51_EXMPLR ;
   dataOut(50) <= dataOut_50_EXMPLR ;
   dataOut(49) <= dataOut_49_EXMPLR ;
   dataOut(48) <= dataOut_48_EXMPLR ;
   dataOut(47) <= dataOut_47_EXMPLR ;
   dataOut(46) <= dataOut_46_EXMPLR ;
   dataOut(45) <= dataOut_45_EXMPLR ;
   dataOut(44) <= dataOut_44_EXMPLR ;
   dataOut(43) <= dataOut_43_EXMPLR ;
   dataOut(42) <= dataOut_42_EXMPLR ;
   dataOut(41) <= dataOut_41_EXMPLR ;
   dataOut(40) <= dataOut_40_EXMPLR ;
   dataOut(39) <= dataOut_39_EXMPLR ;
   dataOut(38) <= dataOut_38_EXMPLR ;
   dataOut(37) <= dataOut_37_EXMPLR ;
   dataOut(36) <= dataOut_36_EXMPLR ;
   dataOut(35) <= dataOut_35_EXMPLR ;
   dataOut(34) <= dataOut_34_EXMPLR ;
   dataOut(33) <= dataOut_33_EXMPLR ;
   dataOut(32) <= dataOut_32_EXMPLR ;
   dataOut(31) <= dataOut_31_EXMPLR ;
   dataOut(30) <= dataOut_30_EXMPLR ;
   dataOut(29) <= dataOut_29_EXMPLR ;
   dataOut(28) <= dataOut_28_EXMPLR ;
   dataOut(27) <= dataOut_27_EXMPLR ;
   dataOut(26) <= dataOut_26_EXMPLR ;
   dataOut(25) <= dataOut_25_EXMPLR ;
   dataOut(24) <= dataOut_24_EXMPLR ;
   dataOut(23) <= dataOut_23_EXMPLR ;
   dataOut(22) <= dataOut_22_EXMPLR ;
   dataOut(21) <= dataOut_21_EXMPLR ;
   dataOut(20) <= dataOut_20_EXMPLR ;
   dataOut(19) <= dataOut_19_EXMPLR ;
   dataOut(18) <= dataOut_18_EXMPLR ;
   dataOut(17) <= dataOut_17_EXMPLR ;
   dataOut(16) <= dataOut_16_EXMPLR ;
   dataOut(15) <= dataOut_15_EXMPLR ;
   dataOut(14) <= dataOut_14_EXMPLR ;
   dataOut(13) <= dataOut_13_EXMPLR ;
   dataOut(12) <= dataOut_12_EXMPLR ;
   dataOut(11) <= dataOut_11_EXMPLR ;
   dataOut(10) <= dataOut_10_EXMPLR ;
   dataOut(9) <= dataOut_9_EXMPLR ;
   dataOut(8) <= dataOut_8_EXMPLR ;
   dataOut(7) <= dataOut_7_EXMPLR ;
   dataOut(6) <= dataOut_6_EXMPLR ;
   dataOut(5) <= dataOut_5_EXMPLR ;
   dataOut(4) <= dataOut_4_EXMPLR ;
   dataOut(3) <= dataOut_3_EXMPLR ;
   dataOut(2) <= dataOut_2_EXMPLR ;
   dataOut(1) <= dataOut_1_EXMPLR ;
   dataOut(0) <= dataOut_0_EXMPLR ;
   Ram1Rd : triStateBuffer_448 port map ( D(447)=>nx5655, D(446)=>nx5655, 
      D(445)=>nx5655, D(444)=>nx5655, D(443)=>nx5655, D(442)=>nx5655, D(441)
      =>nx5655, D(440)=>nx5657, D(439)=>nx5657, D(438)=>nx5657, D(437)=>
      nx5657, D(436)=>nx5657, D(435)=>nx5657, D(434)=>nx5657, D(433)=>nx5659, 
      D(432)=>nx5659, D(431)=>nx5659, D(430)=>nx5659, D(429)=>nx5659, D(428)
      =>nx5659, D(427)=>nx5659, D(426)=>nx5661, D(425)=>nx5661, D(424)=>
      nx5661, D(423)=>nx5661, D(422)=>nx5661, D(421)=>nx5661, D(420)=>nx5661, 
      D(419)=>nx5663, D(418)=>nx5663, D(417)=>nx5663, D(416)=>nx5663, D(415)
      =>nx5663, D(414)=>nx5663, D(413)=>nx5663, D(412)=>nx5665, D(411)=>
      nx5665, D(410)=>nx5665, D(409)=>nx5665, D(408)=>nx5665, D(407)=>nx5665, 
      D(406)=>nx5665, D(405)=>nx5667, D(404)=>nx5667, D(403)=>nx5667, D(402)
      =>nx5667, D(401)=>nx5667, D(400)=>nx5667, D(399)=>nx5667, D(398)=>
      nx5669, D(397)=>nx5669, D(396)=>nx5669, D(395)=>nx5669, D(394)=>nx5669, 
      D(393)=>nx5669, D(392)=>nx5669, D(391)=>nx5671, D(390)=>nx5671, D(389)
      =>nx5671, D(388)=>nx5671, D(387)=>nx5671, D(386)=>nx5671, D(385)=>
      nx5671, D(384)=>nx5673, D(383)=>nx5673, D(382)=>nx5673, D(381)=>nx5673, 
      D(380)=>nx5673, D(379)=>nx5673, D(378)=>nx5673, D(377)=>nx5675, D(376)
      =>nx5675, D(375)=>nx5675, D(374)=>nx5675, D(373)=>nx5675, D(372)=>
      nx5675, D(371)=>nx5675, D(370)=>nx5677, D(369)=>nx5677, D(368)=>nx5677, 
      D(367)=>nx5677, D(366)=>nx5677, D(365)=>nx5677, D(364)=>nx5677, D(363)
      =>nx5679, D(362)=>nx5679, D(361)=>nx5679, D(360)=>nx5679, D(359)=>
      nx5679, D(358)=>nx5679, D(357)=>nx5679, D(356)=>nx5681, D(355)=>nx5681, 
      D(354)=>nx5681, D(353)=>nx5681, D(352)=>nx5681, D(351)=>nx5681, D(350)
      =>nx5681, D(349)=>nx5683, D(348)=>nx5683, D(347)=>nx5683, D(346)=>
      nx5683, D(345)=>nx5683, D(344)=>nx5683, D(343)=>nx5683, D(342)=>nx5685, 
      D(341)=>nx5685, D(340)=>nx5685, D(339)=>nx5685, D(338)=>nx5685, D(337)
      =>nx5685, D(336)=>nx5685, D(335)=>nx5687, D(334)=>nx5687, D(333)=>
      nx5687, D(332)=>nx5687, D(331)=>nx5687, D(330)=>nx5687, D(329)=>nx5687, 
      D(328)=>nx5689, D(327)=>nx5689, D(326)=>nx5689, D(325)=>nx5689, D(324)
      =>nx5689, D(323)=>nx5689, D(322)=>nx5689, D(321)=>nx5691, D(320)=>
      nx5691, D(319)=>nx5691, D(318)=>nx5691, D(317)=>nx5691, D(316)=>nx5691, 
      D(315)=>nx5691, D(314)=>nx5693, D(313)=>nx5693, D(312)=>nx5693, D(311)
      =>nx5693, D(310)=>nx5693, D(309)=>nx5693, D(308)=>nx5693, D(307)=>
      nx5695, D(306)=>nx5695, D(305)=>nx5695, D(304)=>nx5695, D(303)=>nx5695, 
      D(302)=>nx5695, D(301)=>nx5695, D(300)=>nx5697, D(299)=>nx5697, D(298)
      =>nx5697, D(297)=>nx5697, D(296)=>nx5697, D(295)=>nx5697, D(294)=>
      nx5697, D(293)=>nx5699, D(292)=>nx5699, D(291)=>nx5699, D(290)=>nx5699, 
      D(289)=>nx5699, D(288)=>nx5699, D(287)=>nx5699, D(286)=>nx5701, D(285)
      =>nx5701, D(284)=>nx5701, D(283)=>nx5701, D(282)=>nx5701, D(281)=>
      nx5701, D(280)=>nx5701, D(279)=>nx5703, D(278)=>nx5703, D(277)=>nx5703, 
      D(276)=>nx5703, D(275)=>nx5703, D(274)=>nx5703, D(273)=>nx5703, D(272)
      =>nx5705, D(271)=>nx5705, D(270)=>nx5705, D(269)=>nx5705, D(268)=>
      nx5705, D(267)=>nx5705, D(266)=>nx5705, D(265)=>nx5707, D(264)=>nx5707, 
      D(263)=>nx5707, D(262)=>nx5707, D(261)=>nx5707, D(260)=>nx5707, D(259)
      =>nx5707, D(258)=>nx5709, D(257)=>nx5709, D(256)=>nx5709, D(255)=>
      nx5709, D(254)=>nx5709, D(253)=>nx5709, D(252)=>nx5709, D(251)=>nx5711, 
      D(250)=>nx5711, D(249)=>nx5711, D(248)=>nx5711, D(247)=>nx5711, D(246)
      =>nx5711, D(245)=>nx5711, D(244)=>nx5713, D(243)=>nx5713, D(242)=>
      nx5713, D(241)=>nx5713, D(240)=>nx5713, D(239)=>nx5713, D(238)=>nx5713, 
      D(237)=>nx5715, D(236)=>nx5715, D(235)=>nx5715, D(234)=>nx5715, D(233)
      =>nx5715, D(232)=>nx5715, D(231)=>nx5715, D(230)=>nx5717, D(229)=>
      nx5717, D(228)=>nx5717, D(227)=>nx5717, D(226)=>nx5717, D(225)=>nx5717, 
      D(224)=>nx5717, D(223)=>nx5719, D(222)=>nx5719, D(221)=>nx5719, D(220)
      =>nx5719, D(219)=>nx5719, D(218)=>nx5719, D(217)=>nx5719, D(216)=>
      nx5721, D(215)=>nx5721, D(214)=>nx5721, D(213)=>nx5721, D(212)=>nx5721, 
      D(211)=>nx5721, D(210)=>nx5721, D(209)=>nx5723, D(208)=>nx5723, D(207)
      =>nx5723, D(206)=>nx5723, D(205)=>nx5723, D(204)=>nx5723, D(203)=>
      nx5723, D(202)=>nx5725, D(201)=>nx5725, D(200)=>nx5725, D(199)=>nx5725, 
      D(198)=>nx5725, D(197)=>nx5725, D(196)=>nx5725, D(195)=>nx5727, D(194)
      =>nx5727, D(193)=>nx5727, D(192)=>nx5727, D(191)=>nx5727, D(190)=>
      nx5727, D(189)=>nx5727, D(188)=>nx5729, D(187)=>nx5729, D(186)=>nx5729, 
      D(185)=>nx5729, D(184)=>nx5729, D(183)=>nx5729, D(182)=>nx5729, D(181)
      =>nx5731, D(180)=>nx5731, D(179)=>nx5731, D(178)=>nx5731, D(177)=>
      nx5731, D(176)=>nx5731, D(175)=>nx5731, D(174)=>nx5733, D(173)=>nx5733, 
      D(172)=>nx5733, D(171)=>nx5733, D(170)=>nx5733, D(169)=>nx5733, D(168)
      =>nx5733, D(167)=>nx5735, D(166)=>nx5735, D(165)=>nx5735, D(164)=>
      nx5735, D(163)=>nx5735, D(162)=>nx5735, D(161)=>nx5735, D(160)=>nx5737, 
      D(159)=>nx5737, D(158)=>nx5737, D(157)=>nx5737, D(156)=>nx5737, D(155)
      =>nx5737, D(154)=>nx5737, D(153)=>nx5739, D(152)=>nx5739, D(151)=>
      nx5739, D(150)=>nx5739, D(149)=>nx5739, D(148)=>nx5739, D(147)=>nx5739, 
      D(146)=>nx5741, D(145)=>nx5741, D(144)=>nx5741, D(143)=>nx5741, D(142)
      =>nx5741, D(141)=>nx5741, D(140)=>nx5741, D(139)=>nx5743, D(138)=>
      nx5743, D(137)=>nx5743, D(136)=>nx5743, D(135)=>nx5743, D(134)=>nx5743, 
      D(133)=>nx5743, D(132)=>nx5745, D(131)=>nx5745, D(130)=>nx5745, D(129)
      =>nx5745, D(128)=>nx5745, D(127)=>nx5745, D(126)=>nx5745, D(125)=>
      nx5747, D(124)=>nx5747, D(123)=>nx5747, D(122)=>nx5747, D(121)=>nx5747, 
      D(120)=>nx5747, D(119)=>nx5747, D(118)=>nx5749, D(117)=>nx5749, D(116)
      =>nx5749, D(115)=>nx5749, D(114)=>nx5749, D(113)=>nx5749, D(112)=>
      nx5749, D(111)=>nx5751, D(110)=>nx5751, D(109)=>nx5751, D(108)=>nx5751, 
      D(107)=>nx5751, D(106)=>nx5751, D(105)=>nx5751, D(104)=>nx5753, D(103)
      =>nx5753, D(102)=>nx5753, D(101)=>nx5753, D(100)=>nx5753, D(99)=>
      nx5753, D(98)=>nx5753, D(97)=>nx5755, D(96)=>nx5755, D(95)=>nx5755, 
      D(94)=>nx5755, D(93)=>nx5755, D(92)=>nx5755, D(91)=>nx5755, D(90)=>
      nx5757, D(89)=>nx5757, D(88)=>nx5757, D(87)=>nx5757, D(86)=>nx5757, 
      D(85)=>nx5757, D(84)=>nx5757, D(83)=>nx5759, D(82)=>nx5759, D(81)=>
      nx5759, D(80)=>nx5759, D(79)=>nx5759, D(78)=>nx5759, D(77)=>nx5759, 
      D(76)=>nx5761, D(75)=>nx5761, D(74)=>nx5761, D(73)=>nx5761, D(72)=>
      nx5761, D(71)=>nx5761, D(70)=>nx5761, D(69)=>nx5763, D(68)=>nx5763, 
      D(67)=>nx5763, D(66)=>nx5763, D(65)=>nx5763, D(64)=>nx5763, D(63)=>
      nx5763, D(62)=>nx5765, D(61)=>nx5765, D(60)=>nx5765, D(59)=>nx5765, 
      D(58)=>nx5765, D(57)=>nx5765, D(56)=>nx5765, D(55)=>nx5767, D(54)=>
      nx5767, D(53)=>nx5767, D(52)=>nx5767, D(51)=>nx5767, D(50)=>nx5767, 
      D(49)=>nx5767, D(48)=>nx5769, D(47)=>nx5769, D(46)=>nx5769, D(45)=>
      nx5769, D(44)=>nx5769, D(43)=>nx5769, D(42)=>nx5769, D(41)=>nx5771, 
      D(40)=>nx5771, D(39)=>nx5771, D(38)=>nx5771, D(37)=>nx5771, D(36)=>
      nx5771, D(35)=>nx5771, D(34)=>nx5773, D(33)=>nx5773, D(32)=>nx5773, 
      D(31)=>nx5773, D(30)=>nx5773, D(29)=>nx5773, D(28)=>nx5773, D(27)=>
      nx5775, D(26)=>nx5775, D(25)=>nx5775, D(24)=>nx5775, D(23)=>nx5775, 
      D(22)=>nx5775, D(21)=>nx5775, D(20)=>nx5777, D(19)=>nx5777, D(18)=>
      nx5777, D(17)=>nx5777, D(16)=>nx5777, D(15)=>nx5777, D(14)=>nx5777, 
      D(13)=>nx5779, D(12)=>nx5779, D(11)=>nx5779, D(10)=>nx5779, D(9)=>
      nx5779, D(8)=>nx5779, D(7)=>nx5779, D(6)=>nx5781, D(5)=>nx5781, D(4)=>
      nx5781, D(3)=>nx5781, D(2)=>nx5781, D(1)=>nx5781, D(0)=>nx5781, EN=>
      test, F(447)=>dataOut_447_EXMPLR, F(446)=>dataOut_446_EXMPLR, F(445)=>
      dataOut_445_EXMPLR, F(444)=>dataOut_444_EXMPLR, F(443)=>
      dataOut_443_EXMPLR, F(442)=>dataOut_442_EXMPLR, F(441)=>
      dataOut_441_EXMPLR, F(440)=>dataOut_440_EXMPLR, F(439)=>
      dataOut_439_EXMPLR, F(438)=>dataOut_438_EXMPLR, F(437)=>
      dataOut_437_EXMPLR, F(436)=>dataOut_436_EXMPLR, F(435)=>
      dataOut_435_EXMPLR, F(434)=>dataOut_434_EXMPLR, F(433)=>
      dataOut_433_EXMPLR, F(432)=>dataOut_432_EXMPLR, F(431)=>
      dataOut_431_EXMPLR, F(430)=>dataOut_430_EXMPLR, F(429)=>
      dataOut_429_EXMPLR, F(428)=>dataOut_428_EXMPLR, F(427)=>
      dataOut_427_EXMPLR, F(426)=>dataOut_426_EXMPLR, F(425)=>
      dataOut_425_EXMPLR, F(424)=>dataOut_424_EXMPLR, F(423)=>
      dataOut_423_EXMPLR, F(422)=>dataOut_422_EXMPLR, F(421)=>
      dataOut_421_EXMPLR, F(420)=>dataOut_420_EXMPLR, F(419)=>
      dataOut_419_EXMPLR, F(418)=>dataOut_418_EXMPLR, F(417)=>
      dataOut_417_EXMPLR, F(416)=>dataOut_416_EXMPLR, F(415)=>
      dataOut_415_EXMPLR, F(414)=>dataOut_414_EXMPLR, F(413)=>
      dataOut_413_EXMPLR, F(412)=>dataOut_412_EXMPLR, F(411)=>
      dataOut_411_EXMPLR, F(410)=>dataOut_410_EXMPLR, F(409)=>
      dataOut_409_EXMPLR, F(408)=>dataOut_408_EXMPLR, F(407)=>
      dataOut_407_EXMPLR, F(406)=>dataOut_406_EXMPLR, F(405)=>
      dataOut_405_EXMPLR, F(404)=>dataOut_404_EXMPLR, F(403)=>
      dataOut_403_EXMPLR, F(402)=>dataOut_402_EXMPLR, F(401)=>
      dataOut_401_EXMPLR, F(400)=>dataOut_400_EXMPLR, F(399)=>
      dataOut_399_EXMPLR, F(398)=>dataOut_398_EXMPLR, F(397)=>
      dataOut_397_EXMPLR, F(396)=>dataOut_396_EXMPLR, F(395)=>
      dataOut_395_EXMPLR, F(394)=>dataOut_394_EXMPLR, F(393)=>
      dataOut_393_EXMPLR, F(392)=>dataOut_392_EXMPLR, F(391)=>
      dataOut_391_EXMPLR, F(390)=>dataOut_390_EXMPLR, F(389)=>
      dataOut_389_EXMPLR, F(388)=>dataOut_388_EXMPLR, F(387)=>
      dataOut_387_EXMPLR, F(386)=>dataOut_386_EXMPLR, F(385)=>
      dataOut_385_EXMPLR, F(384)=>dataOut_384_EXMPLR, F(383)=>
      dataOut_383_EXMPLR, F(382)=>dataOut_382_EXMPLR, F(381)=>
      dataOut_381_EXMPLR, F(380)=>dataOut_380_EXMPLR, F(379)=>
      dataOut_379_EXMPLR, F(378)=>dataOut_378_EXMPLR, F(377)=>
      dataOut_377_EXMPLR, F(376)=>dataOut_376_EXMPLR, F(375)=>
      dataOut_375_EXMPLR, F(374)=>dataOut_374_EXMPLR, F(373)=>
      dataOut_373_EXMPLR, F(372)=>dataOut_372_EXMPLR, F(371)=>
      dataOut_371_EXMPLR, F(370)=>dataOut_370_EXMPLR, F(369)=>
      dataOut_369_EXMPLR, F(368)=>dataOut_368_EXMPLR, F(367)=>
      dataOut_367_EXMPLR, F(366)=>dataOut_366_EXMPLR, F(365)=>
      dataOut_365_EXMPLR, F(364)=>dataOut_364_EXMPLR, F(363)=>
      dataOut_363_EXMPLR, F(362)=>dataOut_362_EXMPLR, F(361)=>
      dataOut_361_EXMPLR, F(360)=>dataOut_360_EXMPLR, F(359)=>
      dataOut_359_EXMPLR, F(358)=>dataOut_358_EXMPLR, F(357)=>
      dataOut_357_EXMPLR, F(356)=>dataOut_356_EXMPLR, F(355)=>
      dataOut_355_EXMPLR, F(354)=>dataOut_354_EXMPLR, F(353)=>
      dataOut_353_EXMPLR, F(352)=>dataOut_352_EXMPLR, F(351)=>
      dataOut_351_EXMPLR, F(350)=>dataOut_350_EXMPLR, F(349)=>
      dataOut_349_EXMPLR, F(348)=>dataOut_348_EXMPLR, F(347)=>
      dataOut_347_EXMPLR, F(346)=>dataOut_346_EXMPLR, F(345)=>
      dataOut_345_EXMPLR, F(344)=>dataOut_344_EXMPLR, F(343)=>
      dataOut_343_EXMPLR, F(342)=>dataOut_342_EXMPLR, F(341)=>
      dataOut_341_EXMPLR, F(340)=>dataOut_340_EXMPLR, F(339)=>
      dataOut_339_EXMPLR, F(338)=>dataOut_338_EXMPLR, F(337)=>
      dataOut_337_EXMPLR, F(336)=>dataOut_336_EXMPLR, F(335)=>
      dataOut_335_EXMPLR, F(334)=>dataOut_334_EXMPLR, F(333)=>
      dataOut_333_EXMPLR, F(332)=>dataOut_332_EXMPLR, F(331)=>
      dataOut_331_EXMPLR, F(330)=>dataOut_330_EXMPLR, F(329)=>
      dataOut_329_EXMPLR, F(328)=>dataOut_328_EXMPLR, F(327)=>
      dataOut_327_EXMPLR, F(326)=>dataOut_326_EXMPLR, F(325)=>
      dataOut_325_EXMPLR, F(324)=>dataOut_324_EXMPLR, F(323)=>
      dataOut_323_EXMPLR, F(322)=>dataOut_322_EXMPLR, F(321)=>
      dataOut_321_EXMPLR, F(320)=>dataOut_320_EXMPLR, F(319)=>
      dataOut_319_EXMPLR, F(318)=>dataOut_318_EXMPLR, F(317)=>
      dataOut_317_EXMPLR, F(316)=>dataOut_316_EXMPLR, F(315)=>
      dataOut_315_EXMPLR, F(314)=>dataOut_314_EXMPLR, F(313)=>
      dataOut_313_EXMPLR, F(312)=>dataOut_312_EXMPLR, F(311)=>
      dataOut_311_EXMPLR, F(310)=>dataOut_310_EXMPLR, F(309)=>
      dataOut_309_EXMPLR, F(308)=>dataOut_308_EXMPLR, F(307)=>
      dataOut_307_EXMPLR, F(306)=>dataOut_306_EXMPLR, F(305)=>
      dataOut_305_EXMPLR, F(304)=>dataOut_304_EXMPLR, F(303)=>
      dataOut_303_EXMPLR, F(302)=>dataOut_302_EXMPLR, F(301)=>
      dataOut_301_EXMPLR, F(300)=>dataOut_300_EXMPLR, F(299)=>
      dataOut_299_EXMPLR, F(298)=>dataOut_298_EXMPLR, F(297)=>
      dataOut_297_EXMPLR, F(296)=>dataOut_296_EXMPLR, F(295)=>
      dataOut_295_EXMPLR, F(294)=>dataOut_294_EXMPLR, F(293)=>
      dataOut_293_EXMPLR, F(292)=>dataOut_292_EXMPLR, F(291)=>
      dataOut_291_EXMPLR, F(290)=>dataOut_290_EXMPLR, F(289)=>
      dataOut_289_EXMPLR, F(288)=>dataOut_288_EXMPLR, F(287)=>
      dataOut_287_EXMPLR, F(286)=>dataOut_286_EXMPLR, F(285)=>
      dataOut_285_EXMPLR, F(284)=>dataOut_284_EXMPLR, F(283)=>
      dataOut_283_EXMPLR, F(282)=>dataOut_282_EXMPLR, F(281)=>
      dataOut_281_EXMPLR, F(280)=>dataOut_280_EXMPLR, F(279)=>
      dataOut_279_EXMPLR, F(278)=>dataOut_278_EXMPLR, F(277)=>
      dataOut_277_EXMPLR, F(276)=>dataOut_276_EXMPLR, F(275)=>
      dataOut_275_EXMPLR, F(274)=>dataOut_274_EXMPLR, F(273)=>
      dataOut_273_EXMPLR, F(272)=>dataOut_272_EXMPLR, F(271)=>
      dataOut_271_EXMPLR, F(270)=>dataOut_270_EXMPLR, F(269)=>
      dataOut_269_EXMPLR, F(268)=>dataOut_268_EXMPLR, F(267)=>
      dataOut_267_EXMPLR, F(266)=>dataOut_266_EXMPLR, F(265)=>
      dataOut_265_EXMPLR, F(264)=>dataOut_264_EXMPLR, F(263)=>
      dataOut_263_EXMPLR, F(262)=>dataOut_262_EXMPLR, F(261)=>
      dataOut_261_EXMPLR, F(260)=>dataOut_260_EXMPLR, F(259)=>
      dataOut_259_EXMPLR, F(258)=>dataOut_258_EXMPLR, F(257)=>
      dataOut_257_EXMPLR, F(256)=>dataOut_256_EXMPLR, F(255)=>
      dataOut_255_EXMPLR, F(254)=>dataOut_254_EXMPLR, F(253)=>
      dataOut_253_EXMPLR, F(252)=>dataOut_252_EXMPLR, F(251)=>
      dataOut_251_EXMPLR, F(250)=>dataOut_250_EXMPLR, F(249)=>
      dataOut_249_EXMPLR, F(248)=>dataOut_248_EXMPLR, F(247)=>
      dataOut_247_EXMPLR, F(246)=>dataOut_246_EXMPLR, F(245)=>
      dataOut_245_EXMPLR, F(244)=>dataOut_244_EXMPLR, F(243)=>
      dataOut_243_EXMPLR, F(242)=>dataOut_242_EXMPLR, F(241)=>
      dataOut_241_EXMPLR, F(240)=>dataOut_240_EXMPLR, F(239)=>
      dataOut_239_EXMPLR, F(238)=>dataOut_238_EXMPLR, F(237)=>
      dataOut_237_EXMPLR, F(236)=>dataOut_236_EXMPLR, F(235)=>
      dataOut_235_EXMPLR, F(234)=>dataOut_234_EXMPLR, F(233)=>
      dataOut_233_EXMPLR, F(232)=>dataOut_232_EXMPLR, F(231)=>
      dataOut_231_EXMPLR, F(230)=>dataOut_230_EXMPLR, F(229)=>
      dataOut_229_EXMPLR, F(228)=>dataOut_228_EXMPLR, F(227)=>
      dataOut_227_EXMPLR, F(226)=>dataOut_226_EXMPLR, F(225)=>
      dataOut_225_EXMPLR, F(224)=>dataOut_224_EXMPLR, F(223)=>
      dataOut_223_EXMPLR, F(222)=>dataOut_222_EXMPLR, F(221)=>
      dataOut_221_EXMPLR, F(220)=>dataOut_220_EXMPLR, F(219)=>
      dataOut_219_EXMPLR, F(218)=>dataOut_218_EXMPLR, F(217)=>
      dataOut_217_EXMPLR, F(216)=>dataOut_216_EXMPLR, F(215)=>
      dataOut_215_EXMPLR, F(214)=>dataOut_214_EXMPLR, F(213)=>
      dataOut_213_EXMPLR, F(212)=>dataOut_212_EXMPLR, F(211)=>
      dataOut_211_EXMPLR, F(210)=>dataOut_210_EXMPLR, F(209)=>
      dataOut_209_EXMPLR, F(208)=>dataOut_208_EXMPLR, F(207)=>
      dataOut_207_EXMPLR, F(206)=>dataOut_206_EXMPLR, F(205)=>
      dataOut_205_EXMPLR, F(204)=>dataOut_204_EXMPLR, F(203)=>
      dataOut_203_EXMPLR, F(202)=>dataOut_202_EXMPLR, F(201)=>
      dataOut_201_EXMPLR, F(200)=>dataOut_200_EXMPLR, F(199)=>
      dataOut_199_EXMPLR, F(198)=>dataOut_198_EXMPLR, F(197)=>
      dataOut_197_EXMPLR, F(196)=>dataOut_196_EXMPLR, F(195)=>
      dataOut_195_EXMPLR, F(194)=>dataOut_194_EXMPLR, F(193)=>
      dataOut_193_EXMPLR, F(192)=>dataOut_192_EXMPLR, F(191)=>
      dataOut_191_EXMPLR, F(190)=>dataOut_190_EXMPLR, F(189)=>
      dataOut_189_EXMPLR, F(188)=>dataOut_188_EXMPLR, F(187)=>
      dataOut_187_EXMPLR, F(186)=>dataOut_186_EXMPLR, F(185)=>
      dataOut_185_EXMPLR, F(184)=>dataOut_184_EXMPLR, F(183)=>
      dataOut_183_EXMPLR, F(182)=>dataOut_182_EXMPLR, F(181)=>
      dataOut_181_EXMPLR, F(180)=>dataOut_180_EXMPLR, F(179)=>
      dataOut_179_EXMPLR, F(178)=>dataOut_178_EXMPLR, F(177)=>
      dataOut_177_EXMPLR, F(176)=>dataOut_176_EXMPLR, F(175)=>
      dataOut_175_EXMPLR, F(174)=>dataOut_174_EXMPLR, F(173)=>
      dataOut_173_EXMPLR, F(172)=>dataOut_172_EXMPLR, F(171)=>
      dataOut_171_EXMPLR, F(170)=>dataOut_170_EXMPLR, F(169)=>
      dataOut_169_EXMPLR, F(168)=>dataOut_168_EXMPLR, F(167)=>
      dataOut_167_EXMPLR, F(166)=>dataOut_166_EXMPLR, F(165)=>
      dataOut_165_EXMPLR, F(164)=>dataOut_164_EXMPLR, F(163)=>
      dataOut_163_EXMPLR, F(162)=>dataOut_162_EXMPLR, F(161)=>
      dataOut_161_EXMPLR, F(160)=>dataOut_160_EXMPLR, F(159)=>
      dataOut_159_EXMPLR, F(158)=>dataOut_158_EXMPLR, F(157)=>
      dataOut_157_EXMPLR, F(156)=>dataOut_156_EXMPLR, F(155)=>
      dataOut_155_EXMPLR, F(154)=>dataOut_154_EXMPLR, F(153)=>
      dataOut_153_EXMPLR, F(152)=>dataOut_152_EXMPLR, F(151)=>
      dataOut_151_EXMPLR, F(150)=>dataOut_150_EXMPLR, F(149)=>
      dataOut_149_EXMPLR, F(148)=>dataOut_148_EXMPLR, F(147)=>
      dataOut_147_EXMPLR, F(146)=>dataOut_146_EXMPLR, F(145)=>
      dataOut_145_EXMPLR, F(144)=>dataOut_144_EXMPLR, F(143)=>
      dataOut_143_EXMPLR, F(142)=>dataOut_142_EXMPLR, F(141)=>
      dataOut_141_EXMPLR, F(140)=>dataOut_140_EXMPLR, F(139)=>
      dataOut_139_EXMPLR, F(138)=>dataOut_138_EXMPLR, F(137)=>
      dataOut_137_EXMPLR, F(136)=>dataOut_136_EXMPLR, F(135)=>
      dataOut_135_EXMPLR, F(134)=>dataOut_134_EXMPLR, F(133)=>
      dataOut_133_EXMPLR, F(132)=>dataOut_132_EXMPLR, F(131)=>
      dataOut_131_EXMPLR, F(130)=>dataOut_130_EXMPLR, F(129)=>
      dataOut_129_EXMPLR, F(128)=>dataOut_128_EXMPLR, F(127)=>
      dataOut_127_EXMPLR, F(126)=>dataOut_126_EXMPLR, F(125)=>
      dataOut_125_EXMPLR, F(124)=>dataOut_124_EXMPLR, F(123)=>
      dataOut_123_EXMPLR, F(122)=>dataOut_122_EXMPLR, F(121)=>
      dataOut_121_EXMPLR, F(120)=>dataOut_120_EXMPLR, F(119)=>
      dataOut_119_EXMPLR, F(118)=>dataOut_118_EXMPLR, F(117)=>
      dataOut_117_EXMPLR, F(116)=>dataOut_116_EXMPLR, F(115)=>
      dataOut_115_EXMPLR, F(114)=>dataOut_114_EXMPLR, F(113)=>
      dataOut_113_EXMPLR, F(112)=>dataOut_112_EXMPLR, F(111)=>
      dataOut_111_EXMPLR, F(110)=>dataOut_110_EXMPLR, F(109)=>
      dataOut_109_EXMPLR, F(108)=>dataOut_108_EXMPLR, F(107)=>
      dataOut_107_EXMPLR, F(106)=>dataOut_106_EXMPLR, F(105)=>
      dataOut_105_EXMPLR, F(104)=>dataOut_104_EXMPLR, F(103)=>
      dataOut_103_EXMPLR, F(102)=>dataOut_102_EXMPLR, F(101)=>
      dataOut_101_EXMPLR, F(100)=>dataOut_100_EXMPLR, F(99)=>
      dataOut_99_EXMPLR, F(98)=>dataOut_98_EXMPLR, F(97)=>dataOut_97_EXMPLR, 
      F(96)=>dataOut_96_EXMPLR, F(95)=>dataOut_95_EXMPLR, F(94)=>
      dataOut_94_EXMPLR, F(93)=>dataOut_93_EXMPLR, F(92)=>dataOut_92_EXMPLR, 
      F(91)=>dataOut_91_EXMPLR, F(90)=>dataOut_90_EXMPLR, F(89)=>
      dataOut_89_EXMPLR, F(88)=>dataOut_88_EXMPLR, F(87)=>dataOut_87_EXMPLR, 
      F(86)=>dataOut_86_EXMPLR, F(85)=>dataOut_85_EXMPLR, F(84)=>
      dataOut_84_EXMPLR, F(83)=>dataOut_83_EXMPLR, F(82)=>dataOut_82_EXMPLR, 
      F(81)=>dataOut_81_EXMPLR, F(80)=>dataOut_80_EXMPLR, F(79)=>
      dataOut_79_EXMPLR, F(78)=>dataOut_78_EXMPLR, F(77)=>dataOut_77_EXMPLR, 
      F(76)=>dataOut_76_EXMPLR, F(75)=>dataOut_75_EXMPLR, F(74)=>
      dataOut_74_EXMPLR, F(73)=>dataOut_73_EXMPLR, F(72)=>dataOut_72_EXMPLR, 
      F(71)=>dataOut_71_EXMPLR, F(70)=>dataOut_70_EXMPLR, F(69)=>
      dataOut_69_EXMPLR, F(68)=>dataOut_68_EXMPLR, F(67)=>dataOut_67_EXMPLR, 
      F(66)=>dataOut_66_EXMPLR, F(65)=>dataOut_65_EXMPLR, F(64)=>
      dataOut_64_EXMPLR, F(63)=>dataOut_63_EXMPLR, F(62)=>dataOut_62_EXMPLR, 
      F(61)=>dataOut_61_EXMPLR, F(60)=>dataOut_60_EXMPLR, F(59)=>
      dataOut_59_EXMPLR, F(58)=>dataOut_58_EXMPLR, F(57)=>dataOut_57_EXMPLR, 
      F(56)=>dataOut_56_EXMPLR, F(55)=>dataOut_55_EXMPLR, F(54)=>
      dataOut_54_EXMPLR, F(53)=>dataOut_53_EXMPLR, F(52)=>dataOut_52_EXMPLR, 
      F(51)=>dataOut_51_EXMPLR, F(50)=>dataOut_50_EXMPLR, F(49)=>
      dataOut_49_EXMPLR, F(48)=>dataOut_48_EXMPLR, F(47)=>dataOut_47_EXMPLR, 
      F(46)=>dataOut_46_EXMPLR, F(45)=>dataOut_45_EXMPLR, F(44)=>
      dataOut_44_EXMPLR, F(43)=>dataOut_43_EXMPLR, F(42)=>dataOut_42_EXMPLR, 
      F(41)=>dataOut_41_EXMPLR, F(40)=>dataOut_40_EXMPLR, F(39)=>
      dataOut_39_EXMPLR, F(38)=>dataOut_38_EXMPLR, F(37)=>dataOut_37_EXMPLR, 
      F(36)=>dataOut_36_EXMPLR, F(35)=>dataOut_35_EXMPLR, F(34)=>
      dataOut_34_EXMPLR, F(33)=>dataOut_33_EXMPLR, F(32)=>dataOut_32_EXMPLR, 
      F(31)=>dataOut_31_EXMPLR, F(30)=>dataOut_30_EXMPLR, F(29)=>
      dataOut_29_EXMPLR, F(28)=>dataOut_28_EXMPLR, F(27)=>dataOut_27_EXMPLR, 
      F(26)=>dataOut_26_EXMPLR, F(25)=>dataOut_25_EXMPLR, F(24)=>
      dataOut_24_EXMPLR, F(23)=>dataOut_23_EXMPLR, F(22)=>dataOut_22_EXMPLR, 
      F(21)=>dataOut_21_EXMPLR, F(20)=>dataOut_20_EXMPLR, F(19)=>
      dataOut_19_EXMPLR, F(18)=>dataOut_18_EXMPLR, F(17)=>dataOut_17_EXMPLR, 
      F(16)=>dataOut_16_EXMPLR, F(15)=>dataOut_15_EXMPLR, F(14)=>
      dataOut_14_EXMPLR, F(13)=>dataOut_13_EXMPLR, F(12)=>dataOut_12_EXMPLR, 
      F(11)=>dataOut_11_EXMPLR, F(10)=>dataOut_10_EXMPLR, F(9)=>
      dataOut_9_EXMPLR, F(8)=>dataOut_8_EXMPLR, F(7)=>dataOut_7_EXMPLR, F(6)
      =>dataOut_6_EXMPLR, F(5)=>dataOut_5_EXMPLR, F(4)=>dataOut_4_EXMPLR, 
      F(3)=>dataOut_3_EXMPLR, F(2)=>dataOut_2_EXMPLR, F(1)=>dataOut_1_EXMPLR, 
      F(0)=>dataOut_0_EXMPLR);
   Ram1Wr : triStateBuffer_16 port map ( D(15)=>dataIn(15), D(14)=>
      dataIn(14), D(13)=>dataIn(13), D(12)=>dataIn(12), D(11)=>dataIn(11), 
      D(10)=>dataIn(10), D(9)=>dataIn(9), D(8)=>dataIn(8), D(7)=>dataIn(7), 
      D(6)=>dataIn(6), D(5)=>dataIn(5), D(4)=>dataIn(4), D(3)=>dataIn(3), 
      D(2)=>dataIn(2), D(1)=>dataIn(1), D(0)=>dataIn(0), EN=>ram1Write, 
      F(15)=>dataToRam1_15, F(14)=>dataToRam1_14, F(13)=>dataToRam1_13, 
      F(12)=>dataToRam1_12, F(11)=>dataToRam1_11, F(10)=>dataToRam1_10, F(9)
      =>dataToRam1_9, F(8)=>dataToRam1_8, F(7)=>dataToRam1_7, F(6)=>
      dataToRam1_6, F(5)=>dataToRam1_5, F(4)=>dataToRam1_4, F(3)=>
      dataToRam1_3, F(2)=>dataToRam1_2, F(1)=>dataToRam1_1, F(0)=>
      dataToRam1_0);
   Ram2Rd : triStateBuffer_448 port map ( D(447)=>nx5785, D(446)=>nx5785, 
      D(445)=>nx5785, D(444)=>nx5785, D(443)=>nx5785, D(442)=>nx5785, D(441)
      =>nx5785, D(440)=>nx5787, D(439)=>nx5787, D(438)=>nx5787, D(437)=>
      nx5787, D(436)=>nx5787, D(435)=>nx5787, D(434)=>nx5787, D(433)=>nx5789, 
      D(432)=>nx5789, D(431)=>nx5789, D(430)=>nx5789, D(429)=>nx5789, D(428)
      =>nx5789, D(427)=>nx5789, D(426)=>nx5791, D(425)=>nx5791, D(424)=>
      nx5791, D(423)=>nx5791, D(422)=>nx5791, D(421)=>nx5791, D(420)=>nx5791, 
      D(419)=>nx5793, D(418)=>nx5793, D(417)=>nx5793, D(416)=>nx5793, D(415)
      =>nx5793, D(414)=>nx5793, D(413)=>nx5793, D(412)=>nx5795, D(411)=>
      nx5795, D(410)=>nx5795, D(409)=>nx5795, D(408)=>nx5795, D(407)=>nx5795, 
      D(406)=>nx5795, D(405)=>nx5797, D(404)=>nx5797, D(403)=>nx5797, D(402)
      =>nx5797, D(401)=>nx5797, D(400)=>nx5797, D(399)=>nx5797, D(398)=>
      nx5799, D(397)=>nx5799, D(396)=>nx5799, D(395)=>nx5799, D(394)=>nx5799, 
      D(393)=>nx5799, D(392)=>nx5799, D(391)=>nx5801, D(390)=>nx5801, D(389)
      =>nx5801, D(388)=>nx5801, D(387)=>nx5801, D(386)=>nx5801, D(385)=>
      nx5801, D(384)=>nx5803, D(383)=>nx5803, D(382)=>nx5803, D(381)=>nx5803, 
      D(380)=>nx5803, D(379)=>nx5803, D(378)=>nx5803, D(377)=>nx5805, D(376)
      =>nx5805, D(375)=>nx5805, D(374)=>nx5805, D(373)=>nx5805, D(372)=>
      nx5805, D(371)=>nx5805, D(370)=>nx5807, D(369)=>nx5807, D(368)=>nx5807, 
      D(367)=>nx5807, D(366)=>nx5807, D(365)=>nx5807, D(364)=>nx5807, D(363)
      =>nx5809, D(362)=>nx5809, D(361)=>nx5809, D(360)=>nx5809, D(359)=>
      nx5809, D(358)=>nx5809, D(357)=>nx5809, D(356)=>nx5811, D(355)=>nx5811, 
      D(354)=>nx5811, D(353)=>nx5811, D(352)=>nx5811, D(351)=>nx5811, D(350)
      =>nx5811, D(349)=>nx5813, D(348)=>nx5813, D(347)=>nx5813, D(346)=>
      nx5813, D(345)=>nx5813, D(344)=>nx5813, D(343)=>nx5813, D(342)=>nx5815, 
      D(341)=>nx5815, D(340)=>nx5815, D(339)=>nx5815, D(338)=>nx5815, D(337)
      =>nx5815, D(336)=>nx5815, D(335)=>nx5817, D(334)=>nx5817, D(333)=>
      nx5817, D(332)=>nx5817, D(331)=>nx5817, D(330)=>nx5817, D(329)=>nx5817, 
      D(328)=>nx5819, D(327)=>nx5819, D(326)=>nx5819, D(325)=>nx5819, D(324)
      =>nx5819, D(323)=>nx5819, D(322)=>nx5819, D(321)=>nx5821, D(320)=>
      nx5821, D(319)=>nx5821, D(318)=>nx5821, D(317)=>nx5821, D(316)=>nx5821, 
      D(315)=>nx5821, D(314)=>nx5823, D(313)=>nx5823, D(312)=>nx5823, D(311)
      =>nx5823, D(310)=>nx5823, D(309)=>nx5823, D(308)=>nx5823, D(307)=>
      nx5825, D(306)=>nx5825, D(305)=>nx5825, D(304)=>nx5825, D(303)=>nx5825, 
      D(302)=>nx5825, D(301)=>nx5825, D(300)=>nx5827, D(299)=>nx5827, D(298)
      =>nx5827, D(297)=>nx5827, D(296)=>nx5827, D(295)=>nx5827, D(294)=>
      nx5827, D(293)=>nx5829, D(292)=>nx5829, D(291)=>nx5829, D(290)=>nx5829, 
      D(289)=>nx5829, D(288)=>nx5829, D(287)=>nx5829, D(286)=>nx5831, D(285)
      =>nx5831, D(284)=>nx5831, D(283)=>nx5831, D(282)=>nx5831, D(281)=>
      nx5831, D(280)=>nx5831, D(279)=>nx5833, D(278)=>nx5833, D(277)=>nx5833, 
      D(276)=>nx5833, D(275)=>nx5833, D(274)=>nx5833, D(273)=>nx5833, D(272)
      =>nx5835, D(271)=>nx5835, D(270)=>nx5835, D(269)=>nx5835, D(268)=>
      nx5835, D(267)=>nx5835, D(266)=>nx5835, D(265)=>nx5837, D(264)=>nx5837, 
      D(263)=>nx5837, D(262)=>nx5837, D(261)=>nx5837, D(260)=>nx5837, D(259)
      =>nx5837, D(258)=>nx5839, D(257)=>nx5839, D(256)=>nx5839, D(255)=>
      nx5839, D(254)=>nx5839, D(253)=>nx5839, D(252)=>nx5839, D(251)=>nx5841, 
      D(250)=>nx5841, D(249)=>nx5841, D(248)=>nx5841, D(247)=>nx5841, D(246)
      =>nx5841, D(245)=>nx5841, D(244)=>nx5843, D(243)=>nx5843, D(242)=>
      nx5843, D(241)=>nx5843, D(240)=>nx5843, D(239)=>nx5843, D(238)=>nx5843, 
      D(237)=>nx5845, D(236)=>nx5845, D(235)=>nx5845, D(234)=>nx5845, D(233)
      =>nx5845, D(232)=>nx5845, D(231)=>nx5845, D(230)=>nx5847, D(229)=>
      nx5847, D(228)=>nx5847, D(227)=>nx5847, D(226)=>nx5847, D(225)=>nx5847, 
      D(224)=>nx5847, D(223)=>nx5849, D(222)=>nx5849, D(221)=>nx5849, D(220)
      =>nx5849, D(219)=>nx5849, D(218)=>nx5849, D(217)=>nx5849, D(216)=>
      nx5851, D(215)=>nx5851, D(214)=>nx5851, D(213)=>nx5851, D(212)=>nx5851, 
      D(211)=>nx5851, D(210)=>nx5851, D(209)=>nx5853, D(208)=>nx5853, D(207)
      =>nx5853, D(206)=>nx5853, D(205)=>nx5853, D(204)=>nx5853, D(203)=>
      nx5853, D(202)=>nx5855, D(201)=>nx5855, D(200)=>nx5855, D(199)=>nx5855, 
      D(198)=>nx5855, D(197)=>nx5855, D(196)=>nx5855, D(195)=>nx5857, D(194)
      =>nx5857, D(193)=>nx5857, D(192)=>nx5857, D(191)=>nx5857, D(190)=>
      nx5857, D(189)=>nx5857, D(188)=>nx5859, D(187)=>nx5859, D(186)=>nx5859, 
      D(185)=>nx5859, D(184)=>nx5859, D(183)=>nx5859, D(182)=>nx5859, D(181)
      =>nx5861, D(180)=>nx5861, D(179)=>nx5861, D(178)=>nx5861, D(177)=>
      nx5861, D(176)=>nx5861, D(175)=>nx5861, D(174)=>nx5863, D(173)=>nx5863, 
      D(172)=>nx5863, D(171)=>nx5863, D(170)=>nx5863, D(169)=>nx5863, D(168)
      =>nx5863, D(167)=>nx5865, D(166)=>nx5865, D(165)=>nx5865, D(164)=>
      nx5865, D(163)=>nx5865, D(162)=>nx5865, D(161)=>nx5865, D(160)=>nx5867, 
      D(159)=>nx5867, D(158)=>nx5867, D(157)=>nx5867, D(156)=>nx5867, D(155)
      =>nx5867, D(154)=>nx5867, D(153)=>nx5869, D(152)=>nx5869, D(151)=>
      nx5869, D(150)=>nx5869, D(149)=>nx5869, D(148)=>nx5869, D(147)=>nx5869, 
      D(146)=>nx5871, D(145)=>nx5871, D(144)=>nx5871, D(143)=>nx5871, D(142)
      =>nx5871, D(141)=>nx5871, D(140)=>nx5871, D(139)=>nx5873, D(138)=>
      nx5873, D(137)=>nx5873, D(136)=>nx5873, D(135)=>nx5873, D(134)=>nx5873, 
      D(133)=>nx5873, D(132)=>nx5875, D(131)=>nx5875, D(130)=>nx5875, D(129)
      =>nx5875, D(128)=>nx5875, D(127)=>nx5875, D(126)=>nx5875, D(125)=>
      nx5877, D(124)=>nx5877, D(123)=>nx5877, D(122)=>nx5877, D(121)=>nx5877, 
      D(120)=>nx5877, D(119)=>nx5877, D(118)=>nx5879, D(117)=>nx5879, D(116)
      =>nx5879, D(115)=>nx5879, D(114)=>nx5879, D(113)=>nx5879, D(112)=>
      nx5879, D(111)=>nx5881, D(110)=>nx5881, D(109)=>nx5881, D(108)=>nx5881, 
      D(107)=>nx5881, D(106)=>nx5881, D(105)=>nx5881, D(104)=>nx5883, D(103)
      =>nx5883, D(102)=>nx5883, D(101)=>nx5883, D(100)=>nx5883, D(99)=>
      nx5883, D(98)=>nx5883, D(97)=>nx5885, D(96)=>nx5885, D(95)=>nx5885, 
      D(94)=>nx5885, D(93)=>nx5885, D(92)=>nx5885, D(91)=>nx5885, D(90)=>
      nx5887, D(89)=>nx5887, D(88)=>nx5887, D(87)=>nx5887, D(86)=>nx5887, 
      D(85)=>nx5887, D(84)=>nx5887, D(83)=>nx5889, D(82)=>nx5889, D(81)=>
      nx5889, D(80)=>nx5889, D(79)=>nx5889, D(78)=>nx5889, D(77)=>nx5889, 
      D(76)=>nx5891, D(75)=>nx5891, D(74)=>nx5891, D(73)=>nx5891, D(72)=>
      nx5891, D(71)=>nx5891, D(70)=>nx5891, D(69)=>nx5893, D(68)=>nx5893, 
      D(67)=>nx5893, D(66)=>nx5893, D(65)=>nx5893, D(64)=>nx5893, D(63)=>
      nx5893, D(62)=>nx5895, D(61)=>nx5895, D(60)=>nx5895, D(59)=>nx5895, 
      D(58)=>nx5895, D(57)=>nx5895, D(56)=>nx5895, D(55)=>nx5897, D(54)=>
      nx5897, D(53)=>nx5897, D(52)=>nx5897, D(51)=>nx5897, D(50)=>nx5897, 
      D(49)=>nx5897, D(48)=>nx5899, D(47)=>nx5899, D(46)=>nx5899, D(45)=>
      nx5899, D(44)=>nx5899, D(43)=>nx5899, D(42)=>nx5899, D(41)=>nx5901, 
      D(40)=>nx5901, D(39)=>nx5901, D(38)=>nx5901, D(37)=>nx5901, D(36)=>
      nx5901, D(35)=>nx5901, D(34)=>nx5903, D(33)=>nx5903, D(32)=>nx5903, 
      D(31)=>nx5903, D(30)=>nx5903, D(29)=>nx5903, D(28)=>nx5903, D(27)=>
      nx5905, D(26)=>nx5905, D(25)=>nx5905, D(24)=>nx5905, D(23)=>nx5905, 
      D(22)=>nx5905, D(21)=>nx5905, D(20)=>nx5907, D(19)=>nx5907, D(18)=>
      nx5907, D(17)=>nx5907, D(16)=>nx5907, D(15)=>nx5907, D(14)=>nx5907, 
      D(13)=>nx5909, D(12)=>nx5909, D(11)=>nx5909, D(10)=>nx5909, D(9)=>
      nx5909, D(8)=>nx5909, D(7)=>nx5909, D(6)=>nx5911, D(5)=>nx5911, D(4)=>
      nx5911, D(3)=>nx5911, D(2)=>nx5911, D(1)=>nx5911, D(0)=>nx5911, EN=>
      DInput, F(447)=>dataOut_447_EXMPLR, F(446)=>dataOut_446_EXMPLR, F(445)
      =>dataOut_445_EXMPLR, F(444)=>dataOut_444_EXMPLR, F(443)=>
      dataOut_443_EXMPLR, F(442)=>dataOut_442_EXMPLR, F(441)=>
      dataOut_441_EXMPLR, F(440)=>dataOut_440_EXMPLR, F(439)=>
      dataOut_439_EXMPLR, F(438)=>dataOut_438_EXMPLR, F(437)=>
      dataOut_437_EXMPLR, F(436)=>dataOut_436_EXMPLR, F(435)=>
      dataOut_435_EXMPLR, F(434)=>dataOut_434_EXMPLR, F(433)=>
      dataOut_433_EXMPLR, F(432)=>dataOut_432_EXMPLR, F(431)=>
      dataOut_431_EXMPLR, F(430)=>dataOut_430_EXMPLR, F(429)=>
      dataOut_429_EXMPLR, F(428)=>dataOut_428_EXMPLR, F(427)=>
      dataOut_427_EXMPLR, F(426)=>dataOut_426_EXMPLR, F(425)=>
      dataOut_425_EXMPLR, F(424)=>dataOut_424_EXMPLR, F(423)=>
      dataOut_423_EXMPLR, F(422)=>dataOut_422_EXMPLR, F(421)=>
      dataOut_421_EXMPLR, F(420)=>dataOut_420_EXMPLR, F(419)=>
      dataOut_419_EXMPLR, F(418)=>dataOut_418_EXMPLR, F(417)=>
      dataOut_417_EXMPLR, F(416)=>dataOut_416_EXMPLR, F(415)=>
      dataOut_415_EXMPLR, F(414)=>dataOut_414_EXMPLR, F(413)=>
      dataOut_413_EXMPLR, F(412)=>dataOut_412_EXMPLR, F(411)=>
      dataOut_411_EXMPLR, F(410)=>dataOut_410_EXMPLR, F(409)=>
      dataOut_409_EXMPLR, F(408)=>dataOut_408_EXMPLR, F(407)=>
      dataOut_407_EXMPLR, F(406)=>dataOut_406_EXMPLR, F(405)=>
      dataOut_405_EXMPLR, F(404)=>dataOut_404_EXMPLR, F(403)=>
      dataOut_403_EXMPLR, F(402)=>dataOut_402_EXMPLR, F(401)=>
      dataOut_401_EXMPLR, F(400)=>dataOut_400_EXMPLR, F(399)=>
      dataOut_399_EXMPLR, F(398)=>dataOut_398_EXMPLR, F(397)=>
      dataOut_397_EXMPLR, F(396)=>dataOut_396_EXMPLR, F(395)=>
      dataOut_395_EXMPLR, F(394)=>dataOut_394_EXMPLR, F(393)=>
      dataOut_393_EXMPLR, F(392)=>dataOut_392_EXMPLR, F(391)=>
      dataOut_391_EXMPLR, F(390)=>dataOut_390_EXMPLR, F(389)=>
      dataOut_389_EXMPLR, F(388)=>dataOut_388_EXMPLR, F(387)=>
      dataOut_387_EXMPLR, F(386)=>dataOut_386_EXMPLR, F(385)=>
      dataOut_385_EXMPLR, F(384)=>dataOut_384_EXMPLR, F(383)=>
      dataOut_383_EXMPLR, F(382)=>dataOut_382_EXMPLR, F(381)=>
      dataOut_381_EXMPLR, F(380)=>dataOut_380_EXMPLR, F(379)=>
      dataOut_379_EXMPLR, F(378)=>dataOut_378_EXMPLR, F(377)=>
      dataOut_377_EXMPLR, F(376)=>dataOut_376_EXMPLR, F(375)=>
      dataOut_375_EXMPLR, F(374)=>dataOut_374_EXMPLR, F(373)=>
      dataOut_373_EXMPLR, F(372)=>dataOut_372_EXMPLR, F(371)=>
      dataOut_371_EXMPLR, F(370)=>dataOut_370_EXMPLR, F(369)=>
      dataOut_369_EXMPLR, F(368)=>dataOut_368_EXMPLR, F(367)=>
      dataOut_367_EXMPLR, F(366)=>dataOut_366_EXMPLR, F(365)=>
      dataOut_365_EXMPLR, F(364)=>dataOut_364_EXMPLR, F(363)=>
      dataOut_363_EXMPLR, F(362)=>dataOut_362_EXMPLR, F(361)=>
      dataOut_361_EXMPLR, F(360)=>dataOut_360_EXMPLR, F(359)=>
      dataOut_359_EXMPLR, F(358)=>dataOut_358_EXMPLR, F(357)=>
      dataOut_357_EXMPLR, F(356)=>dataOut_356_EXMPLR, F(355)=>
      dataOut_355_EXMPLR, F(354)=>dataOut_354_EXMPLR, F(353)=>
      dataOut_353_EXMPLR, F(352)=>dataOut_352_EXMPLR, F(351)=>
      dataOut_351_EXMPLR, F(350)=>dataOut_350_EXMPLR, F(349)=>
      dataOut_349_EXMPLR, F(348)=>dataOut_348_EXMPLR, F(347)=>
      dataOut_347_EXMPLR, F(346)=>dataOut_346_EXMPLR, F(345)=>
      dataOut_345_EXMPLR, F(344)=>dataOut_344_EXMPLR, F(343)=>
      dataOut_343_EXMPLR, F(342)=>dataOut_342_EXMPLR, F(341)=>
      dataOut_341_EXMPLR, F(340)=>dataOut_340_EXMPLR, F(339)=>
      dataOut_339_EXMPLR, F(338)=>dataOut_338_EXMPLR, F(337)=>
      dataOut_337_EXMPLR, F(336)=>dataOut_336_EXMPLR, F(335)=>
      dataOut_335_EXMPLR, F(334)=>dataOut_334_EXMPLR, F(333)=>
      dataOut_333_EXMPLR, F(332)=>dataOut_332_EXMPLR, F(331)=>
      dataOut_331_EXMPLR, F(330)=>dataOut_330_EXMPLR, F(329)=>
      dataOut_329_EXMPLR, F(328)=>dataOut_328_EXMPLR, F(327)=>
      dataOut_327_EXMPLR, F(326)=>dataOut_326_EXMPLR, F(325)=>
      dataOut_325_EXMPLR, F(324)=>dataOut_324_EXMPLR, F(323)=>
      dataOut_323_EXMPLR, F(322)=>dataOut_322_EXMPLR, F(321)=>
      dataOut_321_EXMPLR, F(320)=>dataOut_320_EXMPLR, F(319)=>
      dataOut_319_EXMPLR, F(318)=>dataOut_318_EXMPLR, F(317)=>
      dataOut_317_EXMPLR, F(316)=>dataOut_316_EXMPLR, F(315)=>
      dataOut_315_EXMPLR, F(314)=>dataOut_314_EXMPLR, F(313)=>
      dataOut_313_EXMPLR, F(312)=>dataOut_312_EXMPLR, F(311)=>
      dataOut_311_EXMPLR, F(310)=>dataOut_310_EXMPLR, F(309)=>
      dataOut_309_EXMPLR, F(308)=>dataOut_308_EXMPLR, F(307)=>
      dataOut_307_EXMPLR, F(306)=>dataOut_306_EXMPLR, F(305)=>
      dataOut_305_EXMPLR, F(304)=>dataOut_304_EXMPLR, F(303)=>
      dataOut_303_EXMPLR, F(302)=>dataOut_302_EXMPLR, F(301)=>
      dataOut_301_EXMPLR, F(300)=>dataOut_300_EXMPLR, F(299)=>
      dataOut_299_EXMPLR, F(298)=>dataOut_298_EXMPLR, F(297)=>
      dataOut_297_EXMPLR, F(296)=>dataOut_296_EXMPLR, F(295)=>
      dataOut_295_EXMPLR, F(294)=>dataOut_294_EXMPLR, F(293)=>
      dataOut_293_EXMPLR, F(292)=>dataOut_292_EXMPLR, F(291)=>
      dataOut_291_EXMPLR, F(290)=>dataOut_290_EXMPLR, F(289)=>
      dataOut_289_EXMPLR, F(288)=>dataOut_288_EXMPLR, F(287)=>
      dataOut_287_EXMPLR, F(286)=>dataOut_286_EXMPLR, F(285)=>
      dataOut_285_EXMPLR, F(284)=>dataOut_284_EXMPLR, F(283)=>
      dataOut_283_EXMPLR, F(282)=>dataOut_282_EXMPLR, F(281)=>
      dataOut_281_EXMPLR, F(280)=>dataOut_280_EXMPLR, F(279)=>
      dataOut_279_EXMPLR, F(278)=>dataOut_278_EXMPLR, F(277)=>
      dataOut_277_EXMPLR, F(276)=>dataOut_276_EXMPLR, F(275)=>
      dataOut_275_EXMPLR, F(274)=>dataOut_274_EXMPLR, F(273)=>
      dataOut_273_EXMPLR, F(272)=>dataOut_272_EXMPLR, F(271)=>
      dataOut_271_EXMPLR, F(270)=>dataOut_270_EXMPLR, F(269)=>
      dataOut_269_EXMPLR, F(268)=>dataOut_268_EXMPLR, F(267)=>
      dataOut_267_EXMPLR, F(266)=>dataOut_266_EXMPLR, F(265)=>
      dataOut_265_EXMPLR, F(264)=>dataOut_264_EXMPLR, F(263)=>
      dataOut_263_EXMPLR, F(262)=>dataOut_262_EXMPLR, F(261)=>
      dataOut_261_EXMPLR, F(260)=>dataOut_260_EXMPLR, F(259)=>
      dataOut_259_EXMPLR, F(258)=>dataOut_258_EXMPLR, F(257)=>
      dataOut_257_EXMPLR, F(256)=>dataOut_256_EXMPLR, F(255)=>
      dataOut_255_EXMPLR, F(254)=>dataOut_254_EXMPLR, F(253)=>
      dataOut_253_EXMPLR, F(252)=>dataOut_252_EXMPLR, F(251)=>
      dataOut_251_EXMPLR, F(250)=>dataOut_250_EXMPLR, F(249)=>
      dataOut_249_EXMPLR, F(248)=>dataOut_248_EXMPLR, F(247)=>
      dataOut_247_EXMPLR, F(246)=>dataOut_246_EXMPLR, F(245)=>
      dataOut_245_EXMPLR, F(244)=>dataOut_244_EXMPLR, F(243)=>
      dataOut_243_EXMPLR, F(242)=>dataOut_242_EXMPLR, F(241)=>
      dataOut_241_EXMPLR, F(240)=>dataOut_240_EXMPLR, F(239)=>
      dataOut_239_EXMPLR, F(238)=>dataOut_238_EXMPLR, F(237)=>
      dataOut_237_EXMPLR, F(236)=>dataOut_236_EXMPLR, F(235)=>
      dataOut_235_EXMPLR, F(234)=>dataOut_234_EXMPLR, F(233)=>
      dataOut_233_EXMPLR, F(232)=>dataOut_232_EXMPLR, F(231)=>
      dataOut_231_EXMPLR, F(230)=>dataOut_230_EXMPLR, F(229)=>
      dataOut_229_EXMPLR, F(228)=>dataOut_228_EXMPLR, F(227)=>
      dataOut_227_EXMPLR, F(226)=>dataOut_226_EXMPLR, F(225)=>
      dataOut_225_EXMPLR, F(224)=>dataOut_224_EXMPLR, F(223)=>
      dataOut_223_EXMPLR, F(222)=>dataOut_222_EXMPLR, F(221)=>
      dataOut_221_EXMPLR, F(220)=>dataOut_220_EXMPLR, F(219)=>
      dataOut_219_EXMPLR, F(218)=>dataOut_218_EXMPLR, F(217)=>
      dataOut_217_EXMPLR, F(216)=>dataOut_216_EXMPLR, F(215)=>
      dataOut_215_EXMPLR, F(214)=>dataOut_214_EXMPLR, F(213)=>
      dataOut_213_EXMPLR, F(212)=>dataOut_212_EXMPLR, F(211)=>
      dataOut_211_EXMPLR, F(210)=>dataOut_210_EXMPLR, F(209)=>
      dataOut_209_EXMPLR, F(208)=>dataOut_208_EXMPLR, F(207)=>
      dataOut_207_EXMPLR, F(206)=>dataOut_206_EXMPLR, F(205)=>
      dataOut_205_EXMPLR, F(204)=>dataOut_204_EXMPLR, F(203)=>
      dataOut_203_EXMPLR, F(202)=>dataOut_202_EXMPLR, F(201)=>
      dataOut_201_EXMPLR, F(200)=>dataOut_200_EXMPLR, F(199)=>
      dataOut_199_EXMPLR, F(198)=>dataOut_198_EXMPLR, F(197)=>
      dataOut_197_EXMPLR, F(196)=>dataOut_196_EXMPLR, F(195)=>
      dataOut_195_EXMPLR, F(194)=>dataOut_194_EXMPLR, F(193)=>
      dataOut_193_EXMPLR, F(192)=>dataOut_192_EXMPLR, F(191)=>
      dataOut_191_EXMPLR, F(190)=>dataOut_190_EXMPLR, F(189)=>
      dataOut_189_EXMPLR, F(188)=>dataOut_188_EXMPLR, F(187)=>
      dataOut_187_EXMPLR, F(186)=>dataOut_186_EXMPLR, F(185)=>
      dataOut_185_EXMPLR, F(184)=>dataOut_184_EXMPLR, F(183)=>
      dataOut_183_EXMPLR, F(182)=>dataOut_182_EXMPLR, F(181)=>
      dataOut_181_EXMPLR, F(180)=>dataOut_180_EXMPLR, F(179)=>
      dataOut_179_EXMPLR, F(178)=>dataOut_178_EXMPLR, F(177)=>
      dataOut_177_EXMPLR, F(176)=>dataOut_176_EXMPLR, F(175)=>
      dataOut_175_EXMPLR, F(174)=>dataOut_174_EXMPLR, F(173)=>
      dataOut_173_EXMPLR, F(172)=>dataOut_172_EXMPLR, F(171)=>
      dataOut_171_EXMPLR, F(170)=>dataOut_170_EXMPLR, F(169)=>
      dataOut_169_EXMPLR, F(168)=>dataOut_168_EXMPLR, F(167)=>
      dataOut_167_EXMPLR, F(166)=>dataOut_166_EXMPLR, F(165)=>
      dataOut_165_EXMPLR, F(164)=>dataOut_164_EXMPLR, F(163)=>
      dataOut_163_EXMPLR, F(162)=>dataOut_162_EXMPLR, F(161)=>
      dataOut_161_EXMPLR, F(160)=>dataOut_160_EXMPLR, F(159)=>
      dataOut_159_EXMPLR, F(158)=>dataOut_158_EXMPLR, F(157)=>
      dataOut_157_EXMPLR, F(156)=>dataOut_156_EXMPLR, F(155)=>
      dataOut_155_EXMPLR, F(154)=>dataOut_154_EXMPLR, F(153)=>
      dataOut_153_EXMPLR, F(152)=>dataOut_152_EXMPLR, F(151)=>
      dataOut_151_EXMPLR, F(150)=>dataOut_150_EXMPLR, F(149)=>
      dataOut_149_EXMPLR, F(148)=>dataOut_148_EXMPLR, F(147)=>
      dataOut_147_EXMPLR, F(146)=>dataOut_146_EXMPLR, F(145)=>
      dataOut_145_EXMPLR, F(144)=>dataOut_144_EXMPLR, F(143)=>
      dataOut_143_EXMPLR, F(142)=>dataOut_142_EXMPLR, F(141)=>
      dataOut_141_EXMPLR, F(140)=>dataOut_140_EXMPLR, F(139)=>
      dataOut_139_EXMPLR, F(138)=>dataOut_138_EXMPLR, F(137)=>
      dataOut_137_EXMPLR, F(136)=>dataOut_136_EXMPLR, F(135)=>
      dataOut_135_EXMPLR, F(134)=>dataOut_134_EXMPLR, F(133)=>
      dataOut_133_EXMPLR, F(132)=>dataOut_132_EXMPLR, F(131)=>
      dataOut_131_EXMPLR, F(130)=>dataOut_130_EXMPLR, F(129)=>
      dataOut_129_EXMPLR, F(128)=>dataOut_128_EXMPLR, F(127)=>
      dataOut_127_EXMPLR, F(126)=>dataOut_126_EXMPLR, F(125)=>
      dataOut_125_EXMPLR, F(124)=>dataOut_124_EXMPLR, F(123)=>
      dataOut_123_EXMPLR, F(122)=>dataOut_122_EXMPLR, F(121)=>
      dataOut_121_EXMPLR, F(120)=>dataOut_120_EXMPLR, F(119)=>
      dataOut_119_EXMPLR, F(118)=>dataOut_118_EXMPLR, F(117)=>
      dataOut_117_EXMPLR, F(116)=>dataOut_116_EXMPLR, F(115)=>
      dataOut_115_EXMPLR, F(114)=>dataOut_114_EXMPLR, F(113)=>
      dataOut_113_EXMPLR, F(112)=>dataOut_112_EXMPLR, F(111)=>
      dataOut_111_EXMPLR, F(110)=>dataOut_110_EXMPLR, F(109)=>
      dataOut_109_EXMPLR, F(108)=>dataOut_108_EXMPLR, F(107)=>
      dataOut_107_EXMPLR, F(106)=>dataOut_106_EXMPLR, F(105)=>
      dataOut_105_EXMPLR, F(104)=>dataOut_104_EXMPLR, F(103)=>
      dataOut_103_EXMPLR, F(102)=>dataOut_102_EXMPLR, F(101)=>
      dataOut_101_EXMPLR, F(100)=>dataOut_100_EXMPLR, F(99)=>
      dataOut_99_EXMPLR, F(98)=>dataOut_98_EXMPLR, F(97)=>dataOut_97_EXMPLR, 
      F(96)=>dataOut_96_EXMPLR, F(95)=>dataOut_95_EXMPLR, F(94)=>
      dataOut_94_EXMPLR, F(93)=>dataOut_93_EXMPLR, F(92)=>dataOut_92_EXMPLR, 
      F(91)=>dataOut_91_EXMPLR, F(90)=>dataOut_90_EXMPLR, F(89)=>
      dataOut_89_EXMPLR, F(88)=>dataOut_88_EXMPLR, F(87)=>dataOut_87_EXMPLR, 
      F(86)=>dataOut_86_EXMPLR, F(85)=>dataOut_85_EXMPLR, F(84)=>
      dataOut_84_EXMPLR, F(83)=>dataOut_83_EXMPLR, F(82)=>dataOut_82_EXMPLR, 
      F(81)=>dataOut_81_EXMPLR, F(80)=>dataOut_80_EXMPLR, F(79)=>
      dataOut_79_EXMPLR, F(78)=>dataOut_78_EXMPLR, F(77)=>dataOut_77_EXMPLR, 
      F(76)=>dataOut_76_EXMPLR, F(75)=>dataOut_75_EXMPLR, F(74)=>
      dataOut_74_EXMPLR, F(73)=>dataOut_73_EXMPLR, F(72)=>dataOut_72_EXMPLR, 
      F(71)=>dataOut_71_EXMPLR, F(70)=>dataOut_70_EXMPLR, F(69)=>
      dataOut_69_EXMPLR, F(68)=>dataOut_68_EXMPLR, F(67)=>dataOut_67_EXMPLR, 
      F(66)=>dataOut_66_EXMPLR, F(65)=>dataOut_65_EXMPLR, F(64)=>
      dataOut_64_EXMPLR, F(63)=>dataOut_63_EXMPLR, F(62)=>dataOut_62_EXMPLR, 
      F(61)=>dataOut_61_EXMPLR, F(60)=>dataOut_60_EXMPLR, F(59)=>
      dataOut_59_EXMPLR, F(58)=>dataOut_58_EXMPLR, F(57)=>dataOut_57_EXMPLR, 
      F(56)=>dataOut_56_EXMPLR, F(55)=>dataOut_55_EXMPLR, F(54)=>
      dataOut_54_EXMPLR, F(53)=>dataOut_53_EXMPLR, F(52)=>dataOut_52_EXMPLR, 
      F(51)=>dataOut_51_EXMPLR, F(50)=>dataOut_50_EXMPLR, F(49)=>
      dataOut_49_EXMPLR, F(48)=>dataOut_48_EXMPLR, F(47)=>dataOut_47_EXMPLR, 
      F(46)=>dataOut_46_EXMPLR, F(45)=>dataOut_45_EXMPLR, F(44)=>
      dataOut_44_EXMPLR, F(43)=>dataOut_43_EXMPLR, F(42)=>dataOut_42_EXMPLR, 
      F(41)=>dataOut_41_EXMPLR, F(40)=>dataOut_40_EXMPLR, F(39)=>
      dataOut_39_EXMPLR, F(38)=>dataOut_38_EXMPLR, F(37)=>dataOut_37_EXMPLR, 
      F(36)=>dataOut_36_EXMPLR, F(35)=>dataOut_35_EXMPLR, F(34)=>
      dataOut_34_EXMPLR, F(33)=>dataOut_33_EXMPLR, F(32)=>dataOut_32_EXMPLR, 
      F(31)=>dataOut_31_EXMPLR, F(30)=>dataOut_30_EXMPLR, F(29)=>
      dataOut_29_EXMPLR, F(28)=>dataOut_28_EXMPLR, F(27)=>dataOut_27_EXMPLR, 
      F(26)=>dataOut_26_EXMPLR, F(25)=>dataOut_25_EXMPLR, F(24)=>
      dataOut_24_EXMPLR, F(23)=>dataOut_23_EXMPLR, F(22)=>dataOut_22_EXMPLR, 
      F(21)=>dataOut_21_EXMPLR, F(20)=>dataOut_20_EXMPLR, F(19)=>
      dataOut_19_EXMPLR, F(18)=>dataOut_18_EXMPLR, F(17)=>dataOut_17_EXMPLR, 
      F(16)=>dataOut_16_EXMPLR, F(15)=>dataOut_15_EXMPLR, F(14)=>
      dataOut_14_EXMPLR, F(13)=>dataOut_13_EXMPLR, F(12)=>dataOut_12_EXMPLR, 
      F(11)=>dataOut_11_EXMPLR, F(10)=>dataOut_10_EXMPLR, F(9)=>
      dataOut_9_EXMPLR, F(8)=>dataOut_8_EXMPLR, F(7)=>dataOut_7_EXMPLR, F(6)
      =>dataOut_6_EXMPLR, F(5)=>dataOut_5_EXMPLR, F(4)=>dataOut_4_EXMPLR, 
      F(3)=>dataOut_3_EXMPLR, F(2)=>dataOut_2_EXMPLR, F(1)=>dataOut_1_EXMPLR, 
      F(0)=>dataOut_0_EXMPLR);
   Ram2Wr : triStateBuffer_16 port map ( D(15)=>dataIn(15), D(14)=>
      dataIn(14), D(13)=>dataIn(13), D(12)=>dataIn(12), D(11)=>dataIn(11), 
      D(10)=>dataIn(10), D(9)=>dataIn(9), D(8)=>dataIn(8), D(7)=>dataIn(7), 
      D(6)=>dataIn(6), D(5)=>dataIn(5), D(4)=>dataIn(4), D(3)=>dataIn(3), 
      D(2)=>dataIn(2), D(1)=>dataIn(1), D(0)=>dataIn(0), EN=>ram2Write, 
      F(15)=>dataToRam2_15, F(14)=>dataToRam2_14, F(13)=>dataToRam2_13, 
      F(12)=>dataToRam2_12, F(11)=>dataToRam2_11, F(10)=>dataToRam2_10, F(9)
      =>dataToRam2_9, F(8)=>dataToRam2_8, F(7)=>dataToRam2_7, F(6)=>
      dataToRam2_6, F(5)=>dataToRam2_5, F(4)=>dataToRam2_4, F(3)=>
      dataToRam2_3, F(2)=>dataToRam2_2, F(1)=>dataToRam2_1, F(0)=>
      dataToRam2_0);
   Ram1 : RAM_28 port map ( reset=>resetEN, CLK=>CLK, W=>ram1Write, R=>
      ram1Read, address(12)=>AddressIn(12), address(11)=>AddressIn(11), 
      address(10)=>AddressIn(10), address(9)=>AddressIn(9), address(8)=>
      AddressIn(8), address(7)=>AddressIn(7), address(6)=>AddressIn(6), 
      address(5)=>AddressIn(5), address(4)=>AddressIn(4), address(3)=>
      AddressIn(3), address(2)=>AddressIn(2), address(1)=>AddressIn(1), 
      address(0)=>AddressIn(0), dataIn(15)=>dataToRam1_15, dataIn(14)=>
      dataToRam1_14, dataIn(13)=>dataToRam1_13, dataIn(12)=>dataToRam1_12, 
      dataIn(11)=>dataToRam1_11, dataIn(10)=>dataToRam1_10, dataIn(9)=>
      dataToRam1_9, dataIn(8)=>dataToRam1_8, dataIn(7)=>dataToRam1_7, 
      dataIn(6)=>dataToRam1_6, dataIn(5)=>dataToRam1_5, dataIn(4)=>
      dataToRam1_4, dataIn(3)=>dataToRam1_3, dataIn(2)=>dataToRam1_2, 
      dataIn(1)=>dataToRam1_1, dataIn(0)=>dataToRam1_0, dataOut(447)=>
      dataFromRam1_447, dataOut(446)=>DANGLING(0), dataOut(445)=>DANGLING(1), 
      dataOut(444)=>DANGLING(2), dataOut(443)=>DANGLING(3), dataOut(442)=>
      DANGLING(4), dataOut(441)=>DANGLING(5), dataOut(440)=>DANGLING(6), 
      dataOut(439)=>DANGLING(7), dataOut(438)=>DANGLING(8), dataOut(437)=>
      DANGLING(9), dataOut(436)=>DANGLING(10), dataOut(435)=>DANGLING(11), 
      dataOut(434)=>DANGLING(12), dataOut(433)=>DANGLING(13), dataOut(432)=>
      DANGLING(14), dataOut(431)=>DANGLING(15), dataOut(430)=>DANGLING(16), 
      dataOut(429)=>DANGLING(17), dataOut(428)=>DANGLING(18), dataOut(427)=>
      DANGLING(19), dataOut(426)=>DANGLING(20), dataOut(425)=>DANGLING(21), 
      dataOut(424)=>DANGLING(22), dataOut(423)=>DANGLING(23), dataOut(422)=>
      DANGLING(24), dataOut(421)=>DANGLING(25), dataOut(420)=>DANGLING(26), 
      dataOut(419)=>DANGLING(27), dataOut(418)=>DANGLING(28), dataOut(417)=>
      DANGLING(29), dataOut(416)=>DANGLING(30), dataOut(415)=>DANGLING(31), 
      dataOut(414)=>DANGLING(32), dataOut(413)=>DANGLING(33), dataOut(412)=>
      DANGLING(34), dataOut(411)=>DANGLING(35), dataOut(410)=>DANGLING(36), 
      dataOut(409)=>DANGLING(37), dataOut(408)=>DANGLING(38), dataOut(407)=>
      DANGLING(39), dataOut(406)=>DANGLING(40), dataOut(405)=>DANGLING(41), 
      dataOut(404)=>DANGLING(42), dataOut(403)=>DANGLING(43), dataOut(402)=>
      DANGLING(44), dataOut(401)=>DANGLING(45), dataOut(400)=>DANGLING(46), 
      dataOut(399)=>DANGLING(47), dataOut(398)=>DANGLING(48), dataOut(397)=>
      DANGLING(49), dataOut(396)=>DANGLING(50), dataOut(395)=>DANGLING(51), 
      dataOut(394)=>DANGLING(52), dataOut(393)=>DANGLING(53), dataOut(392)=>
      DANGLING(54), dataOut(391)=>DANGLING(55), dataOut(390)=>DANGLING(56), 
      dataOut(389)=>DANGLING(57), dataOut(388)=>DANGLING(58), dataOut(387)=>
      DANGLING(59), dataOut(386)=>DANGLING(60), dataOut(385)=>DANGLING(61), 
      dataOut(384)=>DANGLING(62), dataOut(383)=>DANGLING(63), dataOut(382)=>
      DANGLING(64), dataOut(381)=>DANGLING(65), dataOut(380)=>DANGLING(66), 
      dataOut(379)=>DANGLING(67), dataOut(378)=>DANGLING(68), dataOut(377)=>
      DANGLING(69), dataOut(376)=>DANGLING(70), dataOut(375)=>DANGLING(71), 
      dataOut(374)=>DANGLING(72), dataOut(373)=>DANGLING(73), dataOut(372)=>
      DANGLING(74), dataOut(371)=>DANGLING(75), dataOut(370)=>DANGLING(76), 
      dataOut(369)=>DANGLING(77), dataOut(368)=>DANGLING(78), dataOut(367)=>
      DANGLING(79), dataOut(366)=>DANGLING(80), dataOut(365)=>DANGLING(81), 
      dataOut(364)=>DANGLING(82), dataOut(363)=>DANGLING(83), dataOut(362)=>
      DANGLING(84), dataOut(361)=>DANGLING(85), dataOut(360)=>DANGLING(86), 
      dataOut(359)=>DANGLING(87), dataOut(358)=>DANGLING(88), dataOut(357)=>
      DANGLING(89), dataOut(356)=>DANGLING(90), dataOut(355)=>DANGLING(91), 
      dataOut(354)=>DANGLING(92), dataOut(353)=>DANGLING(93), dataOut(352)=>
      DANGLING(94), dataOut(351)=>DANGLING(95), dataOut(350)=>DANGLING(96), 
      dataOut(349)=>DANGLING(97), dataOut(348)=>DANGLING(98), dataOut(347)=>
      DANGLING(99), dataOut(346)=>DANGLING(100), dataOut(345)=>DANGLING(101), 
      dataOut(344)=>DANGLING(102), dataOut(343)=>DANGLING(103), dataOut(342)
      =>DANGLING(104), dataOut(341)=>DANGLING(105), dataOut(340)=>DANGLING(
      106), dataOut(339)=>DANGLING(107), dataOut(338)=>DANGLING(108), 
      dataOut(337)=>DANGLING(109), dataOut(336)=>DANGLING(110), dataOut(335)
      =>DANGLING(111), dataOut(334)=>DANGLING(112), dataOut(333)=>DANGLING(
      113), dataOut(332)=>DANGLING(114), dataOut(331)=>DANGLING(115), 
      dataOut(330)=>DANGLING(116), dataOut(329)=>DANGLING(117), dataOut(328)
      =>DANGLING(118), dataOut(327)=>DANGLING(119), dataOut(326)=>DANGLING(
      120), dataOut(325)=>DANGLING(121), dataOut(324)=>DANGLING(122), 
      dataOut(323)=>DANGLING(123), dataOut(322)=>DANGLING(124), dataOut(321)
      =>DANGLING(125), dataOut(320)=>DANGLING(126), dataOut(319)=>DANGLING(
      127), dataOut(318)=>DANGLING(128), dataOut(317)=>DANGLING(129), 
      dataOut(316)=>DANGLING(130), dataOut(315)=>DANGLING(131), dataOut(314)
      =>DANGLING(132), dataOut(313)=>DANGLING(133), dataOut(312)=>DANGLING(
      134), dataOut(311)=>DANGLING(135), dataOut(310)=>DANGLING(136), 
      dataOut(309)=>DANGLING(137), dataOut(308)=>DANGLING(138), dataOut(307)
      =>DANGLING(139), dataOut(306)=>DANGLING(140), dataOut(305)=>DANGLING(
      141), dataOut(304)=>DANGLING(142), dataOut(303)=>DANGLING(143), 
      dataOut(302)=>DANGLING(144), dataOut(301)=>DANGLING(145), dataOut(300)
      =>DANGLING(146), dataOut(299)=>DANGLING(147), dataOut(298)=>DANGLING(
      148), dataOut(297)=>DANGLING(149), dataOut(296)=>DANGLING(150), 
      dataOut(295)=>DANGLING(151), dataOut(294)=>DANGLING(152), dataOut(293)
      =>DANGLING(153), dataOut(292)=>DANGLING(154), dataOut(291)=>DANGLING(
      155), dataOut(290)=>DANGLING(156), dataOut(289)=>DANGLING(157), 
      dataOut(288)=>DANGLING(158), dataOut(287)=>DANGLING(159), dataOut(286)
      =>DANGLING(160), dataOut(285)=>DANGLING(161), dataOut(284)=>DANGLING(
      162), dataOut(283)=>DANGLING(163), dataOut(282)=>DANGLING(164), 
      dataOut(281)=>DANGLING(165), dataOut(280)=>DANGLING(166), dataOut(279)
      =>DANGLING(167), dataOut(278)=>DANGLING(168), dataOut(277)=>DANGLING(
      169), dataOut(276)=>DANGLING(170), dataOut(275)=>DANGLING(171), 
      dataOut(274)=>DANGLING(172), dataOut(273)=>DANGLING(173), dataOut(272)
      =>DANGLING(174), dataOut(271)=>DANGLING(175), dataOut(270)=>DANGLING(
      176), dataOut(269)=>DANGLING(177), dataOut(268)=>DANGLING(178), 
      dataOut(267)=>DANGLING(179), dataOut(266)=>DANGLING(180), dataOut(265)
      =>DANGLING(181), dataOut(264)=>DANGLING(182), dataOut(263)=>DANGLING(
      183), dataOut(262)=>DANGLING(184), dataOut(261)=>DANGLING(185), 
      dataOut(260)=>DANGLING(186), dataOut(259)=>DANGLING(187), dataOut(258)
      =>DANGLING(188), dataOut(257)=>DANGLING(189), dataOut(256)=>DANGLING(
      190), dataOut(255)=>DANGLING(191), dataOut(254)=>DANGLING(192), 
      dataOut(253)=>DANGLING(193), dataOut(252)=>DANGLING(194), dataOut(251)
      =>DANGLING(195), dataOut(250)=>DANGLING(196), dataOut(249)=>DANGLING(
      197), dataOut(248)=>DANGLING(198), dataOut(247)=>DANGLING(199), 
      dataOut(246)=>DANGLING(200), dataOut(245)=>DANGLING(201), dataOut(244)
      =>DANGLING(202), dataOut(243)=>DANGLING(203), dataOut(242)=>DANGLING(
      204), dataOut(241)=>DANGLING(205), dataOut(240)=>DANGLING(206), 
      dataOut(239)=>DANGLING(207), dataOut(238)=>DANGLING(208), dataOut(237)
      =>DANGLING(209), dataOut(236)=>DANGLING(210), dataOut(235)=>DANGLING(
      211), dataOut(234)=>DANGLING(212), dataOut(233)=>DANGLING(213), 
      dataOut(232)=>DANGLING(214), dataOut(231)=>DANGLING(215), dataOut(230)
      =>DANGLING(216), dataOut(229)=>DANGLING(217), dataOut(228)=>DANGLING(
      218), dataOut(227)=>DANGLING(219), dataOut(226)=>DANGLING(220), 
      dataOut(225)=>DANGLING(221), dataOut(224)=>DANGLING(222), dataOut(223)
      =>DANGLING(223), dataOut(222)=>DANGLING(224), dataOut(221)=>DANGLING(
      225), dataOut(220)=>DANGLING(226), dataOut(219)=>DANGLING(227), 
      dataOut(218)=>DANGLING(228), dataOut(217)=>DANGLING(229), dataOut(216)
      =>DANGLING(230), dataOut(215)=>DANGLING(231), dataOut(214)=>DANGLING(
      232), dataOut(213)=>DANGLING(233), dataOut(212)=>DANGLING(234), 
      dataOut(211)=>DANGLING(235), dataOut(210)=>DANGLING(236), dataOut(209)
      =>DANGLING(237), dataOut(208)=>DANGLING(238), dataOut(207)=>DANGLING(
      239), dataOut(206)=>DANGLING(240), dataOut(205)=>DANGLING(241), 
      dataOut(204)=>DANGLING(242), dataOut(203)=>DANGLING(243), dataOut(202)
      =>DANGLING(244), dataOut(201)=>DANGLING(245), dataOut(200)=>DANGLING(
      246), dataOut(199)=>DANGLING(247), dataOut(198)=>DANGLING(248), 
      dataOut(197)=>DANGLING(249), dataOut(196)=>DANGLING(250), dataOut(195)
      =>DANGLING(251), dataOut(194)=>DANGLING(252), dataOut(193)=>DANGLING(
      253), dataOut(192)=>DANGLING(254), dataOut(191)=>DANGLING(255), 
      dataOut(190)=>DANGLING(256), dataOut(189)=>DANGLING(257), dataOut(188)
      =>DANGLING(258), dataOut(187)=>DANGLING(259), dataOut(186)=>DANGLING(
      260), dataOut(185)=>DANGLING(261), dataOut(184)=>DANGLING(262), 
      dataOut(183)=>DANGLING(263), dataOut(182)=>DANGLING(264), dataOut(181)
      =>DANGLING(265), dataOut(180)=>DANGLING(266), dataOut(179)=>DANGLING(
      267), dataOut(178)=>DANGLING(268), dataOut(177)=>DANGLING(269), 
      dataOut(176)=>DANGLING(270), dataOut(175)=>DANGLING(271), dataOut(174)
      =>DANGLING(272), dataOut(173)=>DANGLING(273), dataOut(172)=>DANGLING(
      274), dataOut(171)=>DANGLING(275), dataOut(170)=>DANGLING(276), 
      dataOut(169)=>DANGLING(277), dataOut(168)=>DANGLING(278), dataOut(167)
      =>DANGLING(279), dataOut(166)=>DANGLING(280), dataOut(165)=>DANGLING(
      281), dataOut(164)=>DANGLING(282), dataOut(163)=>DANGLING(283), 
      dataOut(162)=>DANGLING(284), dataOut(161)=>DANGLING(285), dataOut(160)
      =>DANGLING(286), dataOut(159)=>DANGLING(287), dataOut(158)=>DANGLING(
      288), dataOut(157)=>DANGLING(289), dataOut(156)=>DANGLING(290), 
      dataOut(155)=>DANGLING(291), dataOut(154)=>DANGLING(292), dataOut(153)
      =>DANGLING(293), dataOut(152)=>DANGLING(294), dataOut(151)=>DANGLING(
      295), dataOut(150)=>DANGLING(296), dataOut(149)=>DANGLING(297), 
      dataOut(148)=>DANGLING(298), dataOut(147)=>DANGLING(299), dataOut(146)
      =>DANGLING(300), dataOut(145)=>DANGLING(301), dataOut(144)=>DANGLING(
      302), dataOut(143)=>DANGLING(303), dataOut(142)=>DANGLING(304), 
      dataOut(141)=>DANGLING(305), dataOut(140)=>DANGLING(306), dataOut(139)
      =>DANGLING(307), dataOut(138)=>DANGLING(308), dataOut(137)=>DANGLING(
      309), dataOut(136)=>DANGLING(310), dataOut(135)=>DANGLING(311), 
      dataOut(134)=>DANGLING(312), dataOut(133)=>DANGLING(313), dataOut(132)
      =>DANGLING(314), dataOut(131)=>DANGLING(315), dataOut(130)=>DANGLING(
      316), dataOut(129)=>DANGLING(317), dataOut(128)=>DANGLING(318), 
      dataOut(127)=>DANGLING(319), dataOut(126)=>DANGLING(320), dataOut(125)
      =>DANGLING(321), dataOut(124)=>DANGLING(322), dataOut(123)=>DANGLING(
      323), dataOut(122)=>DANGLING(324), dataOut(121)=>DANGLING(325), 
      dataOut(120)=>DANGLING(326), dataOut(119)=>DANGLING(327), dataOut(118)
      =>DANGLING(328), dataOut(117)=>DANGLING(329), dataOut(116)=>DANGLING(
      330), dataOut(115)=>DANGLING(331), dataOut(114)=>DANGLING(332), 
      dataOut(113)=>DANGLING(333), dataOut(112)=>DANGLING(334), dataOut(111)
      =>DANGLING(335), dataOut(110)=>DANGLING(336), dataOut(109)=>DANGLING(
      337), dataOut(108)=>DANGLING(338), dataOut(107)=>DANGLING(339), 
      dataOut(106)=>DANGLING(340), dataOut(105)=>DANGLING(341), dataOut(104)
      =>DANGLING(342), dataOut(103)=>DANGLING(343), dataOut(102)=>DANGLING(
      344), dataOut(101)=>DANGLING(345), dataOut(100)=>DANGLING(346), 
      dataOut(99)=>DANGLING(347), dataOut(98)=>DANGLING(348), dataOut(97)=>
      DANGLING(349), dataOut(96)=>DANGLING(350), dataOut(95)=>DANGLING(351), 
      dataOut(94)=>DANGLING(352), dataOut(93)=>DANGLING(353), dataOut(92)=>
      DANGLING(354), dataOut(91)=>DANGLING(355), dataOut(90)=>DANGLING(356), 
      dataOut(89)=>DANGLING(357), dataOut(88)=>DANGLING(358), dataOut(87)=>
      DANGLING(359), dataOut(86)=>DANGLING(360), dataOut(85)=>DANGLING(361), 
      dataOut(84)=>DANGLING(362), dataOut(83)=>DANGLING(363), dataOut(82)=>
      DANGLING(364), dataOut(81)=>DANGLING(365), dataOut(80)=>DANGLING(366), 
      dataOut(79)=>DANGLING(367), dataOut(78)=>DANGLING(368), dataOut(77)=>
      DANGLING(369), dataOut(76)=>DANGLING(370), dataOut(75)=>DANGLING(371), 
      dataOut(74)=>DANGLING(372), dataOut(73)=>DANGLING(373), dataOut(72)=>
      DANGLING(374), dataOut(71)=>DANGLING(375), dataOut(70)=>DANGLING(376), 
      dataOut(69)=>DANGLING(377), dataOut(68)=>DANGLING(378), dataOut(67)=>
      DANGLING(379), dataOut(66)=>DANGLING(380), dataOut(65)=>DANGLING(381), 
      dataOut(64)=>DANGLING(382), dataOut(63)=>DANGLING(383), dataOut(62)=>
      DANGLING(384), dataOut(61)=>DANGLING(385), dataOut(60)=>DANGLING(386), 
      dataOut(59)=>DANGLING(387), dataOut(58)=>DANGLING(388), dataOut(57)=>
      DANGLING(389), dataOut(56)=>DANGLING(390), dataOut(55)=>DANGLING(391), 
      dataOut(54)=>DANGLING(392), dataOut(53)=>DANGLING(393), dataOut(52)=>
      DANGLING(394), dataOut(51)=>DANGLING(395), dataOut(50)=>DANGLING(396), 
      dataOut(49)=>DANGLING(397), dataOut(48)=>DANGLING(398), dataOut(47)=>
      DANGLING(399), dataOut(46)=>DANGLING(400), dataOut(45)=>DANGLING(401), 
      dataOut(44)=>DANGLING(402), dataOut(43)=>DANGLING(403), dataOut(42)=>
      DANGLING(404), dataOut(41)=>DANGLING(405), dataOut(40)=>DANGLING(406), 
      dataOut(39)=>DANGLING(407), dataOut(38)=>DANGLING(408), dataOut(37)=>
      DANGLING(409), dataOut(36)=>DANGLING(410), dataOut(35)=>DANGLING(411), 
      dataOut(34)=>DANGLING(412), dataOut(33)=>DANGLING(413), dataOut(32)=>
      DANGLING(414), dataOut(31)=>DANGLING(415), dataOut(30)=>DANGLING(416), 
      dataOut(29)=>DANGLING(417), dataOut(28)=>DANGLING(418), dataOut(27)=>
      DANGLING(419), dataOut(26)=>DANGLING(420), dataOut(25)=>DANGLING(421), 
      dataOut(24)=>DANGLING(422), dataOut(23)=>DANGLING(423), dataOut(22)=>
      DANGLING(424), dataOut(21)=>DANGLING(425), dataOut(20)=>DANGLING(426), 
      dataOut(19)=>DANGLING(427), dataOut(18)=>DANGLING(428), dataOut(17)=>
      DANGLING(429), dataOut(16)=>DANGLING(430), dataOut(15)=>DANGLING(431), 
      dataOut(14)=>DANGLING(432), dataOut(13)=>DANGLING(433), dataOut(12)=>
      DANGLING(434), dataOut(11)=>DANGLING(435), dataOut(10)=>DANGLING(436), 
      dataOut(9)=>DANGLING(437), dataOut(8)=>DANGLING(438), dataOut(7)=>
      DANGLING(439), dataOut(6)=>DANGLING(440), dataOut(5)=>DANGLING(441), 
      dataOut(4)=>DANGLING(442), dataOut(3)=>DANGLING(443), dataOut(2)=>
      DANGLING(444), dataOut(1)=>DANGLING(445), dataOut(0)=>DANGLING(446), 
      MFC=>mfcOfRam1, counterOut(3)=>DANGLING(447), counterOut(2)=>DANGLING(
      448), counterOut(1)=>DANGLING(449), counterOut(0)=>DANGLING(450));
   Ram2 : RAM_28 port map ( reset=>resetEN, CLK=>CLK, W=>ram2Write, R=>
      ram2Read, address(12)=>AddressIn(12), address(11)=>AddressIn(11), 
      address(10)=>AddressIn(10), address(9)=>AddressIn(9), address(8)=>
      AddressIn(8), address(7)=>AddressIn(7), address(6)=>AddressIn(6), 
      address(5)=>AddressIn(5), address(4)=>AddressIn(4), address(3)=>
      AddressIn(3), address(2)=>AddressIn(2), address(1)=>AddressIn(1), 
      address(0)=>AddressIn(0), dataIn(15)=>dataToRam2_15, dataIn(14)=>
      dataToRam2_14, dataIn(13)=>dataToRam2_13, dataIn(12)=>dataToRam2_12, 
      dataIn(11)=>dataToRam2_11, dataIn(10)=>dataToRam2_10, dataIn(9)=>
      dataToRam2_9, dataIn(8)=>dataToRam2_8, dataIn(7)=>dataToRam2_7, 
      dataIn(6)=>dataToRam2_6, dataIn(5)=>dataToRam2_5, dataIn(4)=>
      dataToRam2_4, dataIn(3)=>dataToRam2_3, dataIn(2)=>dataToRam2_2, 
      dataIn(1)=>dataToRam2_1, dataIn(0)=>dataToRam2_0, dataOut(447)=>
      dataFromRam2_447, dataOut(446)=>DANGLING(451), dataOut(445)=>DANGLING(
      452), dataOut(444)=>DANGLING(453), dataOut(443)=>DANGLING(454), 
      dataOut(442)=>DANGLING(455), dataOut(441)=>DANGLING(456), dataOut(440)
      =>DANGLING(457), dataOut(439)=>DANGLING(458), dataOut(438)=>DANGLING(
      459), dataOut(437)=>DANGLING(460), dataOut(436)=>DANGLING(461), 
      dataOut(435)=>DANGLING(462), dataOut(434)=>DANGLING(463), dataOut(433)
      =>DANGLING(464), dataOut(432)=>DANGLING(465), dataOut(431)=>DANGLING(
      466), dataOut(430)=>DANGLING(467), dataOut(429)=>DANGLING(468), 
      dataOut(428)=>DANGLING(469), dataOut(427)=>DANGLING(470), dataOut(426)
      =>DANGLING(471), dataOut(425)=>DANGLING(472), dataOut(424)=>DANGLING(
      473), dataOut(423)=>DANGLING(474), dataOut(422)=>DANGLING(475), 
      dataOut(421)=>DANGLING(476), dataOut(420)=>DANGLING(477), dataOut(419)
      =>DANGLING(478), dataOut(418)=>DANGLING(479), dataOut(417)=>DANGLING(
      480), dataOut(416)=>DANGLING(481), dataOut(415)=>DANGLING(482), 
      dataOut(414)=>DANGLING(483), dataOut(413)=>DANGLING(484), dataOut(412)
      =>DANGLING(485), dataOut(411)=>DANGLING(486), dataOut(410)=>DANGLING(
      487), dataOut(409)=>DANGLING(488), dataOut(408)=>DANGLING(489), 
      dataOut(407)=>DANGLING(490), dataOut(406)=>DANGLING(491), dataOut(405)
      =>DANGLING(492), dataOut(404)=>DANGLING(493), dataOut(403)=>DANGLING(
      494), dataOut(402)=>DANGLING(495), dataOut(401)=>DANGLING(496), 
      dataOut(400)=>DANGLING(497), dataOut(399)=>DANGLING(498), dataOut(398)
      =>DANGLING(499), dataOut(397)=>DANGLING(500), dataOut(396)=>DANGLING(
      501), dataOut(395)=>DANGLING(502), dataOut(394)=>DANGLING(503), 
      dataOut(393)=>DANGLING(504), dataOut(392)=>DANGLING(505), dataOut(391)
      =>DANGLING(506), dataOut(390)=>DANGLING(507), dataOut(389)=>DANGLING(
      508), dataOut(388)=>DANGLING(509), dataOut(387)=>DANGLING(510), 
      dataOut(386)=>DANGLING(511), dataOut(385)=>DANGLING(512), dataOut(384)
      =>DANGLING(513), dataOut(383)=>DANGLING(514), dataOut(382)=>DANGLING(
      515), dataOut(381)=>DANGLING(516), dataOut(380)=>DANGLING(517), 
      dataOut(379)=>DANGLING(518), dataOut(378)=>DANGLING(519), dataOut(377)
      =>DANGLING(520), dataOut(376)=>DANGLING(521), dataOut(375)=>DANGLING(
      522), dataOut(374)=>DANGLING(523), dataOut(373)=>DANGLING(524), 
      dataOut(372)=>DANGLING(525), dataOut(371)=>DANGLING(526), dataOut(370)
      =>DANGLING(527), dataOut(369)=>DANGLING(528), dataOut(368)=>DANGLING(
      529), dataOut(367)=>DANGLING(530), dataOut(366)=>DANGLING(531), 
      dataOut(365)=>DANGLING(532), dataOut(364)=>DANGLING(533), dataOut(363)
      =>DANGLING(534), dataOut(362)=>DANGLING(535), dataOut(361)=>DANGLING(
      536), dataOut(360)=>DANGLING(537), dataOut(359)=>DANGLING(538), 
      dataOut(358)=>DANGLING(539), dataOut(357)=>DANGLING(540), dataOut(356)
      =>DANGLING(541), dataOut(355)=>DANGLING(542), dataOut(354)=>DANGLING(
      543), dataOut(353)=>DANGLING(544), dataOut(352)=>DANGLING(545), 
      dataOut(351)=>DANGLING(546), dataOut(350)=>DANGLING(547), dataOut(349)
      =>DANGLING(548), dataOut(348)=>DANGLING(549), dataOut(347)=>DANGLING(
      550), dataOut(346)=>DANGLING(551), dataOut(345)=>DANGLING(552), 
      dataOut(344)=>DANGLING(553), dataOut(343)=>DANGLING(554), dataOut(342)
      =>DANGLING(555), dataOut(341)=>DANGLING(556), dataOut(340)=>DANGLING(
      557), dataOut(339)=>DANGLING(558), dataOut(338)=>DANGLING(559), 
      dataOut(337)=>DANGLING(560), dataOut(336)=>DANGLING(561), dataOut(335)
      =>DANGLING(562), dataOut(334)=>DANGLING(563), dataOut(333)=>DANGLING(
      564), dataOut(332)=>DANGLING(565), dataOut(331)=>DANGLING(566), 
      dataOut(330)=>DANGLING(567), dataOut(329)=>DANGLING(568), dataOut(328)
      =>DANGLING(569), dataOut(327)=>DANGLING(570), dataOut(326)=>DANGLING(
      571), dataOut(325)=>DANGLING(572), dataOut(324)=>DANGLING(573), 
      dataOut(323)=>DANGLING(574), dataOut(322)=>DANGLING(575), dataOut(321)
      =>DANGLING(576), dataOut(320)=>DANGLING(577), dataOut(319)=>DANGLING(
      578), dataOut(318)=>DANGLING(579), dataOut(317)=>DANGLING(580), 
      dataOut(316)=>DANGLING(581), dataOut(315)=>DANGLING(582), dataOut(314)
      =>DANGLING(583), dataOut(313)=>DANGLING(584), dataOut(312)=>DANGLING(
      585), dataOut(311)=>DANGLING(586), dataOut(310)=>DANGLING(587), 
      dataOut(309)=>DANGLING(588), dataOut(308)=>DANGLING(589), dataOut(307)
      =>DANGLING(590), dataOut(306)=>DANGLING(591), dataOut(305)=>DANGLING(
      592), dataOut(304)=>DANGLING(593), dataOut(303)=>DANGLING(594), 
      dataOut(302)=>DANGLING(595), dataOut(301)=>DANGLING(596), dataOut(300)
      =>DANGLING(597), dataOut(299)=>DANGLING(598), dataOut(298)=>DANGLING(
      599), dataOut(297)=>DANGLING(600), dataOut(296)=>DANGLING(601), 
      dataOut(295)=>DANGLING(602), dataOut(294)=>DANGLING(603), dataOut(293)
      =>DANGLING(604), dataOut(292)=>DANGLING(605), dataOut(291)=>DANGLING(
      606), dataOut(290)=>DANGLING(607), dataOut(289)=>DANGLING(608), 
      dataOut(288)=>DANGLING(609), dataOut(287)=>DANGLING(610), dataOut(286)
      =>DANGLING(611), dataOut(285)=>DANGLING(612), dataOut(284)=>DANGLING(
      613), dataOut(283)=>DANGLING(614), dataOut(282)=>DANGLING(615), 
      dataOut(281)=>DANGLING(616), dataOut(280)=>DANGLING(617), dataOut(279)
      =>DANGLING(618), dataOut(278)=>DANGLING(619), dataOut(277)=>DANGLING(
      620), dataOut(276)=>DANGLING(621), dataOut(275)=>DANGLING(622), 
      dataOut(274)=>DANGLING(623), dataOut(273)=>DANGLING(624), dataOut(272)
      =>DANGLING(625), dataOut(271)=>DANGLING(626), dataOut(270)=>DANGLING(
      627), dataOut(269)=>DANGLING(628), dataOut(268)=>DANGLING(629), 
      dataOut(267)=>DANGLING(630), dataOut(266)=>DANGLING(631), dataOut(265)
      =>DANGLING(632), dataOut(264)=>DANGLING(633), dataOut(263)=>DANGLING(
      634), dataOut(262)=>DANGLING(635), dataOut(261)=>DANGLING(636), 
      dataOut(260)=>DANGLING(637), dataOut(259)=>DANGLING(638), dataOut(258)
      =>DANGLING(639), dataOut(257)=>DANGLING(640), dataOut(256)=>DANGLING(
      641), dataOut(255)=>DANGLING(642), dataOut(254)=>DANGLING(643), 
      dataOut(253)=>DANGLING(644), dataOut(252)=>DANGLING(645), dataOut(251)
      =>DANGLING(646), dataOut(250)=>DANGLING(647), dataOut(249)=>DANGLING(
      648), dataOut(248)=>DANGLING(649), dataOut(247)=>DANGLING(650), 
      dataOut(246)=>DANGLING(651), dataOut(245)=>DANGLING(652), dataOut(244)
      =>DANGLING(653), dataOut(243)=>DANGLING(654), dataOut(242)=>DANGLING(
      655), dataOut(241)=>DANGLING(656), dataOut(240)=>DANGLING(657), 
      dataOut(239)=>DANGLING(658), dataOut(238)=>DANGLING(659), dataOut(237)
      =>DANGLING(660), dataOut(236)=>DANGLING(661), dataOut(235)=>DANGLING(
      662), dataOut(234)=>DANGLING(663), dataOut(233)=>DANGLING(664), 
      dataOut(232)=>DANGLING(665), dataOut(231)=>DANGLING(666), dataOut(230)
      =>DANGLING(667), dataOut(229)=>DANGLING(668), dataOut(228)=>DANGLING(
      669), dataOut(227)=>DANGLING(670), dataOut(226)=>DANGLING(671), 
      dataOut(225)=>DANGLING(672), dataOut(224)=>DANGLING(673), dataOut(223)
      =>DANGLING(674), dataOut(222)=>DANGLING(675), dataOut(221)=>DANGLING(
      676), dataOut(220)=>DANGLING(677), dataOut(219)=>DANGLING(678), 
      dataOut(218)=>DANGLING(679), dataOut(217)=>DANGLING(680), dataOut(216)
      =>DANGLING(681), dataOut(215)=>DANGLING(682), dataOut(214)=>DANGLING(
      683), dataOut(213)=>DANGLING(684), dataOut(212)=>DANGLING(685), 
      dataOut(211)=>DANGLING(686), dataOut(210)=>DANGLING(687), dataOut(209)
      =>DANGLING(688), dataOut(208)=>DANGLING(689), dataOut(207)=>DANGLING(
      690), dataOut(206)=>DANGLING(691), dataOut(205)=>DANGLING(692), 
      dataOut(204)=>DANGLING(693), dataOut(203)=>DANGLING(694), dataOut(202)
      =>DANGLING(695), dataOut(201)=>DANGLING(696), dataOut(200)=>DANGLING(
      697), dataOut(199)=>DANGLING(698), dataOut(198)=>DANGLING(699), 
      dataOut(197)=>DANGLING(700), dataOut(196)=>DANGLING(701), dataOut(195)
      =>DANGLING(702), dataOut(194)=>DANGLING(703), dataOut(193)=>DANGLING(
      704), dataOut(192)=>DANGLING(705), dataOut(191)=>DANGLING(706), 
      dataOut(190)=>DANGLING(707), dataOut(189)=>DANGLING(708), dataOut(188)
      =>DANGLING(709), dataOut(187)=>DANGLING(710), dataOut(186)=>DANGLING(
      711), dataOut(185)=>DANGLING(712), dataOut(184)=>DANGLING(713), 
      dataOut(183)=>DANGLING(714), dataOut(182)=>DANGLING(715), dataOut(181)
      =>DANGLING(716), dataOut(180)=>DANGLING(717), dataOut(179)=>DANGLING(
      718), dataOut(178)=>DANGLING(719), dataOut(177)=>DANGLING(720), 
      dataOut(176)=>DANGLING(721), dataOut(175)=>DANGLING(722), dataOut(174)
      =>DANGLING(723), dataOut(173)=>DANGLING(724), dataOut(172)=>DANGLING(
      725), dataOut(171)=>DANGLING(726), dataOut(170)=>DANGLING(727), 
      dataOut(169)=>DANGLING(728), dataOut(168)=>DANGLING(729), dataOut(167)
      =>DANGLING(730), dataOut(166)=>DANGLING(731), dataOut(165)=>DANGLING(
      732), dataOut(164)=>DANGLING(733), dataOut(163)=>DANGLING(734), 
      dataOut(162)=>DANGLING(735), dataOut(161)=>DANGLING(736), dataOut(160)
      =>DANGLING(737), dataOut(159)=>DANGLING(738), dataOut(158)=>DANGLING(
      739), dataOut(157)=>DANGLING(740), dataOut(156)=>DANGLING(741), 
      dataOut(155)=>DANGLING(742), dataOut(154)=>DANGLING(743), dataOut(153)
      =>DANGLING(744), dataOut(152)=>DANGLING(745), dataOut(151)=>DANGLING(
      746), dataOut(150)=>DANGLING(747), dataOut(149)=>DANGLING(748), 
      dataOut(148)=>DANGLING(749), dataOut(147)=>DANGLING(750), dataOut(146)
      =>DANGLING(751), dataOut(145)=>DANGLING(752), dataOut(144)=>DANGLING(
      753), dataOut(143)=>DANGLING(754), dataOut(142)=>DANGLING(755), 
      dataOut(141)=>DANGLING(756), dataOut(140)=>DANGLING(757), dataOut(139)
      =>DANGLING(758), dataOut(138)=>DANGLING(759), dataOut(137)=>DANGLING(
      760), dataOut(136)=>DANGLING(761), dataOut(135)=>DANGLING(762), 
      dataOut(134)=>DANGLING(763), dataOut(133)=>DANGLING(764), dataOut(132)
      =>DANGLING(765), dataOut(131)=>DANGLING(766), dataOut(130)=>DANGLING(
      767), dataOut(129)=>DANGLING(768), dataOut(128)=>DANGLING(769), 
      dataOut(127)=>DANGLING(770), dataOut(126)=>DANGLING(771), dataOut(125)
      =>DANGLING(772), dataOut(124)=>DANGLING(773), dataOut(123)=>DANGLING(
      774), dataOut(122)=>DANGLING(775), dataOut(121)=>DANGLING(776), 
      dataOut(120)=>DANGLING(777), dataOut(119)=>DANGLING(778), dataOut(118)
      =>DANGLING(779), dataOut(117)=>DANGLING(780), dataOut(116)=>DANGLING(
      781), dataOut(115)=>DANGLING(782), dataOut(114)=>DANGLING(783), 
      dataOut(113)=>DANGLING(784), dataOut(112)=>DANGLING(785), dataOut(111)
      =>DANGLING(786), dataOut(110)=>DANGLING(787), dataOut(109)=>DANGLING(
      788), dataOut(108)=>DANGLING(789), dataOut(107)=>DANGLING(790), 
      dataOut(106)=>DANGLING(791), dataOut(105)=>DANGLING(792), dataOut(104)
      =>DANGLING(793), dataOut(103)=>DANGLING(794), dataOut(102)=>DANGLING(
      795), dataOut(101)=>DANGLING(796), dataOut(100)=>DANGLING(797), 
      dataOut(99)=>DANGLING(798), dataOut(98)=>DANGLING(799), dataOut(97)=>
      DANGLING(800), dataOut(96)=>DANGLING(801), dataOut(95)=>DANGLING(802), 
      dataOut(94)=>DANGLING(803), dataOut(93)=>DANGLING(804), dataOut(92)=>
      DANGLING(805), dataOut(91)=>DANGLING(806), dataOut(90)=>DANGLING(807), 
      dataOut(89)=>DANGLING(808), dataOut(88)=>DANGLING(809), dataOut(87)=>
      DANGLING(810), dataOut(86)=>DANGLING(811), dataOut(85)=>DANGLING(812), 
      dataOut(84)=>DANGLING(813), dataOut(83)=>DANGLING(814), dataOut(82)=>
      DANGLING(815), dataOut(81)=>DANGLING(816), dataOut(80)=>DANGLING(817), 
      dataOut(79)=>DANGLING(818), dataOut(78)=>DANGLING(819), dataOut(77)=>
      DANGLING(820), dataOut(76)=>DANGLING(821), dataOut(75)=>DANGLING(822), 
      dataOut(74)=>DANGLING(823), dataOut(73)=>DANGLING(824), dataOut(72)=>
      DANGLING(825), dataOut(71)=>DANGLING(826), dataOut(70)=>DANGLING(827), 
      dataOut(69)=>DANGLING(828), dataOut(68)=>DANGLING(829), dataOut(67)=>
      DANGLING(830), dataOut(66)=>DANGLING(831), dataOut(65)=>DANGLING(832), 
      dataOut(64)=>DANGLING(833), dataOut(63)=>DANGLING(834), dataOut(62)=>
      DANGLING(835), dataOut(61)=>DANGLING(836), dataOut(60)=>DANGLING(837), 
      dataOut(59)=>DANGLING(838), dataOut(58)=>DANGLING(839), dataOut(57)=>
      DANGLING(840), dataOut(56)=>DANGLING(841), dataOut(55)=>DANGLING(842), 
      dataOut(54)=>DANGLING(843), dataOut(53)=>DANGLING(844), dataOut(52)=>
      DANGLING(845), dataOut(51)=>DANGLING(846), dataOut(50)=>DANGLING(847), 
      dataOut(49)=>DANGLING(848), dataOut(48)=>DANGLING(849), dataOut(47)=>
      DANGLING(850), dataOut(46)=>DANGLING(851), dataOut(45)=>DANGLING(852), 
      dataOut(44)=>DANGLING(853), dataOut(43)=>DANGLING(854), dataOut(42)=>
      DANGLING(855), dataOut(41)=>DANGLING(856), dataOut(40)=>DANGLING(857), 
      dataOut(39)=>DANGLING(858), dataOut(38)=>DANGLING(859), dataOut(37)=>
      DANGLING(860), dataOut(36)=>DANGLING(861), dataOut(35)=>DANGLING(862), 
      dataOut(34)=>DANGLING(863), dataOut(33)=>DANGLING(864), dataOut(32)=>
      DANGLING(865), dataOut(31)=>DANGLING(866), dataOut(30)=>DANGLING(867), 
      dataOut(29)=>DANGLING(868), dataOut(28)=>DANGLING(869), dataOut(27)=>
      DANGLING(870), dataOut(26)=>DANGLING(871), dataOut(25)=>DANGLING(872), 
      dataOut(24)=>DANGLING(873), dataOut(23)=>DANGLING(874), dataOut(22)=>
      DANGLING(875), dataOut(21)=>DANGLING(876), dataOut(20)=>DANGLING(877), 
      dataOut(19)=>DANGLING(878), dataOut(18)=>DANGLING(879), dataOut(17)=>
      DANGLING(880), dataOut(16)=>DANGLING(881), dataOut(15)=>DANGLING(882), 
      dataOut(14)=>DANGLING(883), dataOut(13)=>DANGLING(884), dataOut(12)=>
      DANGLING(885), dataOut(11)=>DANGLING(886), dataOut(10)=>DANGLING(887), 
      dataOut(9)=>DANGLING(888), dataOut(8)=>DANGLING(889), dataOut(7)=>
      DANGLING(890), dataOut(6)=>DANGLING(891), dataOut(5)=>DANGLING(892), 
      dataOut(4)=>DANGLING(893), dataOut(3)=>DANGLING(894), dataOut(2)=>
      DANGLING(895), dataOut(1)=>DANGLING(896), dataOut(0)=>DANGLING(897), 
      MFC=>mfcOfRam2, counterOut(3)=>DANGLING(898), counterOut(2)=>DANGLING(
      899), counterOut(1)=>DANGLING(900), counterOut(0)=>DANGLING(901));
   ix5633 : fake_vcc port map ( Y=>nx5632);
   ix5636 : xnor2 port map ( Y=>test, A0=>switcherEN, A1=>ramSelector);
   ix5623 : fake_gnd port map ( Y=>GND);
   tri_counterOut_0 : tri01 port map ( Y=>counterOut(0), A=>nx5632, E=>GND);
   tri_counterOut_1 : tri01 port map ( Y=>counterOut(1), A=>nx5632, E=>GND);
   tri_counterOut_2 : tri01 port map ( Y=>counterOut(2), A=>nx5632, E=>GND);
   tri_counterOut_3 : tri01 port map ( Y=>counterOut(3), A=>nx5632, E=>GND);
   ix1 : inv01 port map ( Y=>DInput, A=>test);
   ix5652 : inv01 port map ( Y=>nx5653, A=>dataFromRam1_447);
   ix5654 : inv01 port map ( Y=>nx5655, A=>nx5913);
   ix5656 : inv01 port map ( Y=>nx5657, A=>nx5913);
   ix5658 : inv01 port map ( Y=>nx5659, A=>nx5913);
   ix5660 : inv01 port map ( Y=>nx5661, A=>nx5913);
   ix5662 : inv01 port map ( Y=>nx5663, A=>nx5913);
   ix5664 : inv01 port map ( Y=>nx5665, A=>nx5913);
   ix5666 : inv01 port map ( Y=>nx5667, A=>nx5913);
   ix5668 : inv01 port map ( Y=>nx5669, A=>nx5915);
   ix5670 : inv01 port map ( Y=>nx5671, A=>nx5915);
   ix5672 : inv01 port map ( Y=>nx5673, A=>nx5915);
   ix5674 : inv01 port map ( Y=>nx5675, A=>nx5915);
   ix5676 : inv01 port map ( Y=>nx5677, A=>nx5915);
   ix5678 : inv01 port map ( Y=>nx5679, A=>nx5915);
   ix5680 : inv01 port map ( Y=>nx5681, A=>nx5915);
   ix5682 : inv01 port map ( Y=>nx5683, A=>nx5917);
   ix5684 : inv01 port map ( Y=>nx5685, A=>nx5917);
   ix5686 : inv01 port map ( Y=>nx5687, A=>nx5917);
   ix5688 : inv01 port map ( Y=>nx5689, A=>nx5917);
   ix5690 : inv01 port map ( Y=>nx5691, A=>nx5917);
   ix5692 : inv01 port map ( Y=>nx5693, A=>nx5917);
   ix5694 : inv01 port map ( Y=>nx5695, A=>nx5917);
   ix5696 : inv01 port map ( Y=>nx5697, A=>nx5919);
   ix5698 : inv01 port map ( Y=>nx5699, A=>nx5919);
   ix5700 : inv01 port map ( Y=>nx5701, A=>nx5919);
   ix5702 : inv01 port map ( Y=>nx5703, A=>nx5919);
   ix5704 : inv01 port map ( Y=>nx5705, A=>nx5919);
   ix5706 : inv01 port map ( Y=>nx5707, A=>nx5919);
   ix5708 : inv01 port map ( Y=>nx5709, A=>nx5919);
   ix5710 : inv01 port map ( Y=>nx5711, A=>nx5921);
   ix5712 : inv01 port map ( Y=>nx5713, A=>nx5921);
   ix5714 : inv01 port map ( Y=>nx5715, A=>nx5921);
   ix5716 : inv01 port map ( Y=>nx5717, A=>nx5921);
   ix5718 : inv01 port map ( Y=>nx5719, A=>nx5921);
   ix5720 : inv01 port map ( Y=>nx5721, A=>nx5921);
   ix5722 : inv01 port map ( Y=>nx5723, A=>nx5921);
   ix5724 : inv01 port map ( Y=>nx5725, A=>nx5923);
   ix5726 : inv01 port map ( Y=>nx5727, A=>nx5923);
   ix5728 : inv01 port map ( Y=>nx5729, A=>nx5923);
   ix5730 : inv01 port map ( Y=>nx5731, A=>nx5923);
   ix5732 : inv01 port map ( Y=>nx5733, A=>nx5923);
   ix5734 : inv01 port map ( Y=>nx5735, A=>nx5923);
   ix5736 : inv01 port map ( Y=>nx5737, A=>nx5923);
   ix5738 : inv01 port map ( Y=>nx5739, A=>nx5925);
   ix5740 : inv01 port map ( Y=>nx5741, A=>nx5925);
   ix5742 : inv01 port map ( Y=>nx5743, A=>nx5925);
   ix5744 : inv01 port map ( Y=>nx5745, A=>nx5925);
   ix5746 : inv01 port map ( Y=>nx5747, A=>nx5925);
   ix5748 : inv01 port map ( Y=>nx5749, A=>nx5925);
   ix5750 : inv01 port map ( Y=>nx5751, A=>nx5925);
   ix5752 : inv01 port map ( Y=>nx5753, A=>nx5927);
   ix5754 : inv01 port map ( Y=>nx5755, A=>nx5927);
   ix5756 : inv01 port map ( Y=>nx5757, A=>nx5927);
   ix5758 : inv01 port map ( Y=>nx5759, A=>nx5927);
   ix5760 : inv01 port map ( Y=>nx5761, A=>nx5927);
   ix5762 : inv01 port map ( Y=>nx5763, A=>nx5927);
   ix5764 : inv01 port map ( Y=>nx5765, A=>nx5927);
   ix5766 : inv01 port map ( Y=>nx5767, A=>nx5929);
   ix5768 : inv01 port map ( Y=>nx5769, A=>nx5929);
   ix5770 : inv01 port map ( Y=>nx5771, A=>nx5929);
   ix5772 : inv01 port map ( Y=>nx5773, A=>nx5929);
   ix5774 : inv01 port map ( Y=>nx5775, A=>nx5929);
   ix5776 : inv01 port map ( Y=>nx5777, A=>nx5929);
   ix5778 : inv01 port map ( Y=>nx5779, A=>nx5929);
   ix5780 : inv01 port map ( Y=>nx5781, A=>nx5653);
   ix5782 : inv01 port map ( Y=>nx5783, A=>dataFromRam2_447);
   ix5784 : inv01 port map ( Y=>nx5785, A=>nx5931);
   ix5786 : inv01 port map ( Y=>nx5787, A=>nx5931);
   ix5788 : inv01 port map ( Y=>nx5789, A=>nx5931);
   ix5790 : inv01 port map ( Y=>nx5791, A=>nx5931);
   ix5792 : inv01 port map ( Y=>nx5793, A=>nx5931);
   ix5794 : inv01 port map ( Y=>nx5795, A=>nx5931);
   ix5796 : inv01 port map ( Y=>nx5797, A=>nx5931);
   ix5798 : inv01 port map ( Y=>nx5799, A=>nx5933);
   ix5800 : inv01 port map ( Y=>nx5801, A=>nx5933);
   ix5802 : inv01 port map ( Y=>nx5803, A=>nx5933);
   ix5804 : inv01 port map ( Y=>nx5805, A=>nx5933);
   ix5806 : inv01 port map ( Y=>nx5807, A=>nx5933);
   ix5808 : inv01 port map ( Y=>nx5809, A=>nx5933);
   ix5810 : inv01 port map ( Y=>nx5811, A=>nx5933);
   ix5812 : inv01 port map ( Y=>nx5813, A=>nx5935);
   ix5814 : inv01 port map ( Y=>nx5815, A=>nx5935);
   ix5816 : inv01 port map ( Y=>nx5817, A=>nx5935);
   ix5818 : inv01 port map ( Y=>nx5819, A=>nx5935);
   ix5820 : inv01 port map ( Y=>nx5821, A=>nx5935);
   ix5822 : inv01 port map ( Y=>nx5823, A=>nx5935);
   ix5824 : inv01 port map ( Y=>nx5825, A=>nx5935);
   ix5826 : inv01 port map ( Y=>nx5827, A=>nx5937);
   ix5828 : inv01 port map ( Y=>nx5829, A=>nx5937);
   ix5830 : inv01 port map ( Y=>nx5831, A=>nx5937);
   ix5832 : inv01 port map ( Y=>nx5833, A=>nx5937);
   ix5834 : inv01 port map ( Y=>nx5835, A=>nx5937);
   ix5836 : inv01 port map ( Y=>nx5837, A=>nx5937);
   ix5838 : inv01 port map ( Y=>nx5839, A=>nx5937);
   ix5840 : inv01 port map ( Y=>nx5841, A=>nx5939);
   ix5842 : inv01 port map ( Y=>nx5843, A=>nx5939);
   ix5844 : inv01 port map ( Y=>nx5845, A=>nx5939);
   ix5846 : inv01 port map ( Y=>nx5847, A=>nx5939);
   ix5848 : inv01 port map ( Y=>nx5849, A=>nx5939);
   ix5850 : inv01 port map ( Y=>nx5851, A=>nx5939);
   ix5852 : inv01 port map ( Y=>nx5853, A=>nx5939);
   ix5854 : inv01 port map ( Y=>nx5855, A=>nx5941);
   ix5856 : inv01 port map ( Y=>nx5857, A=>nx5941);
   ix5858 : inv01 port map ( Y=>nx5859, A=>nx5941);
   ix5860 : inv01 port map ( Y=>nx5861, A=>nx5941);
   ix5862 : inv01 port map ( Y=>nx5863, A=>nx5941);
   ix5864 : inv01 port map ( Y=>nx5865, A=>nx5941);
   ix5866 : inv01 port map ( Y=>nx5867, A=>nx5941);
   ix5868 : inv01 port map ( Y=>nx5869, A=>nx5943);
   ix5870 : inv01 port map ( Y=>nx5871, A=>nx5943);
   ix5872 : inv01 port map ( Y=>nx5873, A=>nx5943);
   ix5874 : inv01 port map ( Y=>nx5875, A=>nx5943);
   ix5876 : inv01 port map ( Y=>nx5877, A=>nx5943);
   ix5878 : inv01 port map ( Y=>nx5879, A=>nx5943);
   ix5880 : inv01 port map ( Y=>nx5881, A=>nx5943);
   ix5882 : inv01 port map ( Y=>nx5883, A=>nx5945);
   ix5884 : inv01 port map ( Y=>nx5885, A=>nx5945);
   ix5886 : inv01 port map ( Y=>nx5887, A=>nx5945);
   ix5888 : inv01 port map ( Y=>nx5889, A=>nx5945);
   ix5890 : inv01 port map ( Y=>nx5891, A=>nx5945);
   ix5892 : inv01 port map ( Y=>nx5893, A=>nx5945);
   ix5894 : inv01 port map ( Y=>nx5895, A=>nx5945);
   ix5896 : inv01 port map ( Y=>nx5897, A=>nx5947);
   ix5898 : inv01 port map ( Y=>nx5899, A=>nx5947);
   ix5900 : inv01 port map ( Y=>nx5901, A=>nx5947);
   ix5902 : inv01 port map ( Y=>nx5903, A=>nx5947);
   ix5904 : inv01 port map ( Y=>nx5905, A=>nx5947);
   ix5906 : inv01 port map ( Y=>nx5907, A=>nx5947);
   ix5908 : inv01 port map ( Y=>nx5909, A=>nx5947);
   ix5910 : inv01 port map ( Y=>nx5911, A=>nx5783);
   ix5912 : inv01 port map ( Y=>nx5913, A=>nx5953);
   ix5914 : inv01 port map ( Y=>nx5915, A=>nx5953);
   ix5916 : inv01 port map ( Y=>nx5917, A=>nx5953);
   ix5918 : inv01 port map ( Y=>nx5919, A=>nx5953);
   ix5920 : inv01 port map ( Y=>nx5921, A=>nx5953);
   ix5922 : inv01 port map ( Y=>nx5923, A=>nx5953);
   ix5924 : inv01 port map ( Y=>nx5925, A=>nx5953);
   ix5926 : inv01 port map ( Y=>nx5927, A=>nx5955);
   ix5928 : inv01 port map ( Y=>nx5929, A=>nx5955);
   ix5930 : inv01 port map ( Y=>nx5931, A=>nx5957);
   ix5932 : inv01 port map ( Y=>nx5933, A=>nx5957);
   ix5934 : inv01 port map ( Y=>nx5935, A=>nx5957);
   ix5936 : inv01 port map ( Y=>nx5937, A=>nx5957);
   ix5938 : inv01 port map ( Y=>nx5939, A=>nx5957);
   ix5940 : inv01 port map ( Y=>nx5941, A=>nx5957);
   ix5942 : inv01 port map ( Y=>nx5943, A=>nx5957);
   ix5944 : inv01 port map ( Y=>nx5945, A=>nx5959);
   ix5946 : inv01 port map ( Y=>nx5947, A=>nx5959);
   ix5952 : inv01 port map ( Y=>nx5953, A=>nx5653);
   ix5954 : inv01 port map ( Y=>nx5955, A=>nx5653);
   ix5956 : inv01 port map ( Y=>nx5957, A=>nx5783);
   ix5958 : inv01 port map ( Y=>nx5959, A=>nx5783);
   ix13 : and02 port map ( Y=>ram1Write, A0=>test, A1=>writeEn);
   ix15 : nor02ii port map ( Y=>ram2Write, A0=>test, A1=>writeEn);
   ix19 : and02 port map ( Y=>ram1Read, A0=>test, A1=>readEn);
   ix21 : nor02ii port map ( Y=>ram2Read, A0=>test, A1=>readEn);
   ix9 : mux21_ni port map ( Y=>MFC, A0=>mfcOfRam2, A1=>mfcOfRam1, S0=>test
   );
end DMAmemory ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity nBitRegister_16 is
   port (
      D : IN std_logic_vector (15 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      EN : IN std_logic ;
      Q : OUT std_logic_vector (15 DOWNTO 0)) ;
end nBitRegister_16 ;

architecture Data_flow of nBitRegister_16 is
   signal Q_15_EXMPLR, Q_14_EXMPLR, Q_13_EXMPLR, Q_12_EXMPLR, Q_11_EXMPLR, 
      Q_10_EXMPLR, Q_9_EXMPLR, Q_8_EXMPLR, Q_7_EXMPLR, Q_6_EXMPLR, 
      Q_5_EXMPLR, Q_4_EXMPLR, Q_3_EXMPLR, Q_2_EXMPLR, Q_1_EXMPLR, Q_0_EXMPLR, 
      nx230, nx240, nx250, nx260, nx270, nx280, nx290, nx300, nx310, nx320, 
      nx330, nx340, nx350, nx360, nx370, nx380, nx445, nx447, nx449, nx455, 
      nx457, nx459, nx461: std_logic ;

begin
   Q(15) <= Q_15_EXMPLR ;
   Q(14) <= Q_14_EXMPLR ;
   Q(13) <= Q_13_EXMPLR ;
   Q(12) <= Q_12_EXMPLR ;
   Q(11) <= Q_11_EXMPLR ;
   Q(10) <= Q_10_EXMPLR ;
   Q(9) <= Q_9_EXMPLR ;
   Q(8) <= Q_8_EXMPLR ;
   Q(7) <= Q_7_EXMPLR ;
   Q(6) <= Q_6_EXMPLR ;
   Q(5) <= Q_5_EXMPLR ;
   Q(4) <= Q_4_EXMPLR ;
   Q(3) <= Q_3_EXMPLR ;
   Q(2) <= Q_2_EXMPLR ;
   Q(1) <= Q_1_EXMPLR ;
   Q(0) <= Q_0_EXMPLR ;
   reg_Q_0 : dffr port map ( Q=>Q_0_EXMPLR, QB=>OPEN, D=>nx230, CLK=>nx445, 
      R=>RST);
   ix231 : mux21_ni port map ( Y=>nx230, A0=>Q_0_EXMPLR, A1=>D(0), S0=>nx457
   );
   reg_Q_1 : dffr port map ( Q=>Q_1_EXMPLR, QB=>OPEN, D=>nx240, CLK=>nx445, 
      R=>RST);
   ix241 : mux21_ni port map ( Y=>nx240, A0=>Q_1_EXMPLR, A1=>D(1), S0=>nx457
   );
   reg_Q_2 : dffr port map ( Q=>Q_2_EXMPLR, QB=>OPEN, D=>nx250, CLK=>nx445, 
      R=>RST);
   ix251 : mux21_ni port map ( Y=>nx250, A0=>Q_2_EXMPLR, A1=>D(2), S0=>nx457
   );
   reg_Q_3 : dffr port map ( Q=>Q_3_EXMPLR, QB=>OPEN, D=>nx260, CLK=>nx445, 
      R=>RST);
   ix261 : mux21_ni port map ( Y=>nx260, A0=>Q_3_EXMPLR, A1=>D(3), S0=>nx457
   );
   reg_Q_4 : dffr port map ( Q=>Q_4_EXMPLR, QB=>OPEN, D=>nx270, CLK=>nx445, 
      R=>RST);
   ix271 : mux21_ni port map ( Y=>nx270, A0=>Q_4_EXMPLR, A1=>D(4), S0=>nx457
   );
   reg_Q_5 : dffr port map ( Q=>Q_5_EXMPLR, QB=>OPEN, D=>nx280, CLK=>nx445, 
      R=>RST);
   ix281 : mux21_ni port map ( Y=>nx280, A0=>Q_5_EXMPLR, A1=>D(5), S0=>nx457
   );
   reg_Q_6 : dffr port map ( Q=>Q_6_EXMPLR, QB=>OPEN, D=>nx290, CLK=>nx445, 
      R=>RST);
   ix291 : mux21_ni port map ( Y=>nx290, A0=>Q_6_EXMPLR, A1=>D(6), S0=>nx457
   );
   reg_Q_7 : dffr port map ( Q=>Q_7_EXMPLR, QB=>OPEN, D=>nx300, CLK=>nx447, 
      R=>RST);
   ix301 : mux21_ni port map ( Y=>nx300, A0=>Q_7_EXMPLR, A1=>D(7), S0=>nx459
   );
   reg_Q_8 : dffr port map ( Q=>Q_8_EXMPLR, QB=>OPEN, D=>nx310, CLK=>nx447, 
      R=>RST);
   ix311 : mux21_ni port map ( Y=>nx310, A0=>Q_8_EXMPLR, A1=>D(8), S0=>nx459
   );
   reg_Q_9 : dffr port map ( Q=>Q_9_EXMPLR, QB=>OPEN, D=>nx320, CLK=>nx447, 
      R=>RST);
   ix321 : mux21_ni port map ( Y=>nx320, A0=>Q_9_EXMPLR, A1=>D(9), S0=>nx459
   );
   reg_Q_10 : dffr port map ( Q=>Q_10_EXMPLR, QB=>OPEN, D=>nx330, CLK=>nx447, 
      R=>RST);
   ix331 : mux21_ni port map ( Y=>nx330, A0=>Q_10_EXMPLR, A1=>D(10), S0=>
      nx459);
   reg_Q_11 : dffr port map ( Q=>Q_11_EXMPLR, QB=>OPEN, D=>nx340, CLK=>nx447, 
      R=>RST);
   ix341 : mux21_ni port map ( Y=>nx340, A0=>Q_11_EXMPLR, A1=>D(11), S0=>
      nx459);
   reg_Q_12 : dffr port map ( Q=>Q_12_EXMPLR, QB=>OPEN, D=>nx350, CLK=>nx447, 
      R=>RST);
   ix351 : mux21_ni port map ( Y=>nx350, A0=>Q_12_EXMPLR, A1=>D(12), S0=>
      nx459);
   reg_Q_13 : dffr port map ( Q=>Q_13_EXMPLR, QB=>OPEN, D=>nx360, CLK=>nx447, 
      R=>RST);
   ix361 : mux21_ni port map ( Y=>nx360, A0=>Q_13_EXMPLR, A1=>D(13), S0=>
      nx459);
   reg_Q_14 : dffr port map ( Q=>Q_14_EXMPLR, QB=>OPEN, D=>nx370, CLK=>nx449, 
      R=>RST);
   ix371 : mux21_ni port map ( Y=>nx370, A0=>Q_14_EXMPLR, A1=>D(14), S0=>
      nx461);
   reg_Q_15 : dffr port map ( Q=>Q_15_EXMPLR, QB=>OPEN, D=>nx380, CLK=>nx449, 
      R=>RST);
   ix381 : mux21_ni port map ( Y=>nx380, A0=>Q_15_EXMPLR, A1=>D(15), S0=>
      nx461);
   ix444 : inv02 port map ( Y=>nx445, A=>CLK);
   ix446 : inv02 port map ( Y=>nx447, A=>CLK);
   ix448 : inv02 port map ( Y=>nx449, A=>CLK);
   ix454 : inv01 port map ( Y=>nx455, A=>EN);
   ix456 : inv02 port map ( Y=>nx457, A=>nx455);
   ix458 : inv02 port map ( Y=>nx459, A=>nx455);
   ix460 : inv02 port map ( Y=>nx461, A=>nx455);
end Data_flow ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity ReadInfoState is
   port (
      CLK : IN std_logic ;
      S : IN std_logic_vector (14 DOWNTO 0) ;
      reset : IN std_logic ;
      MFC : IN std_logic ;
      filterAddressReg_out : IN std_logic_vector (12 DOWNTO 0) ;
      filterRamData : IN std_logic_vector (15 DOWNTO 0) ;
      noOfLayersReg_out : OUT std_logic_vector (15 DOWNTO 0) ;
      filterRamAddress : OUT std_logic_vector (12 DOWNTO 0)) ;
end ReadInfoState ;

architecture archReadInfoState of ReadInfoState is
   component nBitRegister_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
begin
   noOfLayersReg : nBitRegister_16 port map ( D(15)=>filterRamData(15), 
      D(14)=>filterRamData(14), D(13)=>filterRamData(13), D(12)=>
      filterRamData(12), D(11)=>filterRamData(11), D(10)=>filterRamData(10), 
      D(9)=>filterRamData(9), D(8)=>filterRamData(8), D(7)=>filterRamData(7), 
      D(6)=>filterRamData(6), D(5)=>filterRamData(5), D(4)=>filterRamData(4), 
      D(3)=>filterRamData(3), D(2)=>filterRamData(2), D(1)=>filterRamData(1), 
      D(0)=>filterRamData(0), CLK=>CLK, RST=>reset, EN=>S(0), Q(15)=>
      noOfLayersReg_out(15), Q(14)=>noOfLayersReg_out(14), Q(13)=>
      noOfLayersReg_out(13), Q(12)=>noOfLayersReg_out(12), Q(11)=>
      noOfLayersReg_out(11), Q(10)=>noOfLayersReg_out(10), Q(9)=>
      noOfLayersReg_out(9), Q(8)=>noOfLayersReg_out(8), Q(7)=>
      noOfLayersReg_out(7), Q(6)=>noOfLayersReg_out(6), Q(5)=>
      noOfLayersReg_out(5), Q(4)=>noOfLayersReg_out(4), Q(3)=>
      noOfLayersReg_out(3), Q(2)=>noOfLayersReg_out(2), Q(1)=>
      noOfLayersReg_out(1), Q(0)=>noOfLayersReg_out(0));
   dmaOut : triStateBuffer_13 port map ( D(12)=>filterAddressReg_out(12), 
      D(11)=>filterAddressReg_out(11), D(10)=>filterAddressReg_out(10), D(9)
      =>filterAddressReg_out(9), D(8)=>filterAddressReg_out(8), D(7)=>
      filterAddressReg_out(7), D(6)=>filterAddressReg_out(6), D(5)=>
      filterAddressReg_out(5), D(4)=>filterAddressReg_out(4), D(3)=>
      filterAddressReg_out(3), D(2)=>filterAddressReg_out(2), D(1)=>
      filterAddressReg_out(1), D(0)=>filterAddressReg_out(0), EN=>S(0), 
      F(12)=>filterRamAddress(12), F(11)=>filterRamAddress(11), F(10)=>
      filterRamAddress(10), F(9)=>filterRamAddress(9), F(8)=>
      filterRamAddress(8), F(7)=>filterRamAddress(7), F(6)=>
      filterRamAddress(6), F(5)=>filterRamAddress(5), F(4)=>
      filterRamAddress(4), F(3)=>filterRamAddress(3), F(2)=>
      filterRamAddress(2), F(1)=>filterRamAddress(1), F(0)=>
      filterRamAddress(0));
end archReadInfoState ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity my_adder is
   port (
      a : IN std_logic ;
      b : IN std_logic ;
      cin : IN std_logic ;
      s : OUT std_logic ;
      cout : OUT std_logic) ;
end my_adder ;

architecture a_my_adder of my_adder is
   signal nx0, nx69: std_logic ;

begin
   ix7 : ao22 port map ( Y=>cout, A0=>b, A1=>a, B0=>cin, B1=>nx0);
   ix9 : xnor2 port map ( Y=>s, A0=>nx69, A1=>cin);
   ix70 : xnor2 port map ( Y=>nx69, A0=>a, A1=>b);
   ix1 : inv01 port map ( Y=>nx0, A=>nx69);
end a_my_adder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity my_nadder_13 is
   port (
      a : IN std_logic_vector (12 DOWNTO 0) ;
      b : IN std_logic_vector (12 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (12 DOWNTO 0) ;
      cout : OUT std_logic) ;
end my_nadder_13 ;

architecture a_my_nadder of my_nadder_13 is
   component my_adder
      port (
         a : IN std_logic ;
         b : IN std_logic ;
         cin : IN std_logic ;
         s : OUT std_logic ;
         cout : OUT std_logic) ;
   end component ;
   signal temp_11, temp_10, temp_9, temp_8, temp_7, temp_6, temp_5, temp_4, 
      temp_3, temp_2, temp_1, temp_0: std_logic ;

begin
   f0 : my_adder port map ( a=>a(0), b=>b(0), cin=>cin, s=>s(0), cout=>
      temp_0);
   loop1_1_fx : my_adder port map ( a=>a(1), b=>b(1), cin=>temp_0, s=>s(1), 
      cout=>temp_1);
   loop1_2_fx : my_adder port map ( a=>a(2), b=>b(2), cin=>temp_1, s=>s(2), 
      cout=>temp_2);
   loop1_3_fx : my_adder port map ( a=>a(3), b=>b(3), cin=>temp_2, s=>s(3), 
      cout=>temp_3);
   loop1_4_fx : my_adder port map ( a=>a(4), b=>b(4), cin=>temp_3, s=>s(4), 
      cout=>temp_4);
   loop1_5_fx : my_adder port map ( a=>a(5), b=>b(5), cin=>temp_4, s=>s(5), 
      cout=>temp_5);
   loop1_6_fx : my_adder port map ( a=>a(6), b=>b(6), cin=>temp_5, s=>s(6), 
      cout=>temp_6);
   loop1_7_fx : my_adder port map ( a=>a(7), b=>b(7), cin=>temp_6, s=>s(7), 
      cout=>temp_7);
   loop1_8_fx : my_adder port map ( a=>a(8), b=>b(8), cin=>temp_7, s=>s(8), 
      cout=>temp_8);
   loop1_9_fx : my_adder port map ( a=>a(9), b=>b(9), cin=>temp_8, s=>s(9), 
      cout=>temp_9);
   loop1_10_fx : my_adder port map ( a=>a(10), b=>b(10), cin=>temp_9, s=>
      s(10), cout=>temp_10);
   loop1_11_fx : my_adder port map ( a=>a(11), b=>b(11), cin=>temp_10, s=>
      s(11), cout=>temp_11);
   loop1_12_fx : my_adder port map ( a=>a(12), b=>b(12), cin=>temp_11, s=>
      s(12), cout=>cout);
end a_my_nadder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity ReadLayerInfo is
   port (
      LayerInfoIn : IN std_logic_vector (15 DOWNTO 0) ;
      ImgWidthIn : IN std_logic_vector (15 DOWNTO 0) ;
      FilterAdd : IN std_logic_vector (12 DOWNTO 0) ;
      ImgAdd : IN std_logic_vector (12 DOWNTO 0) ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      ACKF : IN std_logic ;
      ACKI : IN std_logic ;
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      LayerInfoOut : OUT std_logic_vector (15 DOWNTO 0) ;
      ImgWidthOut : OUT std_logic_vector (15 DOWNTO 0) ;
      FilterAddToDMA : OUT std_logic_vector (12 DOWNTO 0) ;
      ImgAddToDMA : OUT std_logic_vector (12 DOWNTO 0)) ;
end ReadLayerInfo ;

architecture LayerInfo of ReadLayerInfo is
   component nBitRegister_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   signal LayerInfEN, ImgWidthEN: std_logic ;

begin
   LayerInf : nBitRegister_16 port map ( D(15)=>LayerInfoIn(15), D(14)=>
      LayerInfoIn(14), D(13)=>LayerInfoIn(13), D(12)=>LayerInfoIn(12), D(11)
      =>LayerInfoIn(11), D(10)=>LayerInfoIn(10), D(9)=>LayerInfoIn(9), D(8)
      =>LayerInfoIn(8), D(7)=>LayerInfoIn(7), D(6)=>LayerInfoIn(6), D(5)=>
      LayerInfoIn(5), D(4)=>LayerInfoIn(4), D(3)=>LayerInfoIn(3), D(2)=>
      LayerInfoIn(2), D(1)=>LayerInfoIn(1), D(0)=>LayerInfoIn(0), CLK=>clk, 
      RST=>rst, EN=>LayerInfEN, Q(15)=>LayerInfoOut(15), Q(14)=>
      LayerInfoOut(14), Q(13)=>LayerInfoOut(13), Q(12)=>LayerInfoOut(12), 
      Q(11)=>LayerInfoOut(11), Q(10)=>LayerInfoOut(10), Q(9)=>
      LayerInfoOut(9), Q(8)=>LayerInfoOut(8), Q(7)=>LayerInfoOut(7), Q(6)=>
      LayerInfoOut(6), Q(5)=>LayerInfoOut(5), Q(4)=>LayerInfoOut(4), Q(3)=>
      LayerInfoOut(3), Q(2)=>LayerInfoOut(2), Q(1)=>LayerInfoOut(1), Q(0)=>
      LayerInfoOut(0));
   ImgWidth : nBitRegister_16 port map ( D(15)=>ImgWidthIn(15), D(14)=>
      ImgWidthIn(14), D(13)=>ImgWidthIn(13), D(12)=>ImgWidthIn(12), D(11)=>
      ImgWidthIn(11), D(10)=>ImgWidthIn(10), D(9)=>ImgWidthIn(9), D(8)=>
      ImgWidthIn(8), D(7)=>ImgWidthIn(7), D(6)=>ImgWidthIn(6), D(5)=>
      ImgWidthIn(5), D(4)=>ImgWidthIn(4), D(3)=>ImgWidthIn(3), D(2)=>
      ImgWidthIn(2), D(1)=>ImgWidthIn(1), D(0)=>ImgWidthIn(0), CLK=>clk, RST
      =>rst, EN=>ImgWidthEN, Q(15)=>ImgWidthOut(15), Q(14)=>ImgWidthOut(14), 
      Q(13)=>ImgWidthOut(13), Q(12)=>ImgWidthOut(12), Q(11)=>ImgWidthOut(11), 
      Q(10)=>ImgWidthOut(10), Q(9)=>ImgWidthOut(9), Q(8)=>ImgWidthOut(8), 
      Q(7)=>ImgWidthOut(7), Q(6)=>ImgWidthOut(6), Q(5)=>ImgWidthOut(5), Q(4)
      =>ImgWidthOut(4), Q(3)=>ImgWidthOut(3), Q(2)=>ImgWidthOut(2), Q(1)=>
      ImgWidthOut(1), Q(0)=>ImgWidthOut(0));
   FilterAddTriDMA : triStateBuffer_13 port map ( D(12)=>FilterAdd(12), 
      D(11)=>FilterAdd(11), D(10)=>FilterAdd(10), D(9)=>FilterAdd(9), D(8)=>
      FilterAdd(8), D(7)=>FilterAdd(7), D(6)=>FilterAdd(6), D(5)=>
      FilterAdd(5), D(4)=>FilterAdd(4), D(3)=>FilterAdd(3), D(2)=>
      FilterAdd(2), D(1)=>FilterAdd(1), D(0)=>FilterAdd(0), EN=>
      current_state(1), F(12)=>FilterAddToDMA(12), F(11)=>FilterAddToDMA(11), 
      F(10)=>FilterAddToDMA(10), F(9)=>FilterAddToDMA(9), F(8)=>
      FilterAddToDMA(8), F(7)=>FilterAddToDMA(7), F(6)=>FilterAddToDMA(6), 
      F(5)=>FilterAddToDMA(5), F(4)=>FilterAddToDMA(4), F(3)=>
      FilterAddToDMA(3), F(2)=>FilterAddToDMA(2), F(1)=>FilterAddToDMA(1), 
      F(0)=>FilterAddToDMA(0));
   ImgAddTriDMA : triStateBuffer_13 port map ( D(12)=>ImgAdd(12), D(11)=>
      ImgAdd(11), D(10)=>ImgAdd(10), D(9)=>ImgAdd(9), D(8)=>ImgAdd(8), D(7)
      =>ImgAdd(7), D(6)=>ImgAdd(6), D(5)=>ImgAdd(5), D(4)=>ImgAdd(4), D(3)=>
      ImgAdd(3), D(2)=>ImgAdd(2), D(1)=>ImgAdd(1), D(0)=>ImgAdd(0), EN=>
      current_state(1), F(12)=>ImgAddToDMA(12), F(11)=>ImgAddToDMA(11), 
      F(10)=>ImgAddToDMA(10), F(9)=>ImgAddToDMA(9), F(8)=>ImgAddToDMA(8), 
      F(7)=>ImgAddToDMA(7), F(6)=>ImgAddToDMA(6), F(5)=>ImgAddToDMA(5), F(4)
      =>ImgAddToDMA(4), F(3)=>ImgAddToDMA(3), F(2)=>ImgAddToDMA(2), F(1)=>
      ImgAddToDMA(1), F(0)=>ImgAddToDMA(0));
   ix1 : and02 port map ( Y=>ImgWidthEN, A0=>ACKI, A1=>current_state(1));
   ix3 : and02 port map ( Y=>LayerInfEN, A0=>ACKF, A1=>current_state(1));

end LayerInfo ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity my_nadder_5 is
   port (
      a : IN std_logic_vector (4 DOWNTO 0) ;
      b : IN std_logic_vector (4 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (4 DOWNTO 0) ;
      cout : OUT std_logic) ;
end my_nadder_5 ;

architecture a_my_nadder of my_nadder_5 is
   component my_adder
      port (
         a : IN std_logic ;
         b : IN std_logic ;
         cin : IN std_logic ;
         s : OUT std_logic ;
         cout : OUT std_logic) ;
   end component ;
   signal temp_3, temp_2, temp_1, temp_0: std_logic ;

begin
   f0 : my_adder port map ( a=>a(0), b=>b(0), cin=>cin, s=>s(0), cout=>
      temp_0);
   loop1_1_fx : my_adder port map ( a=>a(1), b=>b(1), cin=>temp_0, s=>s(1), 
      cout=>temp_1);
   loop1_2_fx : my_adder port map ( a=>a(2), b=>b(2), cin=>temp_1, s=>s(2), 
      cout=>temp_2);
   loop1_3_fx : my_adder port map ( a=>a(3), b=>b(3), cin=>temp_2, s=>s(3), 
      cout=>temp_3);
   loop1_4_fx : my_adder port map ( a=>a(4), b=>b(4), cin=>temp_3, s=>s(4), 
      cout=>cout);
end a_my_nadder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity my_nadder_2 is
   port (
      a : IN std_logic_vector (1 DOWNTO 0) ;
      b : IN std_logic_vector (1 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (1 DOWNTO 0) ;
      cout : OUT std_logic) ;
end my_nadder_2 ;

architecture a_my_nadder of my_nadder_2 is
   component my_adder
      port (
         a : IN std_logic ;
         b : IN std_logic ;
         cin : IN std_logic ;
         s : OUT std_logic ;
         cout : OUT std_logic) ;
   end component ;
   signal temp_0: std_logic ;

begin
   f0 : my_adder port map ( a=>a(0), b=>b(0), cin=>cin, s=>s(0), cout=>
      temp_0);
   loop1_1_fx : my_adder port map ( a=>a(1), b=>b(1), cin=>temp_0, s=>s(1), 
      cout=>cout);
end a_my_nadder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Counter_2 is
   port (
      enable : IN std_logic ;
      reset : IN std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      output : OUT std_logic_vector (1 DOWNTO 0) ;
      input : IN std_logic_vector (1 DOWNTO 0)) ;
end Counter_2 ;

architecture CounterImplementation of Counter_2 is
   component my_nadder_2
      port (
         a : IN std_logic_vector (1 DOWNTO 0) ;
         b : IN std_logic_vector (1 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (1 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal output_1_EXMPLR, output_0_EXMPLR, addResult_1, addResult_0, one_0, 
      one_1, nx28, NOT_clk, nx8, nx12, nx22, nx20, nx25, nx85, nx95, nx104: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   output(1) <= output_1_EXMPLR ;
   output(0) <= output_0_EXMPLR ;
   A1 : my_nadder_2 port map ( a(1)=>output_1_EXMPLR, a(0)=>output_0_EXMPLR, 
      b(1)=>one_1, b(0)=>one_0, cin=>one_1, s(1)=>addResult_1, s(0)=>
      addResult_0, cout=>DANGLING(0));
   ix68 : fake_gnd port map ( Y=>one_1);
   ix66 : fake_vcc port map ( Y=>one_0);
   reg_toOutput_0_dup_1 : dffsr_ni port map ( Q=>output_0_EXMPLR, QB=>OPEN, 
      D=>nx85, CLK=>clk, S=>nx8, R=>nx12);
   ix86 : mux21_ni port map ( Y=>nx85, A0=>output_0_EXMPLR, A1=>addResult_0, 
      S0=>enable);
   ix9 : nor02ii port map ( Y=>nx8, A0=>nx104, A1=>nx28);
   ix105 : nor02_2x port map ( Y=>nx104, A0=>reset, A1=>load);
   ix29 : dffr port map ( Q=>nx28, QB=>OPEN, D=>input(0), CLK=>NOT_clk, R=>
      reset);
   ix108 : inv01 port map ( Y=>NOT_clk, A=>clk);
   ix13 : nor02_2x port map ( Y=>nx12, A0=>nx28, A1=>nx104);
   reg_toOutput_1_dup_1 : dffsr_ni port map ( Q=>output_1_EXMPLR, QB=>OPEN, 
      D=>nx95, CLK=>clk, S=>nx20, R=>nx25);
   ix96 : mux21_ni port map ( Y=>nx95, A0=>output_1_EXMPLR, A1=>addResult_1, 
      S0=>enable);
   ix21 : nor02ii port map ( Y=>nx20, A0=>nx104, A1=>nx22);
   ix23 : dffr port map ( Q=>nx22, QB=>OPEN, D=>input(1), CLK=>NOT_clk, R=>
      reset);
   ix26 : nor02_2x port map ( Y=>nx25, A0=>nx22, A1=>nx104);
end CounterImplementation ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity CalculateInfo is
   port (
      WSquareOut : OUT std_logic_vector (9 DOWNTO 0) ;
      CounOut : OUT std_logic_vector (1 DOWNTO 0) ;
      LayerInfoIn : IN std_logic_vector (15 DOWNTO 0) ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      ACK : OUT std_logic ;
      ACKI : IN std_logic ;
      Wmin1 : OUT std_logic_vector (4 DOWNTO 0)) ;
end CalculateInfo ;

architecture CalInfo of CalculateInfo is
   component my_nadder_5
      port (
         a : IN std_logic_vector (4 DOWNTO 0) ;
         b : IN std_logic_vector (4 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (4 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component Counter_2
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (1 DOWNTO 0) ;
         input : IN std_logic_vector (1 DOWNTO 0)) ;
   end component ;
   signal WSquareOut_0_EXMPLR, CounOut_1_EXMPLR, CounOut_0_EXMPLR, 
      ACK_EXMPLR, Wmin1_4_EXMPLR, Wmin1_3_EXMPLR, Wmin1_2_EXMPLR, 
      Wmin1_1_EXMPLR, Wmin1_0_EXMPLR, CountereEN, CountereRST, GND0, PWR, 
      nx0, nx2, nx12, nx38, nx42, nx46, nx48, nx54, nx58, nx60, nx86, nx88, 
      nx110, nx116, nx130, nx132, nx146, nx148, nx172, nx180, nx182, nx190, 
      nx192, nx206, nx208, nx232, nx236, nx240, nx274, nx290, nx111, nx123, 
      nx129, nx131, nx139, nx141, nx143, nx147, nx157, nx159, nx161, nx163, 
      nx167, nx173, nx183, nx185, nx187, nx189, nx191, nx195, nx197, nx199, 
      nx201, nx203, nx205, nx207, nx209, nx211, nx213, nx215, nx217, nx219, 
      nx227, nx231, nx239, nx241, nx243, nx245, nx247, nx255, nx263, nx265, 
      nx267, nx279, nx291, nx293, nx295, nx297: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   WSquareOut(0) <= WSquareOut_0_EXMPLR ;
   CounOut(1) <= CounOut_1_EXMPLR ;
   CounOut(0) <= CounOut_0_EXMPLR ;
   ACK <= ACK_EXMPLR ;
   Wmin1(4) <= Wmin1_4_EXMPLR ;
   Wmin1(3) <= Wmin1_3_EXMPLR ;
   Wmin1(2) <= Wmin1_2_EXMPLR ;
   Wmin1(1) <= Wmin1_1_EXMPLR ;
   Wmin1(0) <= Wmin1_0_EXMPLR ;
   adder : my_nadder_5 port map ( a(4)=>LayerInfoIn(8), a(3)=>LayerInfoIn(7), 
      a(2)=>LayerInfoIn(6), a(1)=>nx291, a(0)=>nx295, b(4)=>PWR, b(3)=>PWR, 
      b(2)=>PWR, b(1)=>PWR, b(0)=>PWR, cin=>GND0, s(4)=>Wmin1_4_EXMPLR, s(3)
      =>Wmin1_3_EXMPLR, s(2)=>Wmin1_2_EXMPLR, s(1)=>Wmin1_1_EXMPLR, s(0)=>
      Wmin1_0_EXMPLR, cout=>DANGLING(0));
   EndCounter : Counter_2 port map ( enable=>CountereEN, reset=>CountereRST, 
      clk=>clk, load=>GND0, output(1)=>CounOut_1_EXMPLR, output(0)=>
      CounOut_0_EXMPLR, input(1)=>GND0, input(0)=>GND0);
   ix81 : fake_vcc port map ( Y=>PWR);
   ix79 : fake_gnd port map ( Y=>GND0);
   ix285 : ao221 port map ( Y=>CountereRST, A0=>CounOut_1_EXMPLR, A1=>nx111, 
      B0=>ACKI, B1=>nx274, C0=>rst);
   ix112 : inv01 port map ( Y=>nx111, A=>CounOut_0_EXMPLR);
   ix275 : or02 port map ( Y=>nx274, A0=>current_state(2), A1=>
      current_state(4));
   ix301 : nor02_2x port map ( Y=>CountereEN, A0=>ACK_EXMPLR, A1=>nx123);
   reg_ACKW_dup_1 : dffs_ni port map ( Q=>ACK_EXMPLR, QB=>OPEN, D=>GND0, CLK
      =>clk, S=>nx290);
   ix291 : nor02ii port map ( Y=>nx290, A0=>CounOut_1_EXMPLR, A1=>
      CounOut_0_EXMPLR);
   ix124 : nor02_2x port map ( Y=>nx123, A0=>current_state(2), A1=>
      current_state(4));
   ix215 : and02 port map ( Y=>WSquareOut_0_EXMPLR, A0=>Wmin1_0_EXMPLR, A1=>
      nx295);
   ix273 : nor02ii port map ( Y=>WSquareOut(1), A0=>nx129, A1=>nx131);
   ix130 : aoi22 port map ( Y=>nx129, A0=>nx291, A1=>Wmin1_0_EXMPLR, B0=>
      Wmin1_1_EXMPLR, B1=>nx295);
   ix132 : nand03 port map ( Y=>nx131, A0=>WSquareOut_0_EXMPLR, A1=>nx291, 
      A2=>Wmin1_1_EXMPLR);
   ix263 : xnor2 port map ( Y=>WSquareOut(2), A0=>nx131, A1=>nx208);
   ix209 : xnor2 port map ( Y=>nx208, A0=>nx206, A1=>nx143);
   ix207 : nor02ii port map ( Y=>nx206, A0=>nx139, A1=>nx141);
   ix140 : aoi22 port map ( Y=>nx139, A0=>Wmin1_2_EXMPLR, A1=>nx295, B0=>
      nx291, B1=>Wmin1_1_EXMPLR);
   ix142 : nand04 port map ( Y=>nx141, A0=>nx291, A1=>Wmin1_1_EXMPLR, A2=>
      Wmin1_2_EXMPLR, A3=>nx295);
   ix144 : nand02 port map ( Y=>nx143, A0=>LayerInfoIn(6), A1=>
      Wmin1_0_EXMPLR);
   ix261 : xnor2 port map ( Y=>WSquareOut(3), A0=>nx147, A1=>nx192);
   ix148 : mux21_ni port map ( Y=>nx147, A0=>nx143, A1=>nx131, S0=>nx208);
   ix193 : xnor2 port map ( Y=>nx192, A0=>nx190, A1=>nx163);
   ix191 : xnor2 port map ( Y=>nx190, A0=>nx141, A1=>nx148);
   ix149 : xnor2 port map ( Y=>nx148, A0=>nx146, A1=>nx161);
   ix147 : nor02ii port map ( Y=>nx146, A0=>nx157, A1=>nx159);
   ix158 : aoi22 port map ( Y=>nx157, A0=>nx291, A1=>Wmin1_2_EXMPLR, B0=>
      Wmin1_3_EXMPLR, B1=>nx295);
   ix160 : nand04 port map ( Y=>nx159, A0=>Wmin1_3_EXMPLR, A1=>nx297, A2=>
      nx293, A3=>Wmin1_2_EXMPLR);
   ix162 : nand02 port map ( Y=>nx161, A0=>LayerInfoIn(6), A1=>
      Wmin1_1_EXMPLR);
   ix164 : nand02 port map ( Y=>nx163, A0=>LayerInfoIn(7), A1=>
      Wmin1_0_EXMPLR);
   ix259 : xnor2 port map ( Y=>WSquareOut(4), A0=>nx167, A1=>nx182);
   ix168 : mux21_ni port map ( Y=>nx167, A0=>nx163, A1=>nx147, S0=>nx192);
   ix183 : xnor2 port map ( Y=>nx182, A0=>nx180, A1=>nx191);
   ix181 : xnor2 port map ( Y=>nx180, A0=>nx173, A1=>nx132);
   ix174 : mux21_ni port map ( Y=>nx173, A0=>nx161, A1=>nx141, S0=>nx148);
   ix133 : xnor2 port map ( Y=>nx132, A0=>nx130, A1=>nx189);
   ix131 : xnor2 port map ( Y=>nx130, A0=>nx159, A1=>nx88);
   ix89 : xnor2 port map ( Y=>nx88, A0=>nx86, A1=>nx187);
   ix87 : nor02ii port map ( Y=>nx86, A0=>nx183, A1=>nx185);
   ix184 : aoi22 port map ( Y=>nx183, A0=>nx293, A1=>Wmin1_3_EXMPLR, B0=>
      Wmin1_4_EXMPLR, B1=>nx297);
   ix186 : nand04 port map ( Y=>nx185, A0=>nx293, A1=>Wmin1_4_EXMPLR, A2=>
      Wmin1_3_EXMPLR, A3=>nx297);
   ix188 : nand02 port map ( Y=>nx187, A0=>LayerInfoIn(6), A1=>
      Wmin1_2_EXMPLR);
   ix190 : nand02 port map ( Y=>nx189, A0=>LayerInfoIn(7), A1=>
      Wmin1_1_EXMPLR);
   ix192 : nand02 port map ( Y=>nx191, A0=>LayerInfoIn(8), A1=>
      Wmin1_0_EXMPLR);
   ix257 : xor2 port map ( Y=>WSquareOut(5), A0=>nx195, A1=>nx197);
   ix196 : mux21_ni port map ( Y=>nx195, A0=>nx191, A1=>nx167, S0=>nx182);
   ix198 : xnor2 port map ( Y=>nx197, A0=>nx199, A1=>nx201);
   ix200 : mux21_ni port map ( Y=>nx199, A0=>nx189, A1=>nx173, S0=>nx132);
   ix202 : xnor2 port map ( Y=>nx201, A0=>nx203, A1=>nx219);
   ix204 : xnor2 port map ( Y=>nx203, A0=>nx205, A1=>nx207);
   ix206 : mux21_ni port map ( Y=>nx205, A0=>nx187, A1=>nx159, S0=>nx88);
   ix208 : xnor2 port map ( Y=>nx207, A0=>nx209, A1=>nx217);
   ix210 : xnor2 port map ( Y=>nx209, A0=>nx185, A1=>nx211);
   ix212 : xnor2 port map ( Y=>nx211, A0=>nx213, A1=>nx215);
   ix214 : nand02 port map ( Y=>nx213, A0=>nx293, A1=>Wmin1_4_EXMPLR);
   ix216 : nand02 port map ( Y=>nx215, A0=>LayerInfoIn(6), A1=>
      Wmin1_3_EXMPLR);
   ix218 : nand02 port map ( Y=>nx217, A0=>LayerInfoIn(7), A1=>
      Wmin1_2_EXMPLR);
   ix220 : nand02 port map ( Y=>nx219, A0=>LayerInfoIn(8), A1=>
      Wmin1_1_EXMPLR);
   ix251 : xor2 port map ( Y=>WSquareOut(6), A0=>nx232, A1=>nx172);
   ix233 : nor02_2x port map ( Y=>nx232, A0=>nx195, A1=>nx197);
   ix173 : xnor2 port map ( Y=>nx172, A0=>nx227, A1=>nx116);
   ix228 : mux21_ni port map ( Y=>nx227, A0=>nx199, A1=>nx219, S0=>nx201);
   ix117 : xnor2 port map ( Y=>nx116, A0=>nx231, A1=>nx60);
   ix232 : mux21_ni port map ( Y=>nx231, A0=>nx205, A1=>nx217, S0=>nx207);
   ix61 : xnor2 port map ( Y=>nx60, A0=>nx58, A1=>nx247);
   ix59 : xnor2 port map ( Y=>nx58, A0=>nx38, A1=>nx241);
   ix39 : aoi21 port map ( Y=>nx38, A0=>nx239, A1=>nx215, B0=>nx213);
   ix240 : nand02 port map ( Y=>nx239, A0=>Wmin1_3_EXMPLR, A1=>nx297);
   ix242 : xnor2 port map ( Y=>nx241, A0=>nx243, A1=>nx245);
   ix244 : nand02 port map ( Y=>nx243, A0=>LayerInfoIn(6), A1=>
      Wmin1_4_EXMPLR);
   ix246 : nand02 port map ( Y=>nx245, A0=>LayerInfoIn(7), A1=>
      Wmin1_3_EXMPLR);
   ix248 : nand02 port map ( Y=>nx247, A0=>LayerInfoIn(8), A1=>
      Wmin1_2_EXMPLR);
   ix249 : xor2 port map ( Y=>WSquareOut(7), A0=>nx236, A1=>nx110);
   ix237 : mux21_ni port map ( Y=>nx236, A0=>nx116, A1=>nx232, S0=>nx172);
   ix111 : xnor2 port map ( Y=>nx110, A0=>nx255, A1=>nx54);
   ix256 : mux21_ni port map ( Y=>nx255, A0=>nx247, A1=>nx231, S0=>nx60);
   ix55 : xnor2 port map ( Y=>nx54, A0=>nx42, A1=>nx263);
   ix43 : mux21_ni port map ( Y=>nx42, A0=>nx38, A1=>nx12, S0=>nx241);
   ix264 : xnor2 port map ( Y=>nx263, A0=>nx265, A1=>nx267);
   ix266 : nand02 port map ( Y=>nx265, A0=>LayerInfoIn(7), A1=>
      Wmin1_4_EXMPLR);
   ix268 : nand02 port map ( Y=>nx267, A0=>LayerInfoIn(8), A1=>
      Wmin1_3_EXMPLR);
   ix247 : xor2 port map ( Y=>WSquareOut(8), A0=>nx240, A1=>nx48);
   ix241 : mux21_ni port map ( Y=>nx240, A0=>nx54, A1=>nx236, S0=>nx110);
   ix49 : xnor2 port map ( Y=>nx48, A0=>nx46, A1=>nx279);
   ix47 : mux21_ni port map ( Y=>nx46, A0=>nx42, A1=>nx2, S0=>nx263);
   ix280 : nand02 port map ( Y=>nx279, A0=>LayerInfoIn(8), A1=>
      Wmin1_4_EXMPLR);
   ix245 : mux21_ni port map ( Y=>WSquareOut(9), A0=>nx0, A1=>nx240, S0=>
      nx48);
   ix13 : inv01 port map ( Y=>nx12, A=>nx245);
   ix3 : inv01 port map ( Y=>nx2, A=>nx267);
   ix1 : inv01 port map ( Y=>nx0, A=>nx279);
   ix289 : buf02 port map ( Y=>nx291, A=>LayerInfoIn(5));
   ix292 : buf02 port map ( Y=>nx293, A=>LayerInfoIn(5));
   ix294 : buf02 port map ( Y=>nx295, A=>LayerInfoIn(4));
   ix296 : buf02 port map ( Y=>nx297, A=>LayerInfoIn(4));
end CalInfo ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity ReadBias is
   port (
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      BIAS : IN std_logic_vector (399 DOWNTO 0) ;
      FilterAddress : IN std_logic_vector (12 DOWNTO 0) ;
      DMAAddressToFilter : OUT std_logic_vector (12 DOWNTO 0) ;
      UpdatedAddress : OUT std_logic_vector (12 DOWNTO 0) ;
      changerAdd : OUT std_logic_vector (12 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
      outBias0 : OUT std_logic_vector (15 DOWNTO 0) ;
      outBias1 : OUT std_logic_vector (15 DOWNTO 0) ;
      outBias2 : OUT std_logic_vector (15 DOWNTO 0) ;
      outBias3 : OUT std_logic_vector (15 DOWNTO 0) ;
      outBias4 : OUT std_logic_vector (15 DOWNTO 0) ;
      outBias5 : OUT std_logic_vector (15 DOWNTO 0) ;
      outBias6 : OUT std_logic_vector (15 DOWNTO 0) ;
      outBias7 : OUT std_logic_vector (15 DOWNTO 0) ;
      ACKF : IN std_logic) ;
end ReadBias ;

architecture DATA_FLOW of ReadBias is
   component nBitRegister_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component my_nadder_13
      port (
         a : IN std_logic_vector (12 DOWNTO 0) ;
         b : IN std_logic_vector (12 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (12 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal upAddress_12, upAddress_11, upAddress_10, upAddress_9, upAddress_8, 
      upAddress_7, upAddress_6, upAddress_5, upAddress_4, upAddress_3, 
      upAddress_2, upAddress_1, upAddress_0, BiasEnable, Zeros_8, nx370, 
      nx372, nx374, nx376, nx378: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   B0 : nBitRegister_16 port map ( D(15)=>BIAS(15), D(14)=>BIAS(14), D(13)=>
      BIAS(13), D(12)=>BIAS(12), D(11)=>BIAS(11), D(10)=>BIAS(10), D(9)=>
      BIAS(9), D(8)=>BIAS(8), D(7)=>BIAS(7), D(6)=>BIAS(6), D(5)=>BIAS(5), 
      D(4)=>BIAS(4), D(3)=>BIAS(3), D(2)=>BIAS(2), D(1)=>BIAS(1), D(0)=>
      BIAS(0), CLK=>nx372, RST=>RST, EN=>BiasEnable, Q(15)=>outBias0(15), 
      Q(14)=>outBias0(14), Q(13)=>outBias0(13), Q(12)=>outBias0(12), Q(11)=>
      outBias0(11), Q(10)=>outBias0(10), Q(9)=>outBias0(9), Q(8)=>
      outBias0(8), Q(7)=>outBias0(7), Q(6)=>outBias0(6), Q(5)=>outBias0(5), 
      Q(4)=>outBias0(4), Q(3)=>outBias0(3), Q(2)=>outBias0(2), Q(1)=>
      outBias0(1), Q(0)=>outBias0(0));
   B1 : nBitRegister_16 port map ( D(15)=>BIAS(31), D(14)=>BIAS(30), D(13)=>
      BIAS(29), D(12)=>BIAS(28), D(11)=>BIAS(27), D(10)=>BIAS(26), D(9)=>
      BIAS(25), D(8)=>BIAS(24), D(7)=>BIAS(23), D(6)=>BIAS(22), D(5)=>
      BIAS(21), D(4)=>BIAS(20), D(3)=>BIAS(19), D(2)=>BIAS(18), D(1)=>
      BIAS(17), D(0)=>BIAS(16), CLK=>nx372, RST=>RST, EN=>BiasEnable, Q(15)
      =>outBias1(15), Q(14)=>outBias1(14), Q(13)=>outBias1(13), Q(12)=>
      outBias1(12), Q(11)=>outBias1(11), Q(10)=>outBias1(10), Q(9)=>
      outBias1(9), Q(8)=>outBias1(8), Q(7)=>outBias1(7), Q(6)=>outBias1(6), 
      Q(5)=>outBias1(5), Q(4)=>outBias1(4), Q(3)=>outBias1(3), Q(2)=>
      outBias1(2), Q(1)=>outBias1(1), Q(0)=>outBias1(0));
   B2 : nBitRegister_16 port map ( D(15)=>BIAS(47), D(14)=>BIAS(46), D(13)=>
      BIAS(45), D(12)=>BIAS(44), D(11)=>BIAS(43), D(10)=>BIAS(42), D(9)=>
      BIAS(41), D(8)=>BIAS(40), D(7)=>BIAS(39), D(6)=>BIAS(38), D(5)=>
      BIAS(37), D(4)=>BIAS(36), D(3)=>BIAS(35), D(2)=>BIAS(34), D(1)=>
      BIAS(33), D(0)=>BIAS(32), CLK=>nx374, RST=>RST, EN=>BiasEnable, Q(15)
      =>outBias2(15), Q(14)=>outBias2(14), Q(13)=>outBias2(13), Q(12)=>
      outBias2(12), Q(11)=>outBias2(11), Q(10)=>outBias2(10), Q(9)=>
      outBias2(9), Q(8)=>outBias2(8), Q(7)=>outBias2(7), Q(6)=>outBias2(6), 
      Q(5)=>outBias2(5), Q(4)=>outBias2(4), Q(3)=>outBias2(3), Q(2)=>
      outBias2(2), Q(1)=>outBias2(1), Q(0)=>outBias2(0));
   B3 : nBitRegister_16 port map ( D(15)=>BIAS(63), D(14)=>BIAS(62), D(13)=>
      BIAS(61), D(12)=>BIAS(60), D(11)=>BIAS(59), D(10)=>BIAS(58), D(9)=>
      BIAS(57), D(8)=>BIAS(56), D(7)=>BIAS(55), D(6)=>BIAS(54), D(5)=>
      BIAS(53), D(4)=>BIAS(52), D(3)=>BIAS(51), D(2)=>BIAS(50), D(1)=>
      BIAS(49), D(0)=>BIAS(48), CLK=>nx374, RST=>RST, EN=>BiasEnable, Q(15)
      =>outBias3(15), Q(14)=>outBias3(14), Q(13)=>outBias3(13), Q(12)=>
      outBias3(12), Q(11)=>outBias3(11), Q(10)=>outBias3(10), Q(9)=>
      outBias3(9), Q(8)=>outBias3(8), Q(7)=>outBias3(7), Q(6)=>outBias3(6), 
      Q(5)=>outBias3(5), Q(4)=>outBias3(4), Q(3)=>outBias3(3), Q(2)=>
      outBias3(2), Q(1)=>outBias3(1), Q(0)=>outBias3(0));
   B4 : nBitRegister_16 port map ( D(15)=>BIAS(79), D(14)=>BIAS(78), D(13)=>
      BIAS(77), D(12)=>BIAS(76), D(11)=>BIAS(75), D(10)=>BIAS(74), D(9)=>
      BIAS(73), D(8)=>BIAS(72), D(7)=>BIAS(71), D(6)=>BIAS(70), D(5)=>
      BIAS(69), D(4)=>BIAS(68), D(3)=>BIAS(67), D(2)=>BIAS(66), D(1)=>
      BIAS(65), D(0)=>BIAS(64), CLK=>nx376, RST=>RST, EN=>BiasEnable, Q(15)
      =>outBias4(15), Q(14)=>outBias4(14), Q(13)=>outBias4(13), Q(12)=>
      outBias4(12), Q(11)=>outBias4(11), Q(10)=>outBias4(10), Q(9)=>
      outBias4(9), Q(8)=>outBias4(8), Q(7)=>outBias4(7), Q(6)=>outBias4(6), 
      Q(5)=>outBias4(5), Q(4)=>outBias4(4), Q(3)=>outBias4(3), Q(2)=>
      outBias4(2), Q(1)=>outBias4(1), Q(0)=>outBias4(0));
   B5 : nBitRegister_16 port map ( D(15)=>BIAS(95), D(14)=>BIAS(94), D(13)=>
      BIAS(93), D(12)=>BIAS(92), D(11)=>BIAS(91), D(10)=>BIAS(90), D(9)=>
      BIAS(89), D(8)=>BIAS(88), D(7)=>BIAS(87), D(6)=>BIAS(86), D(5)=>
      BIAS(85), D(4)=>BIAS(84), D(3)=>BIAS(83), D(2)=>BIAS(82), D(1)=>
      BIAS(81), D(0)=>BIAS(80), CLK=>nx376, RST=>RST, EN=>BiasEnable, Q(15)
      =>outBias5(15), Q(14)=>outBias5(14), Q(13)=>outBias5(13), Q(12)=>
      outBias5(12), Q(11)=>outBias5(11), Q(10)=>outBias5(10), Q(9)=>
      outBias5(9), Q(8)=>outBias5(8), Q(7)=>outBias5(7), Q(6)=>outBias5(6), 
      Q(5)=>outBias5(5), Q(4)=>outBias5(4), Q(3)=>outBias5(3), Q(2)=>
      outBias5(2), Q(1)=>outBias5(1), Q(0)=>outBias5(0));
   B6 : nBitRegister_16 port map ( D(15)=>BIAS(111), D(14)=>BIAS(110), D(13)
      =>BIAS(109), D(12)=>BIAS(108), D(11)=>BIAS(107), D(10)=>BIAS(106), 
      D(9)=>BIAS(105), D(8)=>BIAS(104), D(7)=>BIAS(103), D(6)=>BIAS(102), 
      D(5)=>BIAS(101), D(4)=>BIAS(100), D(3)=>BIAS(99), D(2)=>BIAS(98), D(1)
      =>BIAS(97), D(0)=>BIAS(96), CLK=>nx378, RST=>RST, EN=>BiasEnable, 
      Q(15)=>outBias6(15), Q(14)=>outBias6(14), Q(13)=>outBias6(13), Q(12)=>
      outBias6(12), Q(11)=>outBias6(11), Q(10)=>outBias6(10), Q(9)=>
      outBias6(9), Q(8)=>outBias6(8), Q(7)=>outBias6(7), Q(6)=>outBias6(6), 
      Q(5)=>outBias6(5), Q(4)=>outBias6(4), Q(3)=>outBias6(3), Q(2)=>
      outBias6(2), Q(1)=>outBias6(1), Q(0)=>outBias6(0));
   B7 : nBitRegister_16 port map ( D(15)=>BIAS(127), D(14)=>BIAS(126), D(13)
      =>BIAS(125), D(12)=>BIAS(124), D(11)=>BIAS(123), D(10)=>BIAS(122), 
      D(9)=>BIAS(121), D(8)=>BIAS(120), D(7)=>BIAS(119), D(6)=>BIAS(118), 
      D(5)=>BIAS(117), D(4)=>BIAS(116), D(3)=>BIAS(115), D(2)=>BIAS(114), 
      D(1)=>BIAS(113), D(0)=>BIAS(112), CLK=>nx378, RST=>RST, EN=>BiasEnable, 
      Q(15)=>outBias7(15), Q(14)=>outBias7(14), Q(13)=>outBias7(13), Q(12)=>
      outBias7(12), Q(11)=>outBias7(11), Q(10)=>outBias7(10), Q(9)=>
      outBias7(9), Q(8)=>outBias7(8), Q(7)=>outBias7(7), Q(6)=>outBias7(6), 
      Q(5)=>outBias7(5), Q(4)=>outBias7(4), Q(3)=>outBias7(3), Q(2)=>
      outBias7(2), Q(1)=>outBias7(1), Q(0)=>outBias7(0));
   tsb0 : triStateBuffer_13 port map ( D(12)=>FilterAddress(12), D(11)=>
      FilterAddress(11), D(10)=>FilterAddress(10), D(9)=>FilterAddress(9), 
      D(8)=>FilterAddress(8), D(7)=>FilterAddress(7), D(6)=>FilterAddress(6), 
      D(5)=>FilterAddress(5), D(4)=>FilterAddress(4), D(3)=>FilterAddress(3), 
      D(2)=>FilterAddress(2), D(1)=>FilterAddress(1), D(0)=>FilterAddress(0), 
      EN=>current_state(4), F(12)=>DMAAddressToFilter(12), F(11)=>
      DMAAddressToFilter(11), F(10)=>DMAAddressToFilter(10), F(9)=>
      DMAAddressToFilter(9), F(8)=>DMAAddressToFilter(8), F(7)=>
      DMAAddressToFilter(7), F(6)=>DMAAddressToFilter(6), F(5)=>
      DMAAddressToFilter(5), F(4)=>DMAAddressToFilter(4), F(3)=>
      DMAAddressToFilter(3), F(2)=>DMAAddressToFilter(2), F(1)=>
      DMAAddressToFilter(1), F(0)=>DMAAddressToFilter(0));
   adder0 : my_nadder_13 port map ( a(12)=>FilterAddress(12), a(11)=>
      FilterAddress(11), a(10)=>FilterAddress(10), a(9)=>FilterAddress(9), 
      a(8)=>FilterAddress(8), a(7)=>FilterAddress(7), a(6)=>FilterAddress(6), 
      a(5)=>FilterAddress(5), a(4)=>FilterAddress(4), a(3)=>FilterAddress(3), 
      a(2)=>FilterAddress(2), a(1)=>FilterAddress(1), a(0)=>FilterAddress(0), 
      b(12)=>Zeros_8, b(11)=>Zeros_8, b(10)=>Zeros_8, b(9)=>Zeros_8, b(8)=>
      Zeros_8, b(7)=>Zeros_8, b(6)=>Zeros_8, b(5)=>Zeros_8, b(4)=>Zeros_8, 
      b(3)=>LayerInfo(3), b(2)=>LayerInfo(2), b(1)=>LayerInfo(1), b(0)=>
      LayerInfo(0), cin=>Zeros_8, s(12)=>upAddress_12, s(11)=>upAddress_11, 
      s(10)=>upAddress_10, s(9)=>upAddress_9, s(8)=>upAddress_8, s(7)=>
      upAddress_7, s(6)=>upAddress_6, s(5)=>upAddress_5, s(4)=>upAddress_4, 
      s(3)=>upAddress_3, s(2)=>upAddress_2, s(1)=>upAddress_1, s(0)=>
      upAddress_0, cout=>DANGLING(0));
   TriStateAdd : triStateBuffer_13 port map ( D(12)=>upAddress_12, D(11)=>
      upAddress_11, D(10)=>upAddress_10, D(9)=>upAddress_9, D(8)=>
      upAddress_8, D(7)=>upAddress_7, D(6)=>upAddress_6, D(5)=>upAddress_5, 
      D(4)=>upAddress_4, D(3)=>upAddress_3, D(2)=>upAddress_2, D(1)=>
      upAddress_1, D(0)=>upAddress_0, EN=>current_state(4), F(12)=>
      UpdatedAddress(12), F(11)=>UpdatedAddress(11), F(10)=>
      UpdatedAddress(10), F(9)=>UpdatedAddress(9), F(8)=>UpdatedAddress(8), 
      F(7)=>UpdatedAddress(7), F(6)=>UpdatedAddress(6), F(5)=>
      UpdatedAddress(5), F(4)=>UpdatedAddress(4), F(3)=>UpdatedAddress(3), 
      F(2)=>UpdatedAddress(2), F(1)=>UpdatedAddress(1), F(0)=>
      UpdatedAddress(0));
   TriStateAddchanger : triStateBuffer_13 port map ( D(12)=>upAddress_12, 
      D(11)=>upAddress_11, D(10)=>upAddress_10, D(9)=>upAddress_9, D(8)=>
      upAddress_8, D(7)=>upAddress_7, D(6)=>upAddress_6, D(5)=>upAddress_5, 
      D(4)=>upAddress_4, D(3)=>upAddress_3, D(2)=>upAddress_2, D(1)=>
      upAddress_1, D(0)=>upAddress_0, EN=>current_state(4), F(12)=>
      changerAdd(12), F(11)=>changerAdd(11), F(10)=>changerAdd(10), F(9)=>
      changerAdd(9), F(8)=>changerAdd(8), F(7)=>changerAdd(7), F(6)=>
      changerAdd(6), F(5)=>changerAdd(5), F(4)=>changerAdd(4), F(3)=>
      changerAdd(3), F(2)=>changerAdd(2), F(1)=>changerAdd(1), F(0)=>
      changerAdd(0));
   ix355 : fake_gnd port map ( Y=>Zeros_8);
   ix1 : and02 port map ( Y=>BiasEnable, A0=>ACKF, A1=>current_state(4));
   ix369 : inv01 port map ( Y=>nx370, A=>CLK);
   ix371 : inv02 port map ( Y=>nx372, A=>nx370);
   ix373 : inv02 port map ( Y=>nx374, A=>nx370);
   ix375 : inv02 port map ( Y=>nx376, A=>nx370);
   ix377 : inv02 port map ( Y=>nx378, A=>nx370);
end DATA_FLOW ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity my_nadder_4 is
   port (
      a : IN std_logic_vector (3 DOWNTO 0) ;
      b : IN std_logic_vector (3 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (3 DOWNTO 0) ;
      cout : OUT std_logic) ;
end my_nadder_4 ;

architecture a_my_nadder of my_nadder_4 is
   component my_adder
      port (
         a : IN std_logic ;
         b : IN std_logic ;
         cin : IN std_logic ;
         s : OUT std_logic ;
         cout : OUT std_logic) ;
   end component ;
   signal temp_2, temp_1, temp_0: std_logic ;

begin
   f0 : my_adder port map ( a=>a(0), b=>b(0), cin=>cin, s=>s(0), cout=>
      temp_0);
   loop1_1_fx : my_adder port map ( a=>a(1), b=>b(1), cin=>temp_0, s=>s(1), 
      cout=>temp_1);
   loop1_2_fx : my_adder port map ( a=>a(2), b=>b(2), cin=>temp_1, s=>s(2), 
      cout=>temp_2);
   loop1_3_fx : my_adder port map ( a=>a(3), b=>b(3), cin=>temp_2, s=>s(3), 
      cout=>cout);
end a_my_nadder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity nBitRegister_400 is
   port (
      D : IN std_logic_vector (399 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      EN : IN std_logic ;
      Q : OUT std_logic_vector (399 DOWNTO 0)) ;
end nBitRegister_400 ;

architecture Data_flow of nBitRegister_400 is
   signal Q_399_EXMPLR, Q_398_EXMPLR, Q_397_EXMPLR, Q_396_EXMPLR, 
      Q_395_EXMPLR, Q_394_EXMPLR, Q_393_EXMPLR, Q_392_EXMPLR, Q_391_EXMPLR, 
      Q_390_EXMPLR, Q_389_EXMPLR, Q_388_EXMPLR, Q_387_EXMPLR, Q_386_EXMPLR, 
      Q_385_EXMPLR, Q_384_EXMPLR, Q_383_EXMPLR, Q_382_EXMPLR, Q_381_EXMPLR, 
      Q_380_EXMPLR, Q_379_EXMPLR, Q_378_EXMPLR, Q_377_EXMPLR, Q_376_EXMPLR, 
      Q_375_EXMPLR, Q_374_EXMPLR, Q_373_EXMPLR, Q_372_EXMPLR, Q_371_EXMPLR, 
      Q_370_EXMPLR, Q_369_EXMPLR, Q_368_EXMPLR, Q_367_EXMPLR, Q_366_EXMPLR, 
      Q_365_EXMPLR, Q_364_EXMPLR, Q_363_EXMPLR, Q_362_EXMPLR, Q_361_EXMPLR, 
      Q_360_EXMPLR, Q_359_EXMPLR, Q_358_EXMPLR, Q_357_EXMPLR, Q_356_EXMPLR, 
      Q_355_EXMPLR, Q_354_EXMPLR, Q_353_EXMPLR, Q_352_EXMPLR, Q_351_EXMPLR, 
      Q_350_EXMPLR, Q_349_EXMPLR, Q_348_EXMPLR, Q_347_EXMPLR, Q_346_EXMPLR, 
      Q_345_EXMPLR, Q_344_EXMPLR, Q_343_EXMPLR, Q_342_EXMPLR, Q_341_EXMPLR, 
      Q_340_EXMPLR, Q_339_EXMPLR, Q_338_EXMPLR, Q_337_EXMPLR, Q_336_EXMPLR, 
      Q_335_EXMPLR, Q_334_EXMPLR, Q_333_EXMPLR, Q_332_EXMPLR, Q_331_EXMPLR, 
      Q_330_EXMPLR, Q_329_EXMPLR, Q_328_EXMPLR, Q_327_EXMPLR, Q_326_EXMPLR, 
      Q_325_EXMPLR, Q_324_EXMPLR, Q_323_EXMPLR, Q_322_EXMPLR, Q_321_EXMPLR, 
      Q_320_EXMPLR, Q_319_EXMPLR, Q_318_EXMPLR, Q_317_EXMPLR, Q_316_EXMPLR, 
      Q_315_EXMPLR, Q_314_EXMPLR, Q_313_EXMPLR, Q_312_EXMPLR, Q_311_EXMPLR, 
      Q_310_EXMPLR, Q_309_EXMPLR, Q_308_EXMPLR, Q_307_EXMPLR, Q_306_EXMPLR, 
      Q_305_EXMPLR, Q_304_EXMPLR, Q_303_EXMPLR, Q_302_EXMPLR, Q_301_EXMPLR, 
      Q_300_EXMPLR, Q_299_EXMPLR, Q_298_EXMPLR, Q_297_EXMPLR, Q_296_EXMPLR, 
      Q_295_EXMPLR, Q_294_EXMPLR, Q_293_EXMPLR, Q_292_EXMPLR, Q_291_EXMPLR, 
      Q_290_EXMPLR, Q_289_EXMPLR, Q_288_EXMPLR, Q_287_EXMPLR, Q_286_EXMPLR, 
      Q_285_EXMPLR, Q_284_EXMPLR, Q_283_EXMPLR, Q_282_EXMPLR, Q_281_EXMPLR, 
      Q_280_EXMPLR, Q_279_EXMPLR, Q_278_EXMPLR, Q_277_EXMPLR, Q_276_EXMPLR, 
      Q_275_EXMPLR, Q_274_EXMPLR, Q_273_EXMPLR, Q_272_EXMPLR, Q_271_EXMPLR, 
      Q_270_EXMPLR, Q_269_EXMPLR, Q_268_EXMPLR, Q_267_EXMPLR, Q_266_EXMPLR, 
      Q_265_EXMPLR, Q_264_EXMPLR, Q_263_EXMPLR, Q_262_EXMPLR, Q_261_EXMPLR, 
      Q_260_EXMPLR, Q_259_EXMPLR, Q_258_EXMPLR, Q_257_EXMPLR, Q_256_EXMPLR, 
      Q_255_EXMPLR, Q_254_EXMPLR, Q_253_EXMPLR, Q_252_EXMPLR, Q_251_EXMPLR, 
      Q_250_EXMPLR, Q_249_EXMPLR, Q_248_EXMPLR, Q_247_EXMPLR, Q_246_EXMPLR, 
      Q_245_EXMPLR, Q_244_EXMPLR, Q_243_EXMPLR, Q_242_EXMPLR, Q_241_EXMPLR, 
      Q_240_EXMPLR, Q_239_EXMPLR, Q_238_EXMPLR, Q_237_EXMPLR, Q_236_EXMPLR, 
      Q_235_EXMPLR, Q_234_EXMPLR, Q_233_EXMPLR, Q_232_EXMPLR, Q_231_EXMPLR, 
      Q_230_EXMPLR, Q_229_EXMPLR, Q_228_EXMPLR, Q_227_EXMPLR, Q_226_EXMPLR, 
      Q_225_EXMPLR, Q_224_EXMPLR, Q_223_EXMPLR, Q_222_EXMPLR, Q_221_EXMPLR, 
      Q_220_EXMPLR, Q_219_EXMPLR, Q_218_EXMPLR, Q_217_EXMPLR, Q_216_EXMPLR, 
      Q_215_EXMPLR, Q_214_EXMPLR, Q_213_EXMPLR, Q_212_EXMPLR, Q_211_EXMPLR, 
      Q_210_EXMPLR, Q_209_EXMPLR, Q_208_EXMPLR, Q_207_EXMPLR, Q_206_EXMPLR, 
      Q_205_EXMPLR, Q_204_EXMPLR, Q_203_EXMPLR, Q_202_EXMPLR, Q_201_EXMPLR, 
      Q_200_EXMPLR, Q_199_EXMPLR, Q_198_EXMPLR, Q_197_EXMPLR, Q_196_EXMPLR, 
      Q_195_EXMPLR, Q_194_EXMPLR, Q_193_EXMPLR, Q_192_EXMPLR, Q_191_EXMPLR, 
      Q_190_EXMPLR, Q_189_EXMPLR, Q_188_EXMPLR, Q_187_EXMPLR, Q_186_EXMPLR, 
      Q_185_EXMPLR, Q_184_EXMPLR, Q_183_EXMPLR, Q_182_EXMPLR, Q_181_EXMPLR, 
      Q_180_EXMPLR, Q_179_EXMPLR, Q_178_EXMPLR, Q_177_EXMPLR, Q_176_EXMPLR, 
      Q_175_EXMPLR, Q_174_EXMPLR, Q_173_EXMPLR, Q_172_EXMPLR, Q_171_EXMPLR, 
      Q_170_EXMPLR, Q_169_EXMPLR, Q_168_EXMPLR, Q_167_EXMPLR, Q_166_EXMPLR, 
      Q_165_EXMPLR, Q_164_EXMPLR, Q_163_EXMPLR, Q_162_EXMPLR, Q_161_EXMPLR, 
      Q_160_EXMPLR, Q_159_EXMPLR, Q_158_EXMPLR, Q_157_EXMPLR, Q_156_EXMPLR, 
      Q_155_EXMPLR, Q_154_EXMPLR, Q_153_EXMPLR, Q_152_EXMPLR, Q_151_EXMPLR, 
      Q_150_EXMPLR, Q_149_EXMPLR, Q_148_EXMPLR, Q_147_EXMPLR, Q_146_EXMPLR, 
      Q_145_EXMPLR, Q_144_EXMPLR, Q_143_EXMPLR, Q_142_EXMPLR, Q_141_EXMPLR, 
      Q_140_EXMPLR, Q_139_EXMPLR, Q_138_EXMPLR, Q_137_EXMPLR, Q_136_EXMPLR, 
      Q_135_EXMPLR, Q_134_EXMPLR, Q_133_EXMPLR, Q_132_EXMPLR, Q_131_EXMPLR, 
      Q_130_EXMPLR, Q_129_EXMPLR, Q_128_EXMPLR, Q_127_EXMPLR, Q_126_EXMPLR, 
      Q_125_EXMPLR, Q_124_EXMPLR, Q_123_EXMPLR, Q_122_EXMPLR, Q_121_EXMPLR, 
      Q_120_EXMPLR, Q_119_EXMPLR, Q_118_EXMPLR, Q_117_EXMPLR, Q_116_EXMPLR, 
      Q_115_EXMPLR, Q_114_EXMPLR, Q_113_EXMPLR, Q_112_EXMPLR, Q_111_EXMPLR, 
      Q_110_EXMPLR, Q_109_EXMPLR, Q_108_EXMPLR, Q_107_EXMPLR, Q_106_EXMPLR, 
      Q_105_EXMPLR, Q_104_EXMPLR, Q_103_EXMPLR, Q_102_EXMPLR, Q_101_EXMPLR, 
      Q_100_EXMPLR, Q_99_EXMPLR, Q_98_EXMPLR, Q_97_EXMPLR, Q_96_EXMPLR, 
      Q_95_EXMPLR, Q_94_EXMPLR, Q_93_EXMPLR, Q_92_EXMPLR, Q_91_EXMPLR, 
      Q_90_EXMPLR, Q_89_EXMPLR, Q_88_EXMPLR, Q_87_EXMPLR, Q_86_EXMPLR, 
      Q_85_EXMPLR, Q_84_EXMPLR, Q_83_EXMPLR, Q_82_EXMPLR, Q_81_EXMPLR, 
      Q_80_EXMPLR, Q_79_EXMPLR, Q_78_EXMPLR, Q_77_EXMPLR, Q_76_EXMPLR, 
      Q_75_EXMPLR, Q_74_EXMPLR, Q_73_EXMPLR, Q_72_EXMPLR, Q_71_EXMPLR, 
      Q_70_EXMPLR, Q_69_EXMPLR, Q_68_EXMPLR, Q_67_EXMPLR, Q_66_EXMPLR, 
      Q_65_EXMPLR, Q_64_EXMPLR, Q_63_EXMPLR, Q_62_EXMPLR, Q_61_EXMPLR, 
      Q_60_EXMPLR, Q_59_EXMPLR, Q_58_EXMPLR, Q_57_EXMPLR, Q_56_EXMPLR, 
      Q_55_EXMPLR, Q_54_EXMPLR, Q_53_EXMPLR, Q_52_EXMPLR, Q_51_EXMPLR, 
      Q_50_EXMPLR, Q_49_EXMPLR, Q_48_EXMPLR, Q_47_EXMPLR, Q_46_EXMPLR, 
      Q_45_EXMPLR, Q_44_EXMPLR, Q_43_EXMPLR, Q_42_EXMPLR, Q_41_EXMPLR, 
      Q_40_EXMPLR, Q_39_EXMPLR, Q_38_EXMPLR, Q_37_EXMPLR, Q_36_EXMPLR, 
      Q_35_EXMPLR, Q_34_EXMPLR, Q_33_EXMPLR, Q_32_EXMPLR, Q_31_EXMPLR, 
      Q_30_EXMPLR, Q_29_EXMPLR, Q_28_EXMPLR, Q_27_EXMPLR, Q_26_EXMPLR, 
      Q_25_EXMPLR, Q_24_EXMPLR, Q_23_EXMPLR, Q_22_EXMPLR, Q_21_EXMPLR, 
      Q_20_EXMPLR, Q_19_EXMPLR, Q_18_EXMPLR, Q_17_EXMPLR, Q_16_EXMPLR, 
      Q_15_EXMPLR, Q_14_EXMPLR, Q_13_EXMPLR, Q_12_EXMPLR, Q_11_EXMPLR, 
      Q_10_EXMPLR, Q_9_EXMPLR, Q_8_EXMPLR, Q_7_EXMPLR, Q_6_EXMPLR, 
      Q_5_EXMPLR, Q_4_EXMPLR, Q_3_EXMPLR, Q_2_EXMPLR, Q_1_EXMPLR, Q_0_EXMPLR, 
      nx4838, nx4848, nx4858, nx4868, nx4878, nx4888, nx4898, nx4908, nx4918, 
      nx4928, nx4938, nx4948, nx4958, nx4968, nx4978, nx4988, nx4998, nx5008, 
      nx5018, nx5028, nx5038, nx5048, nx5058, nx5068, nx5078, nx5088, nx5098, 
      nx5108, nx5118, nx5128, nx5138, nx5148, nx5158, nx5168, nx5178, nx5188, 
      nx5198, nx5208, nx5218, nx5228, nx5238, nx5248, nx5258, nx5268, nx5278, 
      nx5288, nx5298, nx5308, nx5318, nx5328, nx5338, nx5348, nx5358, nx5368, 
      nx5378, nx5388, nx5398, nx5408, nx5418, nx5428, nx5438, nx5448, nx5458, 
      nx5468, nx5478, nx5488, nx5498, nx5508, nx5518, nx5528, nx5538, nx5548, 
      nx5558, nx5568, nx5578, nx5588, nx5598, nx5608, nx5618, nx5628, nx5638, 
      nx5648, nx5658, nx5668, nx5678, nx5688, nx5698, nx5708, nx5718, nx5728, 
      nx5738, nx5748, nx5758, nx5768, nx5778, nx5788, nx5798, nx5808, nx5818, 
      nx5828, nx5838, nx5848, nx5858, nx5868, nx5878, nx5888, nx5898, nx5908, 
      nx5918, nx5928, nx5938, nx5948, nx5958, nx5968, nx5978, nx5988, nx5998, 
      nx6008, nx6018, nx6028, nx6038, nx6048, nx6058, nx6068, nx6078, nx6088, 
      nx6098, nx6108, nx6118, nx6128, nx6138, nx6148, nx6158, nx6168, nx6178, 
      nx6188, nx6198, nx6208, nx6218, nx6228, nx6238, nx6248, nx6258, nx6268, 
      nx6278, nx6288, nx6298, nx6308, nx6318, nx6328, nx6338, nx6348, nx6358, 
      nx6368, nx6378, nx6388, nx6398, nx6408, nx6418, nx6428, nx6438, nx6448, 
      nx6458, nx6468, nx6478, nx6488, nx6498, nx6508, nx6518, nx6528, nx6538, 
      nx6548, nx6558, nx6568, nx6578, nx6588, nx6598, nx6608, nx6618, nx6628, 
      nx6638, nx6648, nx6658, nx6668, nx6678, nx6688, nx6698, nx6708, nx6718, 
      nx6728, nx6738, nx6748, nx6758, nx6768, nx6778, nx6788, nx6798, nx6808, 
      nx6818, nx6828, nx6838, nx6848, nx6858, nx6868, nx6878, nx6888, nx6898, 
      nx6908, nx6918, nx6928, nx6938, nx6948, nx6958, nx6968, nx6978, nx6988, 
      nx6998, nx7008, nx7018, nx7028, nx7038, nx7048, nx7058, nx7068, nx7078, 
      nx7088, nx7098, nx7108, nx7118, nx7128, nx7138, nx7148, nx7158, nx7168, 
      nx7178, nx7188, nx7198, nx7208, nx7218, nx7228, nx7238, nx7248, nx7258, 
      nx7268, nx7278, nx7288, nx7298, nx7308, nx7318, nx7328, nx7338, nx7348, 
      nx7358, nx7368, nx7378, nx7388, nx7398, nx7408, nx7418, nx7428, nx7438, 
      nx7448, nx7458, nx7468, nx7478, nx7488, nx7498, nx7508, nx7518, nx7528, 
      nx7538, nx7548, nx7558, nx7568, nx7578, nx7588, nx7598, nx7608, nx7618, 
      nx7628, nx7638, nx7648, nx7658, nx7668, nx7678, nx7688, nx7698, nx7708, 
      nx7718, nx7728, nx7738, nx7748, nx7758, nx7768, nx7778, nx7788, nx7798, 
      nx7808, nx7818, nx7828, nx7838, nx7848, nx7858, nx7868, nx7878, nx7888, 
      nx7898, nx7908, nx7918, nx7928, nx7938, nx7948, nx7958, nx7968, nx7978, 
      nx7988, nx7998, nx8008, nx8018, nx8028, nx8038, nx8048, nx8058, nx8068, 
      nx8078, nx8088, nx8098, nx8108, nx8118, nx8128, nx8138, nx8148, nx8158, 
      nx8168, nx8178, nx8188, nx8198, nx8208, nx8218, nx8228, nx8238, nx8248, 
      nx8258, nx8268, nx8278, nx8288, nx8298, nx8308, nx8318, nx8328, nx8338, 
      nx8348, nx8358, nx8368, nx8378, nx8388, nx8398, nx8408, nx8418, nx8428, 
      nx8438, nx8448, nx8458, nx8468, nx8478, nx8488, nx8498, nx8508, nx8518, 
      nx8528, nx8538, nx8548, nx8558, nx8568, nx8578, nx8588, nx8598, nx8608, 
      nx8618, nx8628, nx8638, nx8648, nx8658, nx8668, nx8678, nx8688, nx8698, 
      nx8708, nx8718, nx8728, nx8738, nx8748, nx8758, nx8768, nx8778, nx8788, 
      nx8798, nx8808, nx8818, nx8828, nx10045, nx10047, nx10049, nx10051, 
      nx10053, nx10055, nx10057, nx10059, nx10061, nx10063, nx10065, nx10067, 
      nx10069, nx10071, nx10073, nx10075, nx10077, nx10079, nx10081, nx10083, 
      nx10085, nx10087, nx10089, nx10091, nx10093, nx10095, nx10097, nx10099, 
      nx10101, nx10103, nx10105, nx10107, nx10109, nx10111, nx10113, nx10115, 
      nx10117, nx10119, nx10121, nx10123, nx10125, nx10127, nx10129, nx10131, 
      nx10133, nx10135, nx10137, nx10139, nx10141, nx10143, nx10145, nx10147, 
      nx10149, nx10151, nx10153, nx10155, nx10157, nx10159, nx10167, nx10169, 
      nx10171, nx10173, nx10175, nx10177, nx10179, nx10181, nx10183, nx10185, 
      nx10187, nx10189, nx10191, nx10193, nx10195, nx10197, nx10199, nx10201, 
      nx10203, nx10205, nx10207, nx10209, nx10211, nx10213, nx10215, nx10217, 
      nx10219, nx10221, nx10223, nx10225, nx10227, nx10229, nx10231, nx10233, 
      nx10235, nx10237, nx10239, nx10241, nx10243, nx10245, nx10247, nx10249, 
      nx10251, nx10253, nx10255, nx10257, nx10259, nx10261, nx10263, nx10265, 
      nx10267, nx10269, nx10271, nx10273, nx10275, nx10277, nx10279, nx10281, 
      nx10283, nx10285, nx10287, nx10289, nx10291, nx10293, nx10295, nx10297, 
      nx10299, nx10301, nx10303, nx10305, nx10307, nx10309, nx10311, nx10313, 
      nx10315, nx10317, nx10319, nx10321, nx10327, nx10329: std_logic ;

begin
   Q(399) <= Q_399_EXMPLR ;
   Q(398) <= Q_398_EXMPLR ;
   Q(397) <= Q_397_EXMPLR ;
   Q(396) <= Q_396_EXMPLR ;
   Q(395) <= Q_395_EXMPLR ;
   Q(394) <= Q_394_EXMPLR ;
   Q(393) <= Q_393_EXMPLR ;
   Q(392) <= Q_392_EXMPLR ;
   Q(391) <= Q_391_EXMPLR ;
   Q(390) <= Q_390_EXMPLR ;
   Q(389) <= Q_389_EXMPLR ;
   Q(388) <= Q_388_EXMPLR ;
   Q(387) <= Q_387_EXMPLR ;
   Q(386) <= Q_386_EXMPLR ;
   Q(385) <= Q_385_EXMPLR ;
   Q(384) <= Q_384_EXMPLR ;
   Q(383) <= Q_383_EXMPLR ;
   Q(382) <= Q_382_EXMPLR ;
   Q(381) <= Q_381_EXMPLR ;
   Q(380) <= Q_380_EXMPLR ;
   Q(379) <= Q_379_EXMPLR ;
   Q(378) <= Q_378_EXMPLR ;
   Q(377) <= Q_377_EXMPLR ;
   Q(376) <= Q_376_EXMPLR ;
   Q(375) <= Q_375_EXMPLR ;
   Q(374) <= Q_374_EXMPLR ;
   Q(373) <= Q_373_EXMPLR ;
   Q(372) <= Q_372_EXMPLR ;
   Q(371) <= Q_371_EXMPLR ;
   Q(370) <= Q_370_EXMPLR ;
   Q(369) <= Q_369_EXMPLR ;
   Q(368) <= Q_368_EXMPLR ;
   Q(367) <= Q_367_EXMPLR ;
   Q(366) <= Q_366_EXMPLR ;
   Q(365) <= Q_365_EXMPLR ;
   Q(364) <= Q_364_EXMPLR ;
   Q(363) <= Q_363_EXMPLR ;
   Q(362) <= Q_362_EXMPLR ;
   Q(361) <= Q_361_EXMPLR ;
   Q(360) <= Q_360_EXMPLR ;
   Q(359) <= Q_359_EXMPLR ;
   Q(358) <= Q_358_EXMPLR ;
   Q(357) <= Q_357_EXMPLR ;
   Q(356) <= Q_356_EXMPLR ;
   Q(355) <= Q_355_EXMPLR ;
   Q(354) <= Q_354_EXMPLR ;
   Q(353) <= Q_353_EXMPLR ;
   Q(352) <= Q_352_EXMPLR ;
   Q(351) <= Q_351_EXMPLR ;
   Q(350) <= Q_350_EXMPLR ;
   Q(349) <= Q_349_EXMPLR ;
   Q(348) <= Q_348_EXMPLR ;
   Q(347) <= Q_347_EXMPLR ;
   Q(346) <= Q_346_EXMPLR ;
   Q(345) <= Q_345_EXMPLR ;
   Q(344) <= Q_344_EXMPLR ;
   Q(343) <= Q_343_EXMPLR ;
   Q(342) <= Q_342_EXMPLR ;
   Q(341) <= Q_341_EXMPLR ;
   Q(340) <= Q_340_EXMPLR ;
   Q(339) <= Q_339_EXMPLR ;
   Q(338) <= Q_338_EXMPLR ;
   Q(337) <= Q_337_EXMPLR ;
   Q(336) <= Q_336_EXMPLR ;
   Q(335) <= Q_335_EXMPLR ;
   Q(334) <= Q_334_EXMPLR ;
   Q(333) <= Q_333_EXMPLR ;
   Q(332) <= Q_332_EXMPLR ;
   Q(331) <= Q_331_EXMPLR ;
   Q(330) <= Q_330_EXMPLR ;
   Q(329) <= Q_329_EXMPLR ;
   Q(328) <= Q_328_EXMPLR ;
   Q(327) <= Q_327_EXMPLR ;
   Q(326) <= Q_326_EXMPLR ;
   Q(325) <= Q_325_EXMPLR ;
   Q(324) <= Q_324_EXMPLR ;
   Q(323) <= Q_323_EXMPLR ;
   Q(322) <= Q_322_EXMPLR ;
   Q(321) <= Q_321_EXMPLR ;
   Q(320) <= Q_320_EXMPLR ;
   Q(319) <= Q_319_EXMPLR ;
   Q(318) <= Q_318_EXMPLR ;
   Q(317) <= Q_317_EXMPLR ;
   Q(316) <= Q_316_EXMPLR ;
   Q(315) <= Q_315_EXMPLR ;
   Q(314) <= Q_314_EXMPLR ;
   Q(313) <= Q_313_EXMPLR ;
   Q(312) <= Q_312_EXMPLR ;
   Q(311) <= Q_311_EXMPLR ;
   Q(310) <= Q_310_EXMPLR ;
   Q(309) <= Q_309_EXMPLR ;
   Q(308) <= Q_308_EXMPLR ;
   Q(307) <= Q_307_EXMPLR ;
   Q(306) <= Q_306_EXMPLR ;
   Q(305) <= Q_305_EXMPLR ;
   Q(304) <= Q_304_EXMPLR ;
   Q(303) <= Q_303_EXMPLR ;
   Q(302) <= Q_302_EXMPLR ;
   Q(301) <= Q_301_EXMPLR ;
   Q(300) <= Q_300_EXMPLR ;
   Q(299) <= Q_299_EXMPLR ;
   Q(298) <= Q_298_EXMPLR ;
   Q(297) <= Q_297_EXMPLR ;
   Q(296) <= Q_296_EXMPLR ;
   Q(295) <= Q_295_EXMPLR ;
   Q(294) <= Q_294_EXMPLR ;
   Q(293) <= Q_293_EXMPLR ;
   Q(292) <= Q_292_EXMPLR ;
   Q(291) <= Q_291_EXMPLR ;
   Q(290) <= Q_290_EXMPLR ;
   Q(289) <= Q_289_EXMPLR ;
   Q(288) <= Q_288_EXMPLR ;
   Q(287) <= Q_287_EXMPLR ;
   Q(286) <= Q_286_EXMPLR ;
   Q(285) <= Q_285_EXMPLR ;
   Q(284) <= Q_284_EXMPLR ;
   Q(283) <= Q_283_EXMPLR ;
   Q(282) <= Q_282_EXMPLR ;
   Q(281) <= Q_281_EXMPLR ;
   Q(280) <= Q_280_EXMPLR ;
   Q(279) <= Q_279_EXMPLR ;
   Q(278) <= Q_278_EXMPLR ;
   Q(277) <= Q_277_EXMPLR ;
   Q(276) <= Q_276_EXMPLR ;
   Q(275) <= Q_275_EXMPLR ;
   Q(274) <= Q_274_EXMPLR ;
   Q(273) <= Q_273_EXMPLR ;
   Q(272) <= Q_272_EXMPLR ;
   Q(271) <= Q_271_EXMPLR ;
   Q(270) <= Q_270_EXMPLR ;
   Q(269) <= Q_269_EXMPLR ;
   Q(268) <= Q_268_EXMPLR ;
   Q(267) <= Q_267_EXMPLR ;
   Q(266) <= Q_266_EXMPLR ;
   Q(265) <= Q_265_EXMPLR ;
   Q(264) <= Q_264_EXMPLR ;
   Q(263) <= Q_263_EXMPLR ;
   Q(262) <= Q_262_EXMPLR ;
   Q(261) <= Q_261_EXMPLR ;
   Q(260) <= Q_260_EXMPLR ;
   Q(259) <= Q_259_EXMPLR ;
   Q(258) <= Q_258_EXMPLR ;
   Q(257) <= Q_257_EXMPLR ;
   Q(256) <= Q_256_EXMPLR ;
   Q(255) <= Q_255_EXMPLR ;
   Q(254) <= Q_254_EXMPLR ;
   Q(253) <= Q_253_EXMPLR ;
   Q(252) <= Q_252_EXMPLR ;
   Q(251) <= Q_251_EXMPLR ;
   Q(250) <= Q_250_EXMPLR ;
   Q(249) <= Q_249_EXMPLR ;
   Q(248) <= Q_248_EXMPLR ;
   Q(247) <= Q_247_EXMPLR ;
   Q(246) <= Q_246_EXMPLR ;
   Q(245) <= Q_245_EXMPLR ;
   Q(244) <= Q_244_EXMPLR ;
   Q(243) <= Q_243_EXMPLR ;
   Q(242) <= Q_242_EXMPLR ;
   Q(241) <= Q_241_EXMPLR ;
   Q(240) <= Q_240_EXMPLR ;
   Q(239) <= Q_239_EXMPLR ;
   Q(238) <= Q_238_EXMPLR ;
   Q(237) <= Q_237_EXMPLR ;
   Q(236) <= Q_236_EXMPLR ;
   Q(235) <= Q_235_EXMPLR ;
   Q(234) <= Q_234_EXMPLR ;
   Q(233) <= Q_233_EXMPLR ;
   Q(232) <= Q_232_EXMPLR ;
   Q(231) <= Q_231_EXMPLR ;
   Q(230) <= Q_230_EXMPLR ;
   Q(229) <= Q_229_EXMPLR ;
   Q(228) <= Q_228_EXMPLR ;
   Q(227) <= Q_227_EXMPLR ;
   Q(226) <= Q_226_EXMPLR ;
   Q(225) <= Q_225_EXMPLR ;
   Q(224) <= Q_224_EXMPLR ;
   Q(223) <= Q_223_EXMPLR ;
   Q(222) <= Q_222_EXMPLR ;
   Q(221) <= Q_221_EXMPLR ;
   Q(220) <= Q_220_EXMPLR ;
   Q(219) <= Q_219_EXMPLR ;
   Q(218) <= Q_218_EXMPLR ;
   Q(217) <= Q_217_EXMPLR ;
   Q(216) <= Q_216_EXMPLR ;
   Q(215) <= Q_215_EXMPLR ;
   Q(214) <= Q_214_EXMPLR ;
   Q(213) <= Q_213_EXMPLR ;
   Q(212) <= Q_212_EXMPLR ;
   Q(211) <= Q_211_EXMPLR ;
   Q(210) <= Q_210_EXMPLR ;
   Q(209) <= Q_209_EXMPLR ;
   Q(208) <= Q_208_EXMPLR ;
   Q(207) <= Q_207_EXMPLR ;
   Q(206) <= Q_206_EXMPLR ;
   Q(205) <= Q_205_EXMPLR ;
   Q(204) <= Q_204_EXMPLR ;
   Q(203) <= Q_203_EXMPLR ;
   Q(202) <= Q_202_EXMPLR ;
   Q(201) <= Q_201_EXMPLR ;
   Q(200) <= Q_200_EXMPLR ;
   Q(199) <= Q_199_EXMPLR ;
   Q(198) <= Q_198_EXMPLR ;
   Q(197) <= Q_197_EXMPLR ;
   Q(196) <= Q_196_EXMPLR ;
   Q(195) <= Q_195_EXMPLR ;
   Q(194) <= Q_194_EXMPLR ;
   Q(193) <= Q_193_EXMPLR ;
   Q(192) <= Q_192_EXMPLR ;
   Q(191) <= Q_191_EXMPLR ;
   Q(190) <= Q_190_EXMPLR ;
   Q(189) <= Q_189_EXMPLR ;
   Q(188) <= Q_188_EXMPLR ;
   Q(187) <= Q_187_EXMPLR ;
   Q(186) <= Q_186_EXMPLR ;
   Q(185) <= Q_185_EXMPLR ;
   Q(184) <= Q_184_EXMPLR ;
   Q(183) <= Q_183_EXMPLR ;
   Q(182) <= Q_182_EXMPLR ;
   Q(181) <= Q_181_EXMPLR ;
   Q(180) <= Q_180_EXMPLR ;
   Q(179) <= Q_179_EXMPLR ;
   Q(178) <= Q_178_EXMPLR ;
   Q(177) <= Q_177_EXMPLR ;
   Q(176) <= Q_176_EXMPLR ;
   Q(175) <= Q_175_EXMPLR ;
   Q(174) <= Q_174_EXMPLR ;
   Q(173) <= Q_173_EXMPLR ;
   Q(172) <= Q_172_EXMPLR ;
   Q(171) <= Q_171_EXMPLR ;
   Q(170) <= Q_170_EXMPLR ;
   Q(169) <= Q_169_EXMPLR ;
   Q(168) <= Q_168_EXMPLR ;
   Q(167) <= Q_167_EXMPLR ;
   Q(166) <= Q_166_EXMPLR ;
   Q(165) <= Q_165_EXMPLR ;
   Q(164) <= Q_164_EXMPLR ;
   Q(163) <= Q_163_EXMPLR ;
   Q(162) <= Q_162_EXMPLR ;
   Q(161) <= Q_161_EXMPLR ;
   Q(160) <= Q_160_EXMPLR ;
   Q(159) <= Q_159_EXMPLR ;
   Q(158) <= Q_158_EXMPLR ;
   Q(157) <= Q_157_EXMPLR ;
   Q(156) <= Q_156_EXMPLR ;
   Q(155) <= Q_155_EXMPLR ;
   Q(154) <= Q_154_EXMPLR ;
   Q(153) <= Q_153_EXMPLR ;
   Q(152) <= Q_152_EXMPLR ;
   Q(151) <= Q_151_EXMPLR ;
   Q(150) <= Q_150_EXMPLR ;
   Q(149) <= Q_149_EXMPLR ;
   Q(148) <= Q_148_EXMPLR ;
   Q(147) <= Q_147_EXMPLR ;
   Q(146) <= Q_146_EXMPLR ;
   Q(145) <= Q_145_EXMPLR ;
   Q(144) <= Q_144_EXMPLR ;
   Q(143) <= Q_143_EXMPLR ;
   Q(142) <= Q_142_EXMPLR ;
   Q(141) <= Q_141_EXMPLR ;
   Q(140) <= Q_140_EXMPLR ;
   Q(139) <= Q_139_EXMPLR ;
   Q(138) <= Q_138_EXMPLR ;
   Q(137) <= Q_137_EXMPLR ;
   Q(136) <= Q_136_EXMPLR ;
   Q(135) <= Q_135_EXMPLR ;
   Q(134) <= Q_134_EXMPLR ;
   Q(133) <= Q_133_EXMPLR ;
   Q(132) <= Q_132_EXMPLR ;
   Q(131) <= Q_131_EXMPLR ;
   Q(130) <= Q_130_EXMPLR ;
   Q(129) <= Q_129_EXMPLR ;
   Q(128) <= Q_128_EXMPLR ;
   Q(127) <= Q_127_EXMPLR ;
   Q(126) <= Q_126_EXMPLR ;
   Q(125) <= Q_125_EXMPLR ;
   Q(124) <= Q_124_EXMPLR ;
   Q(123) <= Q_123_EXMPLR ;
   Q(122) <= Q_122_EXMPLR ;
   Q(121) <= Q_121_EXMPLR ;
   Q(120) <= Q_120_EXMPLR ;
   Q(119) <= Q_119_EXMPLR ;
   Q(118) <= Q_118_EXMPLR ;
   Q(117) <= Q_117_EXMPLR ;
   Q(116) <= Q_116_EXMPLR ;
   Q(115) <= Q_115_EXMPLR ;
   Q(114) <= Q_114_EXMPLR ;
   Q(113) <= Q_113_EXMPLR ;
   Q(112) <= Q_112_EXMPLR ;
   Q(111) <= Q_111_EXMPLR ;
   Q(110) <= Q_110_EXMPLR ;
   Q(109) <= Q_109_EXMPLR ;
   Q(108) <= Q_108_EXMPLR ;
   Q(107) <= Q_107_EXMPLR ;
   Q(106) <= Q_106_EXMPLR ;
   Q(105) <= Q_105_EXMPLR ;
   Q(104) <= Q_104_EXMPLR ;
   Q(103) <= Q_103_EXMPLR ;
   Q(102) <= Q_102_EXMPLR ;
   Q(101) <= Q_101_EXMPLR ;
   Q(100) <= Q_100_EXMPLR ;
   Q(99) <= Q_99_EXMPLR ;
   Q(98) <= Q_98_EXMPLR ;
   Q(97) <= Q_97_EXMPLR ;
   Q(96) <= Q_96_EXMPLR ;
   Q(95) <= Q_95_EXMPLR ;
   Q(94) <= Q_94_EXMPLR ;
   Q(93) <= Q_93_EXMPLR ;
   Q(92) <= Q_92_EXMPLR ;
   Q(91) <= Q_91_EXMPLR ;
   Q(90) <= Q_90_EXMPLR ;
   Q(89) <= Q_89_EXMPLR ;
   Q(88) <= Q_88_EXMPLR ;
   Q(87) <= Q_87_EXMPLR ;
   Q(86) <= Q_86_EXMPLR ;
   Q(85) <= Q_85_EXMPLR ;
   Q(84) <= Q_84_EXMPLR ;
   Q(83) <= Q_83_EXMPLR ;
   Q(82) <= Q_82_EXMPLR ;
   Q(81) <= Q_81_EXMPLR ;
   Q(80) <= Q_80_EXMPLR ;
   Q(79) <= Q_79_EXMPLR ;
   Q(78) <= Q_78_EXMPLR ;
   Q(77) <= Q_77_EXMPLR ;
   Q(76) <= Q_76_EXMPLR ;
   Q(75) <= Q_75_EXMPLR ;
   Q(74) <= Q_74_EXMPLR ;
   Q(73) <= Q_73_EXMPLR ;
   Q(72) <= Q_72_EXMPLR ;
   Q(71) <= Q_71_EXMPLR ;
   Q(70) <= Q_70_EXMPLR ;
   Q(69) <= Q_69_EXMPLR ;
   Q(68) <= Q_68_EXMPLR ;
   Q(67) <= Q_67_EXMPLR ;
   Q(66) <= Q_66_EXMPLR ;
   Q(65) <= Q_65_EXMPLR ;
   Q(64) <= Q_64_EXMPLR ;
   Q(63) <= Q_63_EXMPLR ;
   Q(62) <= Q_62_EXMPLR ;
   Q(61) <= Q_61_EXMPLR ;
   Q(60) <= Q_60_EXMPLR ;
   Q(59) <= Q_59_EXMPLR ;
   Q(58) <= Q_58_EXMPLR ;
   Q(57) <= Q_57_EXMPLR ;
   Q(56) <= Q_56_EXMPLR ;
   Q(55) <= Q_55_EXMPLR ;
   Q(54) <= Q_54_EXMPLR ;
   Q(53) <= Q_53_EXMPLR ;
   Q(52) <= Q_52_EXMPLR ;
   Q(51) <= Q_51_EXMPLR ;
   Q(50) <= Q_50_EXMPLR ;
   Q(49) <= Q_49_EXMPLR ;
   Q(48) <= Q_48_EXMPLR ;
   Q(47) <= Q_47_EXMPLR ;
   Q(46) <= Q_46_EXMPLR ;
   Q(45) <= Q_45_EXMPLR ;
   Q(44) <= Q_44_EXMPLR ;
   Q(43) <= Q_43_EXMPLR ;
   Q(42) <= Q_42_EXMPLR ;
   Q(41) <= Q_41_EXMPLR ;
   Q(40) <= Q_40_EXMPLR ;
   Q(39) <= Q_39_EXMPLR ;
   Q(38) <= Q_38_EXMPLR ;
   Q(37) <= Q_37_EXMPLR ;
   Q(36) <= Q_36_EXMPLR ;
   Q(35) <= Q_35_EXMPLR ;
   Q(34) <= Q_34_EXMPLR ;
   Q(33) <= Q_33_EXMPLR ;
   Q(32) <= Q_32_EXMPLR ;
   Q(31) <= Q_31_EXMPLR ;
   Q(30) <= Q_30_EXMPLR ;
   Q(29) <= Q_29_EXMPLR ;
   Q(28) <= Q_28_EXMPLR ;
   Q(27) <= Q_27_EXMPLR ;
   Q(26) <= Q_26_EXMPLR ;
   Q(25) <= Q_25_EXMPLR ;
   Q(24) <= Q_24_EXMPLR ;
   Q(23) <= Q_23_EXMPLR ;
   Q(22) <= Q_22_EXMPLR ;
   Q(21) <= Q_21_EXMPLR ;
   Q(20) <= Q_20_EXMPLR ;
   Q(19) <= Q_19_EXMPLR ;
   Q(18) <= Q_18_EXMPLR ;
   Q(17) <= Q_17_EXMPLR ;
   Q(16) <= Q_16_EXMPLR ;
   Q(15) <= Q_15_EXMPLR ;
   Q(14) <= Q_14_EXMPLR ;
   Q(13) <= Q_13_EXMPLR ;
   Q(12) <= Q_12_EXMPLR ;
   Q(11) <= Q_11_EXMPLR ;
   Q(10) <= Q_10_EXMPLR ;
   Q(9) <= Q_9_EXMPLR ;
   Q(8) <= Q_8_EXMPLR ;
   Q(7) <= Q_7_EXMPLR ;
   Q(6) <= Q_6_EXMPLR ;
   Q(5) <= Q_5_EXMPLR ;
   Q(4) <= Q_4_EXMPLR ;
   Q(3) <= Q_3_EXMPLR ;
   Q(2) <= Q_2_EXMPLR ;
   Q(1) <= Q_1_EXMPLR ;
   Q(0) <= Q_0_EXMPLR ;
   reg_Q_0 : dffr port map ( Q=>Q_0_EXMPLR, QB=>OPEN, D=>nx4838, CLK=>
      nx10301, R=>RST);
   ix4839 : mux21_ni port map ( Y=>nx4838, A0=>Q_0_EXMPLR, A1=>D(0), S0=>
      nx10167);
   reg_Q_1 : dffr port map ( Q=>Q_1_EXMPLR, QB=>OPEN, D=>nx4848, CLK=>
      nx10301, R=>RST);
   ix4849 : mux21_ni port map ( Y=>nx4848, A0=>Q_1_EXMPLR, A1=>D(1), S0=>
      nx10167);
   reg_Q_2 : dffr port map ( Q=>Q_2_EXMPLR, QB=>OPEN, D=>nx4858, CLK=>
      nx10301, R=>RST);
   ix4859 : mux21_ni port map ( Y=>nx4858, A0=>Q_2_EXMPLR, A1=>D(2), S0=>
      nx10167);
   reg_Q_3 : dffr port map ( Q=>Q_3_EXMPLR, QB=>OPEN, D=>nx4868, CLK=>
      nx10301, R=>RST);
   ix4869 : mux21_ni port map ( Y=>nx4868, A0=>Q_3_EXMPLR, A1=>D(3), S0=>
      nx10167);
   reg_Q_4 : dffr port map ( Q=>Q_4_EXMPLR, QB=>OPEN, D=>nx4878, CLK=>
      nx10301, R=>RST);
   ix4879 : mux21_ni port map ( Y=>nx4878, A0=>Q_4_EXMPLR, A1=>D(4), S0=>
      nx10167);
   reg_Q_5 : dffr port map ( Q=>Q_5_EXMPLR, QB=>OPEN, D=>nx4888, CLK=>
      nx10301, R=>RST);
   ix4889 : mux21_ni port map ( Y=>nx4888, A0=>Q_5_EXMPLR, A1=>D(5), S0=>
      nx10167);
   reg_Q_6 : dffr port map ( Q=>Q_6_EXMPLR, QB=>OPEN, D=>nx4898, CLK=>
      nx10301, R=>RST);
   ix4899 : mux21_ni port map ( Y=>nx4898, A0=>Q_6_EXMPLR, A1=>D(6), S0=>
      nx10167);
   reg_Q_7 : dffr port map ( Q=>Q_7_EXMPLR, QB=>OPEN, D=>nx4908, CLK=>
      nx10047, R=>RST);
   ix4909 : mux21_ni port map ( Y=>nx4908, A0=>Q_7_EXMPLR, A1=>D(7), S0=>
      nx10169);
   reg_Q_8 : dffr port map ( Q=>Q_8_EXMPLR, QB=>OPEN, D=>nx4918, CLK=>
      nx10047, R=>RST);
   ix4919 : mux21_ni port map ( Y=>nx4918, A0=>Q_8_EXMPLR, A1=>D(8), S0=>
      nx10169);
   reg_Q_9 : dffr port map ( Q=>Q_9_EXMPLR, QB=>OPEN, D=>nx4928, CLK=>
      nx10047, R=>RST);
   ix4929 : mux21_ni port map ( Y=>nx4928, A0=>Q_9_EXMPLR, A1=>D(9), S0=>
      nx10169);
   reg_Q_10 : dffr port map ( Q=>Q_10_EXMPLR, QB=>OPEN, D=>nx4938, CLK=>
      nx10047, R=>RST);
   ix4939 : mux21_ni port map ( Y=>nx4938, A0=>Q_10_EXMPLR, A1=>D(10), S0=>
      nx10169);
   reg_Q_11 : dffr port map ( Q=>Q_11_EXMPLR, QB=>OPEN, D=>nx4948, CLK=>
      nx10047, R=>RST);
   ix4949 : mux21_ni port map ( Y=>nx4948, A0=>Q_11_EXMPLR, A1=>D(11), S0=>
      nx10169);
   reg_Q_12 : dffr port map ( Q=>Q_12_EXMPLR, QB=>OPEN, D=>nx4958, CLK=>
      nx10047, R=>RST);
   ix4959 : mux21_ni port map ( Y=>nx4958, A0=>Q_12_EXMPLR, A1=>D(12), S0=>
      nx10169);
   reg_Q_13 : dffr port map ( Q=>Q_13_EXMPLR, QB=>OPEN, D=>nx4968, CLK=>
      nx10047, R=>RST);
   ix4969 : mux21_ni port map ( Y=>nx4968, A0=>Q_13_EXMPLR, A1=>D(13), S0=>
      nx10169);
   reg_Q_14 : dffr port map ( Q=>Q_14_EXMPLR, QB=>OPEN, D=>nx4978, CLK=>
      nx10049, R=>RST);
   ix4979 : mux21_ni port map ( Y=>nx4978, A0=>Q_14_EXMPLR, A1=>D(14), S0=>
      nx10171);
   reg_Q_15 : dffr port map ( Q=>Q_15_EXMPLR, QB=>OPEN, D=>nx4988, CLK=>
      nx10049, R=>RST);
   ix4989 : mux21_ni port map ( Y=>nx4988, A0=>Q_15_EXMPLR, A1=>D(15), S0=>
      nx10171);
   reg_Q_16 : dffr port map ( Q=>Q_16_EXMPLR, QB=>OPEN, D=>nx4998, CLK=>
      nx10049, R=>RST);
   ix4999 : mux21_ni port map ( Y=>nx4998, A0=>Q_16_EXMPLR, A1=>D(16), S0=>
      nx10171);
   reg_Q_17 : dffr port map ( Q=>Q_17_EXMPLR, QB=>OPEN, D=>nx5008, CLK=>
      nx10049, R=>RST);
   ix5009 : mux21_ni port map ( Y=>nx5008, A0=>Q_17_EXMPLR, A1=>D(17), S0=>
      nx10171);
   reg_Q_18 : dffr port map ( Q=>Q_18_EXMPLR, QB=>OPEN, D=>nx5018, CLK=>
      nx10049, R=>RST);
   ix5019 : mux21_ni port map ( Y=>nx5018, A0=>Q_18_EXMPLR, A1=>D(18), S0=>
      nx10171);
   reg_Q_19 : dffr port map ( Q=>Q_19_EXMPLR, QB=>OPEN, D=>nx5028, CLK=>
      nx10049, R=>RST);
   ix5029 : mux21_ni port map ( Y=>nx5028, A0=>Q_19_EXMPLR, A1=>D(19), S0=>
      nx10171);
   reg_Q_20 : dffr port map ( Q=>Q_20_EXMPLR, QB=>OPEN, D=>nx5038, CLK=>
      nx10049, R=>RST);
   ix5039 : mux21_ni port map ( Y=>nx5038, A0=>Q_20_EXMPLR, A1=>D(20), S0=>
      nx10171);
   reg_Q_21 : dffr port map ( Q=>Q_21_EXMPLR, QB=>OPEN, D=>nx5048, CLK=>
      nx10051, R=>RST);
   ix5049 : mux21_ni port map ( Y=>nx5048, A0=>Q_21_EXMPLR, A1=>D(21), S0=>
      nx10173);
   reg_Q_22 : dffr port map ( Q=>Q_22_EXMPLR, QB=>OPEN, D=>nx5058, CLK=>
      nx10051, R=>RST);
   ix5059 : mux21_ni port map ( Y=>nx5058, A0=>Q_22_EXMPLR, A1=>D(22), S0=>
      nx10173);
   reg_Q_23 : dffr port map ( Q=>Q_23_EXMPLR, QB=>OPEN, D=>nx5068, CLK=>
      nx10051, R=>RST);
   ix5069 : mux21_ni port map ( Y=>nx5068, A0=>Q_23_EXMPLR, A1=>D(23), S0=>
      nx10173);
   reg_Q_24 : dffr port map ( Q=>Q_24_EXMPLR, QB=>OPEN, D=>nx5078, CLK=>
      nx10051, R=>RST);
   ix5079 : mux21_ni port map ( Y=>nx5078, A0=>Q_24_EXMPLR, A1=>D(24), S0=>
      nx10173);
   reg_Q_25 : dffr port map ( Q=>Q_25_EXMPLR, QB=>OPEN, D=>nx5088, CLK=>
      nx10051, R=>RST);
   ix5089 : mux21_ni port map ( Y=>nx5088, A0=>Q_25_EXMPLR, A1=>D(25), S0=>
      nx10173);
   reg_Q_26 : dffr port map ( Q=>Q_26_EXMPLR, QB=>OPEN, D=>nx5098, CLK=>
      nx10051, R=>RST);
   ix5099 : mux21_ni port map ( Y=>nx5098, A0=>Q_26_EXMPLR, A1=>D(26), S0=>
      nx10173);
   reg_Q_27 : dffr port map ( Q=>Q_27_EXMPLR, QB=>OPEN, D=>nx5108, CLK=>
      nx10051, R=>RST);
   ix5109 : mux21_ni port map ( Y=>nx5108, A0=>Q_27_EXMPLR, A1=>D(27), S0=>
      nx10173);
   reg_Q_28 : dffr port map ( Q=>Q_28_EXMPLR, QB=>OPEN, D=>nx5118, CLK=>
      nx10053, R=>RST);
   ix5119 : mux21_ni port map ( Y=>nx5118, A0=>Q_28_EXMPLR, A1=>D(28), S0=>
      nx10175);
   reg_Q_29 : dffr port map ( Q=>Q_29_EXMPLR, QB=>OPEN, D=>nx5128, CLK=>
      nx10053, R=>RST);
   ix5129 : mux21_ni port map ( Y=>nx5128, A0=>Q_29_EXMPLR, A1=>D(29), S0=>
      nx10175);
   reg_Q_30 : dffr port map ( Q=>Q_30_EXMPLR, QB=>OPEN, D=>nx5138, CLK=>
      nx10053, R=>RST);
   ix5139 : mux21_ni port map ( Y=>nx5138, A0=>Q_30_EXMPLR, A1=>D(30), S0=>
      nx10175);
   reg_Q_31 : dffr port map ( Q=>Q_31_EXMPLR, QB=>OPEN, D=>nx5148, CLK=>
      nx10053, R=>RST);
   ix5149 : mux21_ni port map ( Y=>nx5148, A0=>Q_31_EXMPLR, A1=>D(31), S0=>
      nx10175);
   reg_Q_32 : dffr port map ( Q=>Q_32_EXMPLR, QB=>OPEN, D=>nx5158, CLK=>
      nx10053, R=>RST);
   ix5159 : mux21_ni port map ( Y=>nx5158, A0=>Q_32_EXMPLR, A1=>D(32), S0=>
      nx10175);
   reg_Q_33 : dffr port map ( Q=>Q_33_EXMPLR, QB=>OPEN, D=>nx5168, CLK=>
      nx10053, R=>RST);
   ix5169 : mux21_ni port map ( Y=>nx5168, A0=>Q_33_EXMPLR, A1=>D(33), S0=>
      nx10175);
   reg_Q_34 : dffr port map ( Q=>Q_34_EXMPLR, QB=>OPEN, D=>nx5178, CLK=>
      nx10053, R=>RST);
   ix5179 : mux21_ni port map ( Y=>nx5178, A0=>Q_34_EXMPLR, A1=>D(34), S0=>
      nx10175);
   reg_Q_35 : dffr port map ( Q=>Q_35_EXMPLR, QB=>OPEN, D=>nx5188, CLK=>
      nx10055, R=>RST);
   ix5189 : mux21_ni port map ( Y=>nx5188, A0=>Q_35_EXMPLR, A1=>D(35), S0=>
      nx10177);
   reg_Q_36 : dffr port map ( Q=>Q_36_EXMPLR, QB=>OPEN, D=>nx5198, CLK=>
      nx10055, R=>RST);
   ix5199 : mux21_ni port map ( Y=>nx5198, A0=>Q_36_EXMPLR, A1=>D(36), S0=>
      nx10177);
   reg_Q_37 : dffr port map ( Q=>Q_37_EXMPLR, QB=>OPEN, D=>nx5208, CLK=>
      nx10055, R=>RST);
   ix5209 : mux21_ni port map ( Y=>nx5208, A0=>Q_37_EXMPLR, A1=>D(37), S0=>
      nx10177);
   reg_Q_38 : dffr port map ( Q=>Q_38_EXMPLR, QB=>OPEN, D=>nx5218, CLK=>
      nx10055, R=>RST);
   ix5219 : mux21_ni port map ( Y=>nx5218, A0=>Q_38_EXMPLR, A1=>D(38), S0=>
      nx10177);
   reg_Q_39 : dffr port map ( Q=>Q_39_EXMPLR, QB=>OPEN, D=>nx5228, CLK=>
      nx10055, R=>RST);
   ix5229 : mux21_ni port map ( Y=>nx5228, A0=>Q_39_EXMPLR, A1=>D(39), S0=>
      nx10177);
   reg_Q_40 : dffr port map ( Q=>Q_40_EXMPLR, QB=>OPEN, D=>nx5238, CLK=>
      nx10055, R=>RST);
   ix5239 : mux21_ni port map ( Y=>nx5238, A0=>Q_40_EXMPLR, A1=>D(40), S0=>
      nx10177);
   reg_Q_41 : dffr port map ( Q=>Q_41_EXMPLR, QB=>OPEN, D=>nx5248, CLK=>
      nx10055, R=>RST);
   ix5249 : mux21_ni port map ( Y=>nx5248, A0=>Q_41_EXMPLR, A1=>D(41), S0=>
      nx10177);
   reg_Q_42 : dffr port map ( Q=>Q_42_EXMPLR, QB=>OPEN, D=>nx5258, CLK=>
      nx10057, R=>RST);
   ix5259 : mux21_ni port map ( Y=>nx5258, A0=>Q_42_EXMPLR, A1=>D(42), S0=>
      nx10179);
   reg_Q_43 : dffr port map ( Q=>Q_43_EXMPLR, QB=>OPEN, D=>nx5268, CLK=>
      nx10057, R=>RST);
   ix5269 : mux21_ni port map ( Y=>nx5268, A0=>Q_43_EXMPLR, A1=>D(43), S0=>
      nx10179);
   reg_Q_44 : dffr port map ( Q=>Q_44_EXMPLR, QB=>OPEN, D=>nx5278, CLK=>
      nx10057, R=>RST);
   ix5279 : mux21_ni port map ( Y=>nx5278, A0=>Q_44_EXMPLR, A1=>D(44), S0=>
      nx10179);
   reg_Q_45 : dffr port map ( Q=>Q_45_EXMPLR, QB=>OPEN, D=>nx5288, CLK=>
      nx10057, R=>RST);
   ix5289 : mux21_ni port map ( Y=>nx5288, A0=>Q_45_EXMPLR, A1=>D(45), S0=>
      nx10179);
   reg_Q_46 : dffr port map ( Q=>Q_46_EXMPLR, QB=>OPEN, D=>nx5298, CLK=>
      nx10057, R=>RST);
   ix5299 : mux21_ni port map ( Y=>nx5298, A0=>Q_46_EXMPLR, A1=>D(46), S0=>
      nx10179);
   reg_Q_47 : dffr port map ( Q=>Q_47_EXMPLR, QB=>OPEN, D=>nx5308, CLK=>
      nx10057, R=>RST);
   ix5309 : mux21_ni port map ( Y=>nx5308, A0=>Q_47_EXMPLR, A1=>D(47), S0=>
      nx10179);
   reg_Q_48 : dffr port map ( Q=>Q_48_EXMPLR, QB=>OPEN, D=>nx5318, CLK=>
      nx10057, R=>RST);
   ix5319 : mux21_ni port map ( Y=>nx5318, A0=>Q_48_EXMPLR, A1=>D(48), S0=>
      nx10179);
   reg_Q_49 : dffr port map ( Q=>Q_49_EXMPLR, QB=>OPEN, D=>nx5328, CLK=>
      nx10059, R=>RST);
   ix5329 : mux21_ni port map ( Y=>nx5328, A0=>Q_49_EXMPLR, A1=>D(49), S0=>
      nx10181);
   reg_Q_50 : dffr port map ( Q=>Q_50_EXMPLR, QB=>OPEN, D=>nx5338, CLK=>
      nx10059, R=>RST);
   ix5339 : mux21_ni port map ( Y=>nx5338, A0=>Q_50_EXMPLR, A1=>D(50), S0=>
      nx10181);
   reg_Q_51 : dffr port map ( Q=>Q_51_EXMPLR, QB=>OPEN, D=>nx5348, CLK=>
      nx10059, R=>RST);
   ix5349 : mux21_ni port map ( Y=>nx5348, A0=>Q_51_EXMPLR, A1=>D(51), S0=>
      nx10181);
   reg_Q_52 : dffr port map ( Q=>Q_52_EXMPLR, QB=>OPEN, D=>nx5358, CLK=>
      nx10059, R=>RST);
   ix5359 : mux21_ni port map ( Y=>nx5358, A0=>Q_52_EXMPLR, A1=>D(52), S0=>
      nx10181);
   reg_Q_53 : dffr port map ( Q=>Q_53_EXMPLR, QB=>OPEN, D=>nx5368, CLK=>
      nx10059, R=>RST);
   ix5369 : mux21_ni port map ( Y=>nx5368, A0=>Q_53_EXMPLR, A1=>D(53), S0=>
      nx10181);
   reg_Q_54 : dffr port map ( Q=>Q_54_EXMPLR, QB=>OPEN, D=>nx5378, CLK=>
      nx10059, R=>RST);
   ix5379 : mux21_ni port map ( Y=>nx5378, A0=>Q_54_EXMPLR, A1=>D(54), S0=>
      nx10181);
   reg_Q_55 : dffr port map ( Q=>Q_55_EXMPLR, QB=>OPEN, D=>nx5388, CLK=>
      nx10059, R=>RST);
   ix5389 : mux21_ni port map ( Y=>nx5388, A0=>Q_55_EXMPLR, A1=>D(55), S0=>
      nx10181);
   reg_Q_56 : dffr port map ( Q=>Q_56_EXMPLR, QB=>OPEN, D=>nx5398, CLK=>
      nx10061, R=>RST);
   ix5399 : mux21_ni port map ( Y=>nx5398, A0=>Q_56_EXMPLR, A1=>D(56), S0=>
      nx10183);
   reg_Q_57 : dffr port map ( Q=>Q_57_EXMPLR, QB=>OPEN, D=>nx5408, CLK=>
      nx10061, R=>RST);
   ix5409 : mux21_ni port map ( Y=>nx5408, A0=>Q_57_EXMPLR, A1=>D(57), S0=>
      nx10183);
   reg_Q_58 : dffr port map ( Q=>Q_58_EXMPLR, QB=>OPEN, D=>nx5418, CLK=>
      nx10061, R=>RST);
   ix5419 : mux21_ni port map ( Y=>nx5418, A0=>Q_58_EXMPLR, A1=>D(58), S0=>
      nx10183);
   reg_Q_59 : dffr port map ( Q=>Q_59_EXMPLR, QB=>OPEN, D=>nx5428, CLK=>
      nx10061, R=>RST);
   ix5429 : mux21_ni port map ( Y=>nx5428, A0=>Q_59_EXMPLR, A1=>D(59), S0=>
      nx10183);
   reg_Q_60 : dffr port map ( Q=>Q_60_EXMPLR, QB=>OPEN, D=>nx5438, CLK=>
      nx10061, R=>RST);
   ix5439 : mux21_ni port map ( Y=>nx5438, A0=>Q_60_EXMPLR, A1=>D(60), S0=>
      nx10183);
   reg_Q_61 : dffr port map ( Q=>Q_61_EXMPLR, QB=>OPEN, D=>nx5448, CLK=>
      nx10061, R=>RST);
   ix5449 : mux21_ni port map ( Y=>nx5448, A0=>Q_61_EXMPLR, A1=>D(61), S0=>
      nx10183);
   reg_Q_62 : dffr port map ( Q=>Q_62_EXMPLR, QB=>OPEN, D=>nx5458, CLK=>
      nx10061, R=>RST);
   ix5459 : mux21_ni port map ( Y=>nx5458, A0=>Q_62_EXMPLR, A1=>D(62), S0=>
      nx10183);
   reg_Q_63 : dffr port map ( Q=>Q_63_EXMPLR, QB=>OPEN, D=>nx5468, CLK=>
      nx10063, R=>RST);
   ix5469 : mux21_ni port map ( Y=>nx5468, A0=>Q_63_EXMPLR, A1=>D(63), S0=>
      nx10185);
   reg_Q_64 : dffr port map ( Q=>Q_64_EXMPLR, QB=>OPEN, D=>nx5478, CLK=>
      nx10063, R=>RST);
   ix5479 : mux21_ni port map ( Y=>nx5478, A0=>Q_64_EXMPLR, A1=>D(64), S0=>
      nx10185);
   reg_Q_65 : dffr port map ( Q=>Q_65_EXMPLR, QB=>OPEN, D=>nx5488, CLK=>
      nx10063, R=>RST);
   ix5489 : mux21_ni port map ( Y=>nx5488, A0=>Q_65_EXMPLR, A1=>D(65), S0=>
      nx10185);
   reg_Q_66 : dffr port map ( Q=>Q_66_EXMPLR, QB=>OPEN, D=>nx5498, CLK=>
      nx10063, R=>RST);
   ix5499 : mux21_ni port map ( Y=>nx5498, A0=>Q_66_EXMPLR, A1=>D(66), S0=>
      nx10185);
   reg_Q_67 : dffr port map ( Q=>Q_67_EXMPLR, QB=>OPEN, D=>nx5508, CLK=>
      nx10063, R=>RST);
   ix5509 : mux21_ni port map ( Y=>nx5508, A0=>Q_67_EXMPLR, A1=>D(67), S0=>
      nx10185);
   reg_Q_68 : dffr port map ( Q=>Q_68_EXMPLR, QB=>OPEN, D=>nx5518, CLK=>
      nx10063, R=>RST);
   ix5519 : mux21_ni port map ( Y=>nx5518, A0=>Q_68_EXMPLR, A1=>D(68), S0=>
      nx10185);
   reg_Q_69 : dffr port map ( Q=>Q_69_EXMPLR, QB=>OPEN, D=>nx5528, CLK=>
      nx10063, R=>RST);
   ix5529 : mux21_ni port map ( Y=>nx5528, A0=>Q_69_EXMPLR, A1=>D(69), S0=>
      nx10185);
   reg_Q_70 : dffr port map ( Q=>Q_70_EXMPLR, QB=>OPEN, D=>nx5538, CLK=>
      nx10065, R=>RST);
   ix5539 : mux21_ni port map ( Y=>nx5538, A0=>Q_70_EXMPLR, A1=>D(70), S0=>
      nx10187);
   reg_Q_71 : dffr port map ( Q=>Q_71_EXMPLR, QB=>OPEN, D=>nx5548, CLK=>
      nx10065, R=>RST);
   ix5549 : mux21_ni port map ( Y=>nx5548, A0=>Q_71_EXMPLR, A1=>D(71), S0=>
      nx10187);
   reg_Q_72 : dffr port map ( Q=>Q_72_EXMPLR, QB=>OPEN, D=>nx5558, CLK=>
      nx10065, R=>RST);
   ix5559 : mux21_ni port map ( Y=>nx5558, A0=>Q_72_EXMPLR, A1=>D(72), S0=>
      nx10187);
   reg_Q_73 : dffr port map ( Q=>Q_73_EXMPLR, QB=>OPEN, D=>nx5568, CLK=>
      nx10065, R=>RST);
   ix5569 : mux21_ni port map ( Y=>nx5568, A0=>Q_73_EXMPLR, A1=>D(73), S0=>
      nx10187);
   reg_Q_74 : dffr port map ( Q=>Q_74_EXMPLR, QB=>OPEN, D=>nx5578, CLK=>
      nx10065, R=>RST);
   ix5579 : mux21_ni port map ( Y=>nx5578, A0=>Q_74_EXMPLR, A1=>D(74), S0=>
      nx10187);
   reg_Q_75 : dffr port map ( Q=>Q_75_EXMPLR, QB=>OPEN, D=>nx5588, CLK=>
      nx10065, R=>RST);
   ix5589 : mux21_ni port map ( Y=>nx5588, A0=>Q_75_EXMPLR, A1=>D(75), S0=>
      nx10187);
   reg_Q_76 : dffr port map ( Q=>Q_76_EXMPLR, QB=>OPEN, D=>nx5598, CLK=>
      nx10065, R=>RST);
   ix5599 : mux21_ni port map ( Y=>nx5598, A0=>Q_76_EXMPLR, A1=>D(76), S0=>
      nx10187);
   reg_Q_77 : dffr port map ( Q=>Q_77_EXMPLR, QB=>OPEN, D=>nx5608, CLK=>
      nx10067, R=>RST);
   ix5609 : mux21_ni port map ( Y=>nx5608, A0=>Q_77_EXMPLR, A1=>D(77), S0=>
      nx10189);
   reg_Q_78 : dffr port map ( Q=>Q_78_EXMPLR, QB=>OPEN, D=>nx5618, CLK=>
      nx10067, R=>RST);
   ix5619 : mux21_ni port map ( Y=>nx5618, A0=>Q_78_EXMPLR, A1=>D(78), S0=>
      nx10189);
   reg_Q_79 : dffr port map ( Q=>Q_79_EXMPLR, QB=>OPEN, D=>nx5628, CLK=>
      nx10067, R=>RST);
   ix5629 : mux21_ni port map ( Y=>nx5628, A0=>Q_79_EXMPLR, A1=>D(79), S0=>
      nx10189);
   reg_Q_80 : dffr port map ( Q=>Q_80_EXMPLR, QB=>OPEN, D=>nx5638, CLK=>
      nx10067, R=>RST);
   ix5639 : mux21_ni port map ( Y=>nx5638, A0=>Q_80_EXMPLR, A1=>D(80), S0=>
      nx10189);
   reg_Q_81 : dffr port map ( Q=>Q_81_EXMPLR, QB=>OPEN, D=>nx5648, CLK=>
      nx10067, R=>RST);
   ix5649 : mux21_ni port map ( Y=>nx5648, A0=>Q_81_EXMPLR, A1=>D(81), S0=>
      nx10189);
   reg_Q_82 : dffr port map ( Q=>Q_82_EXMPLR, QB=>OPEN, D=>nx5658, CLK=>
      nx10067, R=>RST);
   ix5659 : mux21_ni port map ( Y=>nx5658, A0=>Q_82_EXMPLR, A1=>D(82), S0=>
      nx10189);
   reg_Q_83 : dffr port map ( Q=>Q_83_EXMPLR, QB=>OPEN, D=>nx5668, CLK=>
      nx10067, R=>RST);
   ix5669 : mux21_ni port map ( Y=>nx5668, A0=>Q_83_EXMPLR, A1=>D(83), S0=>
      nx10189);
   reg_Q_84 : dffr port map ( Q=>Q_84_EXMPLR, QB=>OPEN, D=>nx5678, CLK=>
      nx10069, R=>RST);
   ix5679 : mux21_ni port map ( Y=>nx5678, A0=>Q_84_EXMPLR, A1=>D(84), S0=>
      nx10191);
   reg_Q_85 : dffr port map ( Q=>Q_85_EXMPLR, QB=>OPEN, D=>nx5688, CLK=>
      nx10069, R=>RST);
   ix5689 : mux21_ni port map ( Y=>nx5688, A0=>Q_85_EXMPLR, A1=>D(85), S0=>
      nx10191);
   reg_Q_86 : dffr port map ( Q=>Q_86_EXMPLR, QB=>OPEN, D=>nx5698, CLK=>
      nx10069, R=>RST);
   ix5699 : mux21_ni port map ( Y=>nx5698, A0=>Q_86_EXMPLR, A1=>D(86), S0=>
      nx10191);
   reg_Q_87 : dffr port map ( Q=>Q_87_EXMPLR, QB=>OPEN, D=>nx5708, CLK=>
      nx10069, R=>RST);
   ix5709 : mux21_ni port map ( Y=>nx5708, A0=>Q_87_EXMPLR, A1=>D(87), S0=>
      nx10191);
   reg_Q_88 : dffr port map ( Q=>Q_88_EXMPLR, QB=>OPEN, D=>nx5718, CLK=>
      nx10069, R=>RST);
   ix5719 : mux21_ni port map ( Y=>nx5718, A0=>Q_88_EXMPLR, A1=>D(88), S0=>
      nx10191);
   reg_Q_89 : dffr port map ( Q=>Q_89_EXMPLR, QB=>OPEN, D=>nx5728, CLK=>
      nx10069, R=>RST);
   ix5729 : mux21_ni port map ( Y=>nx5728, A0=>Q_89_EXMPLR, A1=>D(89), S0=>
      nx10191);
   reg_Q_90 : dffr port map ( Q=>Q_90_EXMPLR, QB=>OPEN, D=>nx5738, CLK=>
      nx10069, R=>RST);
   ix5739 : mux21_ni port map ( Y=>nx5738, A0=>Q_90_EXMPLR, A1=>D(90), S0=>
      nx10191);
   reg_Q_91 : dffr port map ( Q=>Q_91_EXMPLR, QB=>OPEN, D=>nx5748, CLK=>
      nx10071, R=>RST);
   ix5749 : mux21_ni port map ( Y=>nx5748, A0=>Q_91_EXMPLR, A1=>D(91), S0=>
      nx10193);
   reg_Q_92 : dffr port map ( Q=>Q_92_EXMPLR, QB=>OPEN, D=>nx5758, CLK=>
      nx10071, R=>RST);
   ix5759 : mux21_ni port map ( Y=>nx5758, A0=>Q_92_EXMPLR, A1=>D(92), S0=>
      nx10193);
   reg_Q_93 : dffr port map ( Q=>Q_93_EXMPLR, QB=>OPEN, D=>nx5768, CLK=>
      nx10071, R=>RST);
   ix5769 : mux21_ni port map ( Y=>nx5768, A0=>Q_93_EXMPLR, A1=>D(93), S0=>
      nx10193);
   reg_Q_94 : dffr port map ( Q=>Q_94_EXMPLR, QB=>OPEN, D=>nx5778, CLK=>
      nx10071, R=>RST);
   ix5779 : mux21_ni port map ( Y=>nx5778, A0=>Q_94_EXMPLR, A1=>D(94), S0=>
      nx10193);
   reg_Q_95 : dffr port map ( Q=>Q_95_EXMPLR, QB=>OPEN, D=>nx5788, CLK=>
      nx10071, R=>RST);
   ix5789 : mux21_ni port map ( Y=>nx5788, A0=>Q_95_EXMPLR, A1=>D(95), S0=>
      nx10193);
   reg_Q_96 : dffr port map ( Q=>Q_96_EXMPLR, QB=>OPEN, D=>nx5798, CLK=>
      nx10071, R=>RST);
   ix5799 : mux21_ni port map ( Y=>nx5798, A0=>Q_96_EXMPLR, A1=>D(96), S0=>
      nx10193);
   reg_Q_97 : dffr port map ( Q=>Q_97_EXMPLR, QB=>OPEN, D=>nx5808, CLK=>
      nx10071, R=>RST);
   ix5809 : mux21_ni port map ( Y=>nx5808, A0=>Q_97_EXMPLR, A1=>D(97), S0=>
      nx10193);
   reg_Q_98 : dffr port map ( Q=>Q_98_EXMPLR, QB=>OPEN, D=>nx5818, CLK=>
      nx10073, R=>RST);
   ix5819 : mux21_ni port map ( Y=>nx5818, A0=>Q_98_EXMPLR, A1=>D(98), S0=>
      nx10195);
   reg_Q_99 : dffr port map ( Q=>Q_99_EXMPLR, QB=>OPEN, D=>nx5828, CLK=>
      nx10073, R=>RST);
   ix5829 : mux21_ni port map ( Y=>nx5828, A0=>Q_99_EXMPLR, A1=>D(99), S0=>
      nx10195);
   reg_Q_100 : dffr port map ( Q=>Q_100_EXMPLR, QB=>OPEN, D=>nx5838, CLK=>
      nx10073, R=>RST);
   ix5839 : mux21_ni port map ( Y=>nx5838, A0=>Q_100_EXMPLR, A1=>D(100), S0
      =>nx10195);
   reg_Q_101 : dffr port map ( Q=>Q_101_EXMPLR, QB=>OPEN, D=>nx5848, CLK=>
      nx10073, R=>RST);
   ix5849 : mux21_ni port map ( Y=>nx5848, A0=>Q_101_EXMPLR, A1=>D(101), S0
      =>nx10195);
   reg_Q_102 : dffr port map ( Q=>Q_102_EXMPLR, QB=>OPEN, D=>nx5858, CLK=>
      nx10073, R=>RST);
   ix5859 : mux21_ni port map ( Y=>nx5858, A0=>Q_102_EXMPLR, A1=>D(102), S0
      =>nx10195);
   reg_Q_103 : dffr port map ( Q=>Q_103_EXMPLR, QB=>OPEN, D=>nx5868, CLK=>
      nx10073, R=>RST);
   ix5869 : mux21_ni port map ( Y=>nx5868, A0=>Q_103_EXMPLR, A1=>D(103), S0
      =>nx10195);
   reg_Q_104 : dffr port map ( Q=>Q_104_EXMPLR, QB=>OPEN, D=>nx5878, CLK=>
      nx10073, R=>RST);
   ix5879 : mux21_ni port map ( Y=>nx5878, A0=>Q_104_EXMPLR, A1=>D(104), S0
      =>nx10195);
   reg_Q_105 : dffr port map ( Q=>Q_105_EXMPLR, QB=>OPEN, D=>nx5888, CLK=>
      nx10075, R=>RST);
   ix5889 : mux21_ni port map ( Y=>nx5888, A0=>Q_105_EXMPLR, A1=>D(105), S0
      =>nx10197);
   reg_Q_106 : dffr port map ( Q=>Q_106_EXMPLR, QB=>OPEN, D=>nx5898, CLK=>
      nx10075, R=>RST);
   ix5899 : mux21_ni port map ( Y=>nx5898, A0=>Q_106_EXMPLR, A1=>D(106), S0
      =>nx10197);
   reg_Q_107 : dffr port map ( Q=>Q_107_EXMPLR, QB=>OPEN, D=>nx5908, CLK=>
      nx10075, R=>RST);
   ix5909 : mux21_ni port map ( Y=>nx5908, A0=>Q_107_EXMPLR, A1=>D(107), S0
      =>nx10197);
   reg_Q_108 : dffr port map ( Q=>Q_108_EXMPLR, QB=>OPEN, D=>nx5918, CLK=>
      nx10075, R=>RST);
   ix5919 : mux21_ni port map ( Y=>nx5918, A0=>Q_108_EXMPLR, A1=>D(108), S0
      =>nx10197);
   reg_Q_109 : dffr port map ( Q=>Q_109_EXMPLR, QB=>OPEN, D=>nx5928, CLK=>
      nx10075, R=>RST);
   ix5929 : mux21_ni port map ( Y=>nx5928, A0=>Q_109_EXMPLR, A1=>D(109), S0
      =>nx10197);
   reg_Q_110 : dffr port map ( Q=>Q_110_EXMPLR, QB=>OPEN, D=>nx5938, CLK=>
      nx10075, R=>RST);
   ix5939 : mux21_ni port map ( Y=>nx5938, A0=>Q_110_EXMPLR, A1=>D(110), S0
      =>nx10197);
   reg_Q_111 : dffr port map ( Q=>Q_111_EXMPLR, QB=>OPEN, D=>nx5948, CLK=>
      nx10075, R=>RST);
   ix5949 : mux21_ni port map ( Y=>nx5948, A0=>Q_111_EXMPLR, A1=>D(111), S0
      =>nx10197);
   reg_Q_112 : dffr port map ( Q=>Q_112_EXMPLR, QB=>OPEN, D=>nx5958, CLK=>
      nx10077, R=>RST);
   ix5959 : mux21_ni port map ( Y=>nx5958, A0=>Q_112_EXMPLR, A1=>D(112), S0
      =>nx10199);
   reg_Q_113 : dffr port map ( Q=>Q_113_EXMPLR, QB=>OPEN, D=>nx5968, CLK=>
      nx10077, R=>RST);
   ix5969 : mux21_ni port map ( Y=>nx5968, A0=>Q_113_EXMPLR, A1=>D(113), S0
      =>nx10199);
   reg_Q_114 : dffr port map ( Q=>Q_114_EXMPLR, QB=>OPEN, D=>nx5978, CLK=>
      nx10077, R=>RST);
   ix5979 : mux21_ni port map ( Y=>nx5978, A0=>Q_114_EXMPLR, A1=>D(114), S0
      =>nx10199);
   reg_Q_115 : dffr port map ( Q=>Q_115_EXMPLR, QB=>OPEN, D=>nx5988, CLK=>
      nx10077, R=>RST);
   ix5989 : mux21_ni port map ( Y=>nx5988, A0=>Q_115_EXMPLR, A1=>D(115), S0
      =>nx10199);
   reg_Q_116 : dffr port map ( Q=>Q_116_EXMPLR, QB=>OPEN, D=>nx5998, CLK=>
      nx10077, R=>RST);
   ix5999 : mux21_ni port map ( Y=>nx5998, A0=>Q_116_EXMPLR, A1=>D(116), S0
      =>nx10199);
   reg_Q_117 : dffr port map ( Q=>Q_117_EXMPLR, QB=>OPEN, D=>nx6008, CLK=>
      nx10077, R=>RST);
   ix6009 : mux21_ni port map ( Y=>nx6008, A0=>Q_117_EXMPLR, A1=>D(117), S0
      =>nx10199);
   reg_Q_118 : dffr port map ( Q=>Q_118_EXMPLR, QB=>OPEN, D=>nx6018, CLK=>
      nx10077, R=>RST);
   ix6019 : mux21_ni port map ( Y=>nx6018, A0=>Q_118_EXMPLR, A1=>D(118), S0
      =>nx10199);
   reg_Q_119 : dffr port map ( Q=>Q_119_EXMPLR, QB=>OPEN, D=>nx6028, CLK=>
      nx10079, R=>RST);
   ix6029 : mux21_ni port map ( Y=>nx6028, A0=>Q_119_EXMPLR, A1=>D(119), S0
      =>nx10201);
   reg_Q_120 : dffr port map ( Q=>Q_120_EXMPLR, QB=>OPEN, D=>nx6038, CLK=>
      nx10079, R=>RST);
   ix6039 : mux21_ni port map ( Y=>nx6038, A0=>Q_120_EXMPLR, A1=>D(120), S0
      =>nx10201);
   reg_Q_121 : dffr port map ( Q=>Q_121_EXMPLR, QB=>OPEN, D=>nx6048, CLK=>
      nx10079, R=>RST);
   ix6049 : mux21_ni port map ( Y=>nx6048, A0=>Q_121_EXMPLR, A1=>D(121), S0
      =>nx10201);
   reg_Q_122 : dffr port map ( Q=>Q_122_EXMPLR, QB=>OPEN, D=>nx6058, CLK=>
      nx10079, R=>RST);
   ix6059 : mux21_ni port map ( Y=>nx6058, A0=>Q_122_EXMPLR, A1=>D(122), S0
      =>nx10201);
   reg_Q_123 : dffr port map ( Q=>Q_123_EXMPLR, QB=>OPEN, D=>nx6068, CLK=>
      nx10079, R=>RST);
   ix6069 : mux21_ni port map ( Y=>nx6068, A0=>Q_123_EXMPLR, A1=>D(123), S0
      =>nx10201);
   reg_Q_124 : dffr port map ( Q=>Q_124_EXMPLR, QB=>OPEN, D=>nx6078, CLK=>
      nx10079, R=>RST);
   ix6079 : mux21_ni port map ( Y=>nx6078, A0=>Q_124_EXMPLR, A1=>D(124), S0
      =>nx10201);
   reg_Q_125 : dffr port map ( Q=>Q_125_EXMPLR, QB=>OPEN, D=>nx6088, CLK=>
      nx10079, R=>RST);
   ix6089 : mux21_ni port map ( Y=>nx6088, A0=>Q_125_EXMPLR, A1=>D(125), S0
      =>nx10201);
   reg_Q_126 : dffr port map ( Q=>Q_126_EXMPLR, QB=>OPEN, D=>nx6098, CLK=>
      nx10081, R=>RST);
   ix6099 : mux21_ni port map ( Y=>nx6098, A0=>Q_126_EXMPLR, A1=>D(126), S0
      =>nx10203);
   reg_Q_127 : dffr port map ( Q=>Q_127_EXMPLR, QB=>OPEN, D=>nx6108, CLK=>
      nx10081, R=>RST);
   ix6109 : mux21_ni port map ( Y=>nx6108, A0=>Q_127_EXMPLR, A1=>D(127), S0
      =>nx10203);
   reg_Q_128 : dffr port map ( Q=>Q_128_EXMPLR, QB=>OPEN, D=>nx6118, CLK=>
      nx10081, R=>RST);
   ix6119 : mux21_ni port map ( Y=>nx6118, A0=>Q_128_EXMPLR, A1=>D(128), S0
      =>nx10203);
   reg_Q_129 : dffr port map ( Q=>Q_129_EXMPLR, QB=>OPEN, D=>nx6128, CLK=>
      nx10081, R=>RST);
   ix6129 : mux21_ni port map ( Y=>nx6128, A0=>Q_129_EXMPLR, A1=>D(129), S0
      =>nx10203);
   reg_Q_130 : dffr port map ( Q=>Q_130_EXMPLR, QB=>OPEN, D=>nx6138, CLK=>
      nx10081, R=>RST);
   ix6139 : mux21_ni port map ( Y=>nx6138, A0=>Q_130_EXMPLR, A1=>D(130), S0
      =>nx10203);
   reg_Q_131 : dffr port map ( Q=>Q_131_EXMPLR, QB=>OPEN, D=>nx6148, CLK=>
      nx10081, R=>RST);
   ix6149 : mux21_ni port map ( Y=>nx6148, A0=>Q_131_EXMPLR, A1=>D(131), S0
      =>nx10203);
   reg_Q_132 : dffr port map ( Q=>Q_132_EXMPLR, QB=>OPEN, D=>nx6158, CLK=>
      nx10081, R=>RST);
   ix6159 : mux21_ni port map ( Y=>nx6158, A0=>Q_132_EXMPLR, A1=>D(132), S0
      =>nx10203);
   reg_Q_133 : dffr port map ( Q=>Q_133_EXMPLR, QB=>OPEN, D=>nx6168, CLK=>
      nx10083, R=>RST);
   ix6169 : mux21_ni port map ( Y=>nx6168, A0=>Q_133_EXMPLR, A1=>D(133), S0
      =>nx10205);
   reg_Q_134 : dffr port map ( Q=>Q_134_EXMPLR, QB=>OPEN, D=>nx6178, CLK=>
      nx10083, R=>RST);
   ix6179 : mux21_ni port map ( Y=>nx6178, A0=>Q_134_EXMPLR, A1=>D(134), S0
      =>nx10205);
   reg_Q_135 : dffr port map ( Q=>Q_135_EXMPLR, QB=>OPEN, D=>nx6188, CLK=>
      nx10083, R=>RST);
   ix6189 : mux21_ni port map ( Y=>nx6188, A0=>Q_135_EXMPLR, A1=>D(135), S0
      =>nx10205);
   reg_Q_136 : dffr port map ( Q=>Q_136_EXMPLR, QB=>OPEN, D=>nx6198, CLK=>
      nx10083, R=>RST);
   ix6199 : mux21_ni port map ( Y=>nx6198, A0=>Q_136_EXMPLR, A1=>D(136), S0
      =>nx10205);
   reg_Q_137 : dffr port map ( Q=>Q_137_EXMPLR, QB=>OPEN, D=>nx6208, CLK=>
      nx10083, R=>RST);
   ix6209 : mux21_ni port map ( Y=>nx6208, A0=>Q_137_EXMPLR, A1=>D(137), S0
      =>nx10205);
   reg_Q_138 : dffr port map ( Q=>Q_138_EXMPLR, QB=>OPEN, D=>nx6218, CLK=>
      nx10083, R=>RST);
   ix6219 : mux21_ni port map ( Y=>nx6218, A0=>Q_138_EXMPLR, A1=>D(138), S0
      =>nx10205);
   reg_Q_139 : dffr port map ( Q=>Q_139_EXMPLR, QB=>OPEN, D=>nx6228, CLK=>
      nx10083, R=>RST);
   ix6229 : mux21_ni port map ( Y=>nx6228, A0=>Q_139_EXMPLR, A1=>D(139), S0
      =>nx10205);
   reg_Q_140 : dffr port map ( Q=>Q_140_EXMPLR, QB=>OPEN, D=>nx6238, CLK=>
      nx10085, R=>RST);
   ix6239 : mux21_ni port map ( Y=>nx6238, A0=>Q_140_EXMPLR, A1=>D(140), S0
      =>nx10207);
   reg_Q_141 : dffr port map ( Q=>Q_141_EXMPLR, QB=>OPEN, D=>nx6248, CLK=>
      nx10085, R=>RST);
   ix6249 : mux21_ni port map ( Y=>nx6248, A0=>Q_141_EXMPLR, A1=>D(141), S0
      =>nx10207);
   reg_Q_142 : dffr port map ( Q=>Q_142_EXMPLR, QB=>OPEN, D=>nx6258, CLK=>
      nx10085, R=>RST);
   ix6259 : mux21_ni port map ( Y=>nx6258, A0=>Q_142_EXMPLR, A1=>D(142), S0
      =>nx10207);
   reg_Q_143 : dffr port map ( Q=>Q_143_EXMPLR, QB=>OPEN, D=>nx6268, CLK=>
      nx10085, R=>RST);
   ix6269 : mux21_ni port map ( Y=>nx6268, A0=>Q_143_EXMPLR, A1=>D(143), S0
      =>nx10207);
   reg_Q_144 : dffr port map ( Q=>Q_144_EXMPLR, QB=>OPEN, D=>nx6278, CLK=>
      nx10085, R=>RST);
   ix6279 : mux21_ni port map ( Y=>nx6278, A0=>Q_144_EXMPLR, A1=>D(144), S0
      =>nx10207);
   reg_Q_145 : dffr port map ( Q=>Q_145_EXMPLR, QB=>OPEN, D=>nx6288, CLK=>
      nx10085, R=>RST);
   ix6289 : mux21_ni port map ( Y=>nx6288, A0=>Q_145_EXMPLR, A1=>D(145), S0
      =>nx10207);
   reg_Q_146 : dffr port map ( Q=>Q_146_EXMPLR, QB=>OPEN, D=>nx6298, CLK=>
      nx10085, R=>RST);
   ix6299 : mux21_ni port map ( Y=>nx6298, A0=>Q_146_EXMPLR, A1=>D(146), S0
      =>nx10207);
   reg_Q_147 : dffr port map ( Q=>Q_147_EXMPLR, QB=>OPEN, D=>nx6308, CLK=>
      nx10087, R=>RST);
   ix6309 : mux21_ni port map ( Y=>nx6308, A0=>Q_147_EXMPLR, A1=>D(147), S0
      =>nx10209);
   reg_Q_148 : dffr port map ( Q=>Q_148_EXMPLR, QB=>OPEN, D=>nx6318, CLK=>
      nx10087, R=>RST);
   ix6319 : mux21_ni port map ( Y=>nx6318, A0=>Q_148_EXMPLR, A1=>D(148), S0
      =>nx10209);
   reg_Q_149 : dffr port map ( Q=>Q_149_EXMPLR, QB=>OPEN, D=>nx6328, CLK=>
      nx10087, R=>RST);
   ix6329 : mux21_ni port map ( Y=>nx6328, A0=>Q_149_EXMPLR, A1=>D(149), S0
      =>nx10209);
   reg_Q_150 : dffr port map ( Q=>Q_150_EXMPLR, QB=>OPEN, D=>nx6338, CLK=>
      nx10087, R=>RST);
   ix6339 : mux21_ni port map ( Y=>nx6338, A0=>Q_150_EXMPLR, A1=>D(150), S0
      =>nx10209);
   reg_Q_151 : dffr port map ( Q=>Q_151_EXMPLR, QB=>OPEN, D=>nx6348, CLK=>
      nx10087, R=>RST);
   ix6349 : mux21_ni port map ( Y=>nx6348, A0=>Q_151_EXMPLR, A1=>D(151), S0
      =>nx10209);
   reg_Q_152 : dffr port map ( Q=>Q_152_EXMPLR, QB=>OPEN, D=>nx6358, CLK=>
      nx10087, R=>RST);
   ix6359 : mux21_ni port map ( Y=>nx6358, A0=>Q_152_EXMPLR, A1=>D(152), S0
      =>nx10209);
   reg_Q_153 : dffr port map ( Q=>Q_153_EXMPLR, QB=>OPEN, D=>nx6368, CLK=>
      nx10087, R=>RST);
   ix6369 : mux21_ni port map ( Y=>nx6368, A0=>Q_153_EXMPLR, A1=>D(153), S0
      =>nx10209);
   reg_Q_154 : dffr port map ( Q=>Q_154_EXMPLR, QB=>OPEN, D=>nx6378, CLK=>
      nx10089, R=>RST);
   ix6379 : mux21_ni port map ( Y=>nx6378, A0=>Q_154_EXMPLR, A1=>D(154), S0
      =>nx10211);
   reg_Q_155 : dffr port map ( Q=>Q_155_EXMPLR, QB=>OPEN, D=>nx6388, CLK=>
      nx10089, R=>RST);
   ix6389 : mux21_ni port map ( Y=>nx6388, A0=>Q_155_EXMPLR, A1=>D(155), S0
      =>nx10211);
   reg_Q_156 : dffr port map ( Q=>Q_156_EXMPLR, QB=>OPEN, D=>nx6398, CLK=>
      nx10089, R=>RST);
   ix6399 : mux21_ni port map ( Y=>nx6398, A0=>Q_156_EXMPLR, A1=>D(156), S0
      =>nx10211);
   reg_Q_157 : dffr port map ( Q=>Q_157_EXMPLR, QB=>OPEN, D=>nx6408, CLK=>
      nx10089, R=>RST);
   ix6409 : mux21_ni port map ( Y=>nx6408, A0=>Q_157_EXMPLR, A1=>D(157), S0
      =>nx10211);
   reg_Q_158 : dffr port map ( Q=>Q_158_EXMPLR, QB=>OPEN, D=>nx6418, CLK=>
      nx10089, R=>RST);
   ix6419 : mux21_ni port map ( Y=>nx6418, A0=>Q_158_EXMPLR, A1=>D(158), S0
      =>nx10211);
   reg_Q_159 : dffr port map ( Q=>Q_159_EXMPLR, QB=>OPEN, D=>nx6428, CLK=>
      nx10089, R=>RST);
   ix6429 : mux21_ni port map ( Y=>nx6428, A0=>Q_159_EXMPLR, A1=>D(159), S0
      =>nx10211);
   reg_Q_160 : dffr port map ( Q=>Q_160_EXMPLR, QB=>OPEN, D=>nx6438, CLK=>
      nx10089, R=>RST);
   ix6439 : mux21_ni port map ( Y=>nx6438, A0=>Q_160_EXMPLR, A1=>D(160), S0
      =>nx10211);
   reg_Q_161 : dffr port map ( Q=>Q_161_EXMPLR, QB=>OPEN, D=>nx6448, CLK=>
      nx10091, R=>RST);
   ix6449 : mux21_ni port map ( Y=>nx6448, A0=>Q_161_EXMPLR, A1=>D(161), S0
      =>nx10213);
   reg_Q_162 : dffr port map ( Q=>Q_162_EXMPLR, QB=>OPEN, D=>nx6458, CLK=>
      nx10091, R=>RST);
   ix6459 : mux21_ni port map ( Y=>nx6458, A0=>Q_162_EXMPLR, A1=>D(162), S0
      =>nx10213);
   reg_Q_163 : dffr port map ( Q=>Q_163_EXMPLR, QB=>OPEN, D=>nx6468, CLK=>
      nx10091, R=>RST);
   ix6469 : mux21_ni port map ( Y=>nx6468, A0=>Q_163_EXMPLR, A1=>D(163), S0
      =>nx10213);
   reg_Q_164 : dffr port map ( Q=>Q_164_EXMPLR, QB=>OPEN, D=>nx6478, CLK=>
      nx10091, R=>RST);
   ix6479 : mux21_ni port map ( Y=>nx6478, A0=>Q_164_EXMPLR, A1=>D(164), S0
      =>nx10213);
   reg_Q_165 : dffr port map ( Q=>Q_165_EXMPLR, QB=>OPEN, D=>nx6488, CLK=>
      nx10091, R=>RST);
   ix6489 : mux21_ni port map ( Y=>nx6488, A0=>Q_165_EXMPLR, A1=>D(165), S0
      =>nx10213);
   reg_Q_166 : dffr port map ( Q=>Q_166_EXMPLR, QB=>OPEN, D=>nx6498, CLK=>
      nx10091, R=>RST);
   ix6499 : mux21_ni port map ( Y=>nx6498, A0=>Q_166_EXMPLR, A1=>D(166), S0
      =>nx10213);
   reg_Q_167 : dffr port map ( Q=>Q_167_EXMPLR, QB=>OPEN, D=>nx6508, CLK=>
      nx10091, R=>RST);
   ix6509 : mux21_ni port map ( Y=>nx6508, A0=>Q_167_EXMPLR, A1=>D(167), S0
      =>nx10213);
   reg_Q_168 : dffr port map ( Q=>Q_168_EXMPLR, QB=>OPEN, D=>nx6518, CLK=>
      nx10093, R=>RST);
   ix6519 : mux21_ni port map ( Y=>nx6518, A0=>Q_168_EXMPLR, A1=>D(168), S0
      =>nx10215);
   reg_Q_169 : dffr port map ( Q=>Q_169_EXMPLR, QB=>OPEN, D=>nx6528, CLK=>
      nx10093, R=>RST);
   ix6529 : mux21_ni port map ( Y=>nx6528, A0=>Q_169_EXMPLR, A1=>D(169), S0
      =>nx10215);
   reg_Q_170 : dffr port map ( Q=>Q_170_EXMPLR, QB=>OPEN, D=>nx6538, CLK=>
      nx10093, R=>RST);
   ix6539 : mux21_ni port map ( Y=>nx6538, A0=>Q_170_EXMPLR, A1=>D(170), S0
      =>nx10215);
   reg_Q_171 : dffr port map ( Q=>Q_171_EXMPLR, QB=>OPEN, D=>nx6548, CLK=>
      nx10093, R=>RST);
   ix6549 : mux21_ni port map ( Y=>nx6548, A0=>Q_171_EXMPLR, A1=>D(171), S0
      =>nx10215);
   reg_Q_172 : dffr port map ( Q=>Q_172_EXMPLR, QB=>OPEN, D=>nx6558, CLK=>
      nx10093, R=>RST);
   ix6559 : mux21_ni port map ( Y=>nx6558, A0=>Q_172_EXMPLR, A1=>D(172), S0
      =>nx10215);
   reg_Q_173 : dffr port map ( Q=>Q_173_EXMPLR, QB=>OPEN, D=>nx6568, CLK=>
      nx10093, R=>RST);
   ix6569 : mux21_ni port map ( Y=>nx6568, A0=>Q_173_EXMPLR, A1=>D(173), S0
      =>nx10215);
   reg_Q_174 : dffr port map ( Q=>Q_174_EXMPLR, QB=>OPEN, D=>nx6578, CLK=>
      nx10093, R=>RST);
   ix6579 : mux21_ni port map ( Y=>nx6578, A0=>Q_174_EXMPLR, A1=>D(174), S0
      =>nx10215);
   reg_Q_175 : dffr port map ( Q=>Q_175_EXMPLR, QB=>OPEN, D=>nx6588, CLK=>
      nx10095, R=>RST);
   ix6589 : mux21_ni port map ( Y=>nx6588, A0=>Q_175_EXMPLR, A1=>D(175), S0
      =>nx10217);
   reg_Q_176 : dffr port map ( Q=>Q_176_EXMPLR, QB=>OPEN, D=>nx6598, CLK=>
      nx10095, R=>RST);
   ix6599 : mux21_ni port map ( Y=>nx6598, A0=>Q_176_EXMPLR, A1=>D(176), S0
      =>nx10217);
   reg_Q_177 : dffr port map ( Q=>Q_177_EXMPLR, QB=>OPEN, D=>nx6608, CLK=>
      nx10095, R=>RST);
   ix6609 : mux21_ni port map ( Y=>nx6608, A0=>Q_177_EXMPLR, A1=>D(177), S0
      =>nx10217);
   reg_Q_178 : dffr port map ( Q=>Q_178_EXMPLR, QB=>OPEN, D=>nx6618, CLK=>
      nx10095, R=>RST);
   ix6619 : mux21_ni port map ( Y=>nx6618, A0=>Q_178_EXMPLR, A1=>D(178), S0
      =>nx10217);
   reg_Q_179 : dffr port map ( Q=>Q_179_EXMPLR, QB=>OPEN, D=>nx6628, CLK=>
      nx10095, R=>RST);
   ix6629 : mux21_ni port map ( Y=>nx6628, A0=>Q_179_EXMPLR, A1=>D(179), S0
      =>nx10217);
   reg_Q_180 : dffr port map ( Q=>Q_180_EXMPLR, QB=>OPEN, D=>nx6638, CLK=>
      nx10095, R=>RST);
   ix6639 : mux21_ni port map ( Y=>nx6638, A0=>Q_180_EXMPLR, A1=>D(180), S0
      =>nx10217);
   reg_Q_181 : dffr port map ( Q=>Q_181_EXMPLR, QB=>OPEN, D=>nx6648, CLK=>
      nx10095, R=>RST);
   ix6649 : mux21_ni port map ( Y=>nx6648, A0=>Q_181_EXMPLR, A1=>D(181), S0
      =>nx10217);
   reg_Q_182 : dffr port map ( Q=>Q_182_EXMPLR, QB=>OPEN, D=>nx6658, CLK=>
      nx10097, R=>RST);
   ix6659 : mux21_ni port map ( Y=>nx6658, A0=>Q_182_EXMPLR, A1=>D(182), S0
      =>nx10219);
   reg_Q_183 : dffr port map ( Q=>Q_183_EXMPLR, QB=>OPEN, D=>nx6668, CLK=>
      nx10097, R=>RST);
   ix6669 : mux21_ni port map ( Y=>nx6668, A0=>Q_183_EXMPLR, A1=>D(183), S0
      =>nx10219);
   reg_Q_184 : dffr port map ( Q=>Q_184_EXMPLR, QB=>OPEN, D=>nx6678, CLK=>
      nx10097, R=>RST);
   ix6679 : mux21_ni port map ( Y=>nx6678, A0=>Q_184_EXMPLR, A1=>D(184), S0
      =>nx10219);
   reg_Q_185 : dffr port map ( Q=>Q_185_EXMPLR, QB=>OPEN, D=>nx6688, CLK=>
      nx10097, R=>RST);
   ix6689 : mux21_ni port map ( Y=>nx6688, A0=>Q_185_EXMPLR, A1=>D(185), S0
      =>nx10219);
   reg_Q_186 : dffr port map ( Q=>Q_186_EXMPLR, QB=>OPEN, D=>nx6698, CLK=>
      nx10097, R=>RST);
   ix6699 : mux21_ni port map ( Y=>nx6698, A0=>Q_186_EXMPLR, A1=>D(186), S0
      =>nx10219);
   reg_Q_187 : dffr port map ( Q=>Q_187_EXMPLR, QB=>OPEN, D=>nx6708, CLK=>
      nx10097, R=>RST);
   ix6709 : mux21_ni port map ( Y=>nx6708, A0=>Q_187_EXMPLR, A1=>D(187), S0
      =>nx10219);
   reg_Q_188 : dffr port map ( Q=>Q_188_EXMPLR, QB=>OPEN, D=>nx6718, CLK=>
      nx10097, R=>RST);
   ix6719 : mux21_ni port map ( Y=>nx6718, A0=>Q_188_EXMPLR, A1=>D(188), S0
      =>nx10219);
   reg_Q_189 : dffr port map ( Q=>Q_189_EXMPLR, QB=>OPEN, D=>nx6728, CLK=>
      nx10099, R=>RST);
   ix6729 : mux21_ni port map ( Y=>nx6728, A0=>Q_189_EXMPLR, A1=>D(189), S0
      =>nx10221);
   reg_Q_190 : dffr port map ( Q=>Q_190_EXMPLR, QB=>OPEN, D=>nx6738, CLK=>
      nx10099, R=>RST);
   ix6739 : mux21_ni port map ( Y=>nx6738, A0=>Q_190_EXMPLR, A1=>D(190), S0
      =>nx10221);
   reg_Q_191 : dffr port map ( Q=>Q_191_EXMPLR, QB=>OPEN, D=>nx6748, CLK=>
      nx10099, R=>RST);
   ix6749 : mux21_ni port map ( Y=>nx6748, A0=>Q_191_EXMPLR, A1=>D(191), S0
      =>nx10221);
   reg_Q_192 : dffr port map ( Q=>Q_192_EXMPLR, QB=>OPEN, D=>nx6758, CLK=>
      nx10099, R=>RST);
   ix6759 : mux21_ni port map ( Y=>nx6758, A0=>Q_192_EXMPLR, A1=>D(192), S0
      =>nx10221);
   reg_Q_193 : dffr port map ( Q=>Q_193_EXMPLR, QB=>OPEN, D=>nx6768, CLK=>
      nx10099, R=>RST);
   ix6769 : mux21_ni port map ( Y=>nx6768, A0=>Q_193_EXMPLR, A1=>D(193), S0
      =>nx10221);
   reg_Q_194 : dffr port map ( Q=>Q_194_EXMPLR, QB=>OPEN, D=>nx6778, CLK=>
      nx10099, R=>RST);
   ix6779 : mux21_ni port map ( Y=>nx6778, A0=>Q_194_EXMPLR, A1=>D(194), S0
      =>nx10221);
   reg_Q_195 : dffr port map ( Q=>Q_195_EXMPLR, QB=>OPEN, D=>nx6788, CLK=>
      nx10099, R=>RST);
   ix6789 : mux21_ni port map ( Y=>nx6788, A0=>Q_195_EXMPLR, A1=>D(195), S0
      =>nx10221);
   reg_Q_196 : dffr port map ( Q=>Q_196_EXMPLR, QB=>OPEN, D=>nx6798, CLK=>
      nx10101, R=>RST);
   ix6799 : mux21_ni port map ( Y=>nx6798, A0=>Q_196_EXMPLR, A1=>D(196), S0
      =>nx10223);
   reg_Q_197 : dffr port map ( Q=>Q_197_EXMPLR, QB=>OPEN, D=>nx6808, CLK=>
      nx10101, R=>RST);
   ix6809 : mux21_ni port map ( Y=>nx6808, A0=>Q_197_EXMPLR, A1=>D(197), S0
      =>nx10223);
   reg_Q_198 : dffr port map ( Q=>Q_198_EXMPLR, QB=>OPEN, D=>nx6818, CLK=>
      nx10101, R=>RST);
   ix6819 : mux21_ni port map ( Y=>nx6818, A0=>Q_198_EXMPLR, A1=>D(198), S0
      =>nx10223);
   reg_Q_199 : dffr port map ( Q=>Q_199_EXMPLR, QB=>OPEN, D=>nx6828, CLK=>
      nx10101, R=>RST);
   ix6829 : mux21_ni port map ( Y=>nx6828, A0=>Q_199_EXMPLR, A1=>D(199), S0
      =>nx10223);
   reg_Q_200 : dffr port map ( Q=>Q_200_EXMPLR, QB=>OPEN, D=>nx6838, CLK=>
      nx10101, R=>RST);
   ix6839 : mux21_ni port map ( Y=>nx6838, A0=>Q_200_EXMPLR, A1=>D(200), S0
      =>nx10223);
   reg_Q_201 : dffr port map ( Q=>Q_201_EXMPLR, QB=>OPEN, D=>nx6848, CLK=>
      nx10101, R=>RST);
   ix6849 : mux21_ni port map ( Y=>nx6848, A0=>Q_201_EXMPLR, A1=>D(201), S0
      =>nx10223);
   reg_Q_202 : dffr port map ( Q=>Q_202_EXMPLR, QB=>OPEN, D=>nx6858, CLK=>
      nx10101, R=>RST);
   ix6859 : mux21_ni port map ( Y=>nx6858, A0=>Q_202_EXMPLR, A1=>D(202), S0
      =>nx10223);
   reg_Q_203 : dffr port map ( Q=>Q_203_EXMPLR, QB=>OPEN, D=>nx6868, CLK=>
      nx10103, R=>RST);
   ix6869 : mux21_ni port map ( Y=>nx6868, A0=>Q_203_EXMPLR, A1=>D(203), S0
      =>nx10225);
   reg_Q_204 : dffr port map ( Q=>Q_204_EXMPLR, QB=>OPEN, D=>nx6878, CLK=>
      nx10103, R=>RST);
   ix6879 : mux21_ni port map ( Y=>nx6878, A0=>Q_204_EXMPLR, A1=>D(204), S0
      =>nx10225);
   reg_Q_205 : dffr port map ( Q=>Q_205_EXMPLR, QB=>OPEN, D=>nx6888, CLK=>
      nx10103, R=>RST);
   ix6889 : mux21_ni port map ( Y=>nx6888, A0=>Q_205_EXMPLR, A1=>D(205), S0
      =>nx10225);
   reg_Q_206 : dffr port map ( Q=>Q_206_EXMPLR, QB=>OPEN, D=>nx6898, CLK=>
      nx10103, R=>RST);
   ix6899 : mux21_ni port map ( Y=>nx6898, A0=>Q_206_EXMPLR, A1=>D(206), S0
      =>nx10225);
   reg_Q_207 : dffr port map ( Q=>Q_207_EXMPLR, QB=>OPEN, D=>nx6908, CLK=>
      nx10103, R=>RST);
   ix6909 : mux21_ni port map ( Y=>nx6908, A0=>Q_207_EXMPLR, A1=>D(207), S0
      =>nx10225);
   reg_Q_208 : dffr port map ( Q=>Q_208_EXMPLR, QB=>OPEN, D=>nx6918, CLK=>
      nx10103, R=>RST);
   ix6919 : mux21_ni port map ( Y=>nx6918, A0=>Q_208_EXMPLR, A1=>D(208), S0
      =>nx10225);
   reg_Q_209 : dffr port map ( Q=>Q_209_EXMPLR, QB=>OPEN, D=>nx6928, CLK=>
      nx10103, R=>RST);
   ix6929 : mux21_ni port map ( Y=>nx6928, A0=>Q_209_EXMPLR, A1=>D(209), S0
      =>nx10225);
   reg_Q_210 : dffr port map ( Q=>Q_210_EXMPLR, QB=>OPEN, D=>nx6938, CLK=>
      nx10105, R=>RST);
   ix6939 : mux21_ni port map ( Y=>nx6938, A0=>Q_210_EXMPLR, A1=>D(210), S0
      =>nx10227);
   reg_Q_211 : dffr port map ( Q=>Q_211_EXMPLR, QB=>OPEN, D=>nx6948, CLK=>
      nx10105, R=>RST);
   ix6949 : mux21_ni port map ( Y=>nx6948, A0=>Q_211_EXMPLR, A1=>D(211), S0
      =>nx10227);
   reg_Q_212 : dffr port map ( Q=>Q_212_EXMPLR, QB=>OPEN, D=>nx6958, CLK=>
      nx10105, R=>RST);
   ix6959 : mux21_ni port map ( Y=>nx6958, A0=>Q_212_EXMPLR, A1=>D(212), S0
      =>nx10227);
   reg_Q_213 : dffr port map ( Q=>Q_213_EXMPLR, QB=>OPEN, D=>nx6968, CLK=>
      nx10105, R=>RST);
   ix6969 : mux21_ni port map ( Y=>nx6968, A0=>Q_213_EXMPLR, A1=>D(213), S0
      =>nx10227);
   reg_Q_214 : dffr port map ( Q=>Q_214_EXMPLR, QB=>OPEN, D=>nx6978, CLK=>
      nx10105, R=>RST);
   ix6979 : mux21_ni port map ( Y=>nx6978, A0=>Q_214_EXMPLR, A1=>D(214), S0
      =>nx10227);
   reg_Q_215 : dffr port map ( Q=>Q_215_EXMPLR, QB=>OPEN, D=>nx6988, CLK=>
      nx10105, R=>RST);
   ix6989 : mux21_ni port map ( Y=>nx6988, A0=>Q_215_EXMPLR, A1=>D(215), S0
      =>nx10227);
   reg_Q_216 : dffr port map ( Q=>Q_216_EXMPLR, QB=>OPEN, D=>nx6998, CLK=>
      nx10105, R=>RST);
   ix6999 : mux21_ni port map ( Y=>nx6998, A0=>Q_216_EXMPLR, A1=>D(216), S0
      =>nx10227);
   reg_Q_217 : dffr port map ( Q=>Q_217_EXMPLR, QB=>OPEN, D=>nx7008, CLK=>
      nx10107, R=>RST);
   ix7009 : mux21_ni port map ( Y=>nx7008, A0=>Q_217_EXMPLR, A1=>D(217), S0
      =>nx10229);
   reg_Q_218 : dffr port map ( Q=>Q_218_EXMPLR, QB=>OPEN, D=>nx7018, CLK=>
      nx10107, R=>RST);
   ix7019 : mux21_ni port map ( Y=>nx7018, A0=>Q_218_EXMPLR, A1=>D(218), S0
      =>nx10229);
   reg_Q_219 : dffr port map ( Q=>Q_219_EXMPLR, QB=>OPEN, D=>nx7028, CLK=>
      nx10107, R=>RST);
   ix7029 : mux21_ni port map ( Y=>nx7028, A0=>Q_219_EXMPLR, A1=>D(219), S0
      =>nx10229);
   reg_Q_220 : dffr port map ( Q=>Q_220_EXMPLR, QB=>OPEN, D=>nx7038, CLK=>
      nx10107, R=>RST);
   ix7039 : mux21_ni port map ( Y=>nx7038, A0=>Q_220_EXMPLR, A1=>D(220), S0
      =>nx10229);
   reg_Q_221 : dffr port map ( Q=>Q_221_EXMPLR, QB=>OPEN, D=>nx7048, CLK=>
      nx10107, R=>RST);
   ix7049 : mux21_ni port map ( Y=>nx7048, A0=>Q_221_EXMPLR, A1=>D(221), S0
      =>nx10229);
   reg_Q_222 : dffr port map ( Q=>Q_222_EXMPLR, QB=>OPEN, D=>nx7058, CLK=>
      nx10107, R=>RST);
   ix7059 : mux21_ni port map ( Y=>nx7058, A0=>Q_222_EXMPLR, A1=>D(222), S0
      =>nx10229);
   reg_Q_223 : dffr port map ( Q=>Q_223_EXMPLR, QB=>OPEN, D=>nx7068, CLK=>
      nx10107, R=>RST);
   ix7069 : mux21_ni port map ( Y=>nx7068, A0=>Q_223_EXMPLR, A1=>D(223), S0
      =>nx10229);
   reg_Q_224 : dffr port map ( Q=>Q_224_EXMPLR, QB=>OPEN, D=>nx7078, CLK=>
      nx10109, R=>RST);
   ix7079 : mux21_ni port map ( Y=>nx7078, A0=>Q_224_EXMPLR, A1=>D(224), S0
      =>nx10231);
   reg_Q_225 : dffr port map ( Q=>Q_225_EXMPLR, QB=>OPEN, D=>nx7088, CLK=>
      nx10109, R=>RST);
   ix7089 : mux21_ni port map ( Y=>nx7088, A0=>Q_225_EXMPLR, A1=>D(225), S0
      =>nx10231);
   reg_Q_226 : dffr port map ( Q=>Q_226_EXMPLR, QB=>OPEN, D=>nx7098, CLK=>
      nx10109, R=>RST);
   ix7099 : mux21_ni port map ( Y=>nx7098, A0=>Q_226_EXMPLR, A1=>D(226), S0
      =>nx10231);
   reg_Q_227 : dffr port map ( Q=>Q_227_EXMPLR, QB=>OPEN, D=>nx7108, CLK=>
      nx10109, R=>RST);
   ix7109 : mux21_ni port map ( Y=>nx7108, A0=>Q_227_EXMPLR, A1=>D(227), S0
      =>nx10231);
   reg_Q_228 : dffr port map ( Q=>Q_228_EXMPLR, QB=>OPEN, D=>nx7118, CLK=>
      nx10109, R=>RST);
   ix7119 : mux21_ni port map ( Y=>nx7118, A0=>Q_228_EXMPLR, A1=>D(228), S0
      =>nx10231);
   reg_Q_229 : dffr port map ( Q=>Q_229_EXMPLR, QB=>OPEN, D=>nx7128, CLK=>
      nx10109, R=>RST);
   ix7129 : mux21_ni port map ( Y=>nx7128, A0=>Q_229_EXMPLR, A1=>D(229), S0
      =>nx10231);
   reg_Q_230 : dffr port map ( Q=>Q_230_EXMPLR, QB=>OPEN, D=>nx7138, CLK=>
      nx10109, R=>RST);
   ix7139 : mux21_ni port map ( Y=>nx7138, A0=>Q_230_EXMPLR, A1=>D(230), S0
      =>nx10231);
   reg_Q_231 : dffr port map ( Q=>Q_231_EXMPLR, QB=>OPEN, D=>nx7148, CLK=>
      nx10111, R=>RST);
   ix7149 : mux21_ni port map ( Y=>nx7148, A0=>Q_231_EXMPLR, A1=>D(231), S0
      =>nx10233);
   reg_Q_232 : dffr port map ( Q=>Q_232_EXMPLR, QB=>OPEN, D=>nx7158, CLK=>
      nx10111, R=>RST);
   ix7159 : mux21_ni port map ( Y=>nx7158, A0=>Q_232_EXMPLR, A1=>D(232), S0
      =>nx10233);
   reg_Q_233 : dffr port map ( Q=>Q_233_EXMPLR, QB=>OPEN, D=>nx7168, CLK=>
      nx10111, R=>RST);
   ix7169 : mux21_ni port map ( Y=>nx7168, A0=>Q_233_EXMPLR, A1=>D(233), S0
      =>nx10233);
   reg_Q_234 : dffr port map ( Q=>Q_234_EXMPLR, QB=>OPEN, D=>nx7178, CLK=>
      nx10111, R=>RST);
   ix7179 : mux21_ni port map ( Y=>nx7178, A0=>Q_234_EXMPLR, A1=>D(234), S0
      =>nx10233);
   reg_Q_235 : dffr port map ( Q=>Q_235_EXMPLR, QB=>OPEN, D=>nx7188, CLK=>
      nx10111, R=>RST);
   ix7189 : mux21_ni port map ( Y=>nx7188, A0=>Q_235_EXMPLR, A1=>D(235), S0
      =>nx10233);
   reg_Q_236 : dffr port map ( Q=>Q_236_EXMPLR, QB=>OPEN, D=>nx7198, CLK=>
      nx10111, R=>RST);
   ix7199 : mux21_ni port map ( Y=>nx7198, A0=>Q_236_EXMPLR, A1=>D(236), S0
      =>nx10233);
   reg_Q_237 : dffr port map ( Q=>Q_237_EXMPLR, QB=>OPEN, D=>nx7208, CLK=>
      nx10111, R=>RST);
   ix7209 : mux21_ni port map ( Y=>nx7208, A0=>Q_237_EXMPLR, A1=>D(237), S0
      =>nx10233);
   reg_Q_238 : dffr port map ( Q=>Q_238_EXMPLR, QB=>OPEN, D=>nx7218, CLK=>
      nx10113, R=>RST);
   ix7219 : mux21_ni port map ( Y=>nx7218, A0=>Q_238_EXMPLR, A1=>D(238), S0
      =>nx10235);
   reg_Q_239 : dffr port map ( Q=>Q_239_EXMPLR, QB=>OPEN, D=>nx7228, CLK=>
      nx10113, R=>RST);
   ix7229 : mux21_ni port map ( Y=>nx7228, A0=>Q_239_EXMPLR, A1=>D(239), S0
      =>nx10235);
   reg_Q_240 : dffr port map ( Q=>Q_240_EXMPLR, QB=>OPEN, D=>nx7238, CLK=>
      nx10113, R=>RST);
   ix7239 : mux21_ni port map ( Y=>nx7238, A0=>Q_240_EXMPLR, A1=>D(240), S0
      =>nx10235);
   reg_Q_241 : dffr port map ( Q=>Q_241_EXMPLR, QB=>OPEN, D=>nx7248, CLK=>
      nx10113, R=>RST);
   ix7249 : mux21_ni port map ( Y=>nx7248, A0=>Q_241_EXMPLR, A1=>D(241), S0
      =>nx10235);
   reg_Q_242 : dffr port map ( Q=>Q_242_EXMPLR, QB=>OPEN, D=>nx7258, CLK=>
      nx10113, R=>RST);
   ix7259 : mux21_ni port map ( Y=>nx7258, A0=>Q_242_EXMPLR, A1=>D(242), S0
      =>nx10235);
   reg_Q_243 : dffr port map ( Q=>Q_243_EXMPLR, QB=>OPEN, D=>nx7268, CLK=>
      nx10113, R=>RST);
   ix7269 : mux21_ni port map ( Y=>nx7268, A0=>Q_243_EXMPLR, A1=>D(243), S0
      =>nx10235);
   reg_Q_244 : dffr port map ( Q=>Q_244_EXMPLR, QB=>OPEN, D=>nx7278, CLK=>
      nx10113, R=>RST);
   ix7279 : mux21_ni port map ( Y=>nx7278, A0=>Q_244_EXMPLR, A1=>D(244), S0
      =>nx10235);
   reg_Q_245 : dffr port map ( Q=>Q_245_EXMPLR, QB=>OPEN, D=>nx7288, CLK=>
      nx10115, R=>RST);
   ix7289 : mux21_ni port map ( Y=>nx7288, A0=>Q_245_EXMPLR, A1=>D(245), S0
      =>nx10237);
   reg_Q_246 : dffr port map ( Q=>Q_246_EXMPLR, QB=>OPEN, D=>nx7298, CLK=>
      nx10115, R=>RST);
   ix7299 : mux21_ni port map ( Y=>nx7298, A0=>Q_246_EXMPLR, A1=>D(246), S0
      =>nx10237);
   reg_Q_247 : dffr port map ( Q=>Q_247_EXMPLR, QB=>OPEN, D=>nx7308, CLK=>
      nx10115, R=>RST);
   ix7309 : mux21_ni port map ( Y=>nx7308, A0=>Q_247_EXMPLR, A1=>D(247), S0
      =>nx10237);
   reg_Q_248 : dffr port map ( Q=>Q_248_EXMPLR, QB=>OPEN, D=>nx7318, CLK=>
      nx10115, R=>RST);
   ix7319 : mux21_ni port map ( Y=>nx7318, A0=>Q_248_EXMPLR, A1=>D(248), S0
      =>nx10237);
   reg_Q_249 : dffr port map ( Q=>Q_249_EXMPLR, QB=>OPEN, D=>nx7328, CLK=>
      nx10115, R=>RST);
   ix7329 : mux21_ni port map ( Y=>nx7328, A0=>Q_249_EXMPLR, A1=>D(249), S0
      =>nx10237);
   reg_Q_250 : dffr port map ( Q=>Q_250_EXMPLR, QB=>OPEN, D=>nx7338, CLK=>
      nx10115, R=>RST);
   ix7339 : mux21_ni port map ( Y=>nx7338, A0=>Q_250_EXMPLR, A1=>D(250), S0
      =>nx10237);
   reg_Q_251 : dffr port map ( Q=>Q_251_EXMPLR, QB=>OPEN, D=>nx7348, CLK=>
      nx10115, R=>RST);
   ix7349 : mux21_ni port map ( Y=>nx7348, A0=>Q_251_EXMPLR, A1=>D(251), S0
      =>nx10237);
   reg_Q_252 : dffr port map ( Q=>Q_252_EXMPLR, QB=>OPEN, D=>nx7358, CLK=>
      nx10117, R=>RST);
   ix7359 : mux21_ni port map ( Y=>nx7358, A0=>Q_252_EXMPLR, A1=>D(252), S0
      =>nx10239);
   reg_Q_253 : dffr port map ( Q=>Q_253_EXMPLR, QB=>OPEN, D=>nx7368, CLK=>
      nx10117, R=>RST);
   ix7369 : mux21_ni port map ( Y=>nx7368, A0=>Q_253_EXMPLR, A1=>D(253), S0
      =>nx10239);
   reg_Q_254 : dffr port map ( Q=>Q_254_EXMPLR, QB=>OPEN, D=>nx7378, CLK=>
      nx10117, R=>RST);
   ix7379 : mux21_ni port map ( Y=>nx7378, A0=>Q_254_EXMPLR, A1=>D(254), S0
      =>nx10239);
   reg_Q_255 : dffr port map ( Q=>Q_255_EXMPLR, QB=>OPEN, D=>nx7388, CLK=>
      nx10117, R=>RST);
   ix7389 : mux21_ni port map ( Y=>nx7388, A0=>Q_255_EXMPLR, A1=>D(255), S0
      =>nx10239);
   reg_Q_256 : dffr port map ( Q=>Q_256_EXMPLR, QB=>OPEN, D=>nx7398, CLK=>
      nx10117, R=>RST);
   ix7399 : mux21_ni port map ( Y=>nx7398, A0=>Q_256_EXMPLR, A1=>D(256), S0
      =>nx10239);
   reg_Q_257 : dffr port map ( Q=>Q_257_EXMPLR, QB=>OPEN, D=>nx7408, CLK=>
      nx10117, R=>RST);
   ix7409 : mux21_ni port map ( Y=>nx7408, A0=>Q_257_EXMPLR, A1=>D(257), S0
      =>nx10239);
   reg_Q_258 : dffr port map ( Q=>Q_258_EXMPLR, QB=>OPEN, D=>nx7418, CLK=>
      nx10117, R=>RST);
   ix7419 : mux21_ni port map ( Y=>nx7418, A0=>Q_258_EXMPLR, A1=>D(258), S0
      =>nx10239);
   reg_Q_259 : dffr port map ( Q=>Q_259_EXMPLR, QB=>OPEN, D=>nx7428, CLK=>
      nx10119, R=>RST);
   ix7429 : mux21_ni port map ( Y=>nx7428, A0=>Q_259_EXMPLR, A1=>D(259), S0
      =>nx10241);
   reg_Q_260 : dffr port map ( Q=>Q_260_EXMPLR, QB=>OPEN, D=>nx7438, CLK=>
      nx10119, R=>RST);
   ix7439 : mux21_ni port map ( Y=>nx7438, A0=>Q_260_EXMPLR, A1=>D(260), S0
      =>nx10241);
   reg_Q_261 : dffr port map ( Q=>Q_261_EXMPLR, QB=>OPEN, D=>nx7448, CLK=>
      nx10119, R=>RST);
   ix7449 : mux21_ni port map ( Y=>nx7448, A0=>Q_261_EXMPLR, A1=>D(261), S0
      =>nx10241);
   reg_Q_262 : dffr port map ( Q=>Q_262_EXMPLR, QB=>OPEN, D=>nx7458, CLK=>
      nx10119, R=>RST);
   ix7459 : mux21_ni port map ( Y=>nx7458, A0=>Q_262_EXMPLR, A1=>D(262), S0
      =>nx10241);
   reg_Q_263 : dffr port map ( Q=>Q_263_EXMPLR, QB=>OPEN, D=>nx7468, CLK=>
      nx10119, R=>RST);
   ix7469 : mux21_ni port map ( Y=>nx7468, A0=>Q_263_EXMPLR, A1=>D(263), S0
      =>nx10241);
   reg_Q_264 : dffr port map ( Q=>Q_264_EXMPLR, QB=>OPEN, D=>nx7478, CLK=>
      nx10119, R=>RST);
   ix7479 : mux21_ni port map ( Y=>nx7478, A0=>Q_264_EXMPLR, A1=>D(264), S0
      =>nx10241);
   reg_Q_265 : dffr port map ( Q=>Q_265_EXMPLR, QB=>OPEN, D=>nx7488, CLK=>
      nx10119, R=>RST);
   ix7489 : mux21_ni port map ( Y=>nx7488, A0=>Q_265_EXMPLR, A1=>D(265), S0
      =>nx10241);
   reg_Q_266 : dffr port map ( Q=>Q_266_EXMPLR, QB=>OPEN, D=>nx7498, CLK=>
      nx10121, R=>RST);
   ix7499 : mux21_ni port map ( Y=>nx7498, A0=>Q_266_EXMPLR, A1=>D(266), S0
      =>nx10243);
   reg_Q_267 : dffr port map ( Q=>Q_267_EXMPLR, QB=>OPEN, D=>nx7508, CLK=>
      nx10121, R=>RST);
   ix7509 : mux21_ni port map ( Y=>nx7508, A0=>Q_267_EXMPLR, A1=>D(267), S0
      =>nx10243);
   reg_Q_268 : dffr port map ( Q=>Q_268_EXMPLR, QB=>OPEN, D=>nx7518, CLK=>
      nx10121, R=>RST);
   ix7519 : mux21_ni port map ( Y=>nx7518, A0=>Q_268_EXMPLR, A1=>D(268), S0
      =>nx10243);
   reg_Q_269 : dffr port map ( Q=>Q_269_EXMPLR, QB=>OPEN, D=>nx7528, CLK=>
      nx10121, R=>RST);
   ix7529 : mux21_ni port map ( Y=>nx7528, A0=>Q_269_EXMPLR, A1=>D(269), S0
      =>nx10243);
   reg_Q_270 : dffr port map ( Q=>Q_270_EXMPLR, QB=>OPEN, D=>nx7538, CLK=>
      nx10121, R=>RST);
   ix7539 : mux21_ni port map ( Y=>nx7538, A0=>Q_270_EXMPLR, A1=>D(270), S0
      =>nx10243);
   reg_Q_271 : dffr port map ( Q=>Q_271_EXMPLR, QB=>OPEN, D=>nx7548, CLK=>
      nx10121, R=>RST);
   ix7549 : mux21_ni port map ( Y=>nx7548, A0=>Q_271_EXMPLR, A1=>D(271), S0
      =>nx10243);
   reg_Q_272 : dffr port map ( Q=>Q_272_EXMPLR, QB=>OPEN, D=>nx7558, CLK=>
      nx10121, R=>RST);
   ix7559 : mux21_ni port map ( Y=>nx7558, A0=>Q_272_EXMPLR, A1=>D(272), S0
      =>nx10243);
   reg_Q_273 : dffr port map ( Q=>Q_273_EXMPLR, QB=>OPEN, D=>nx7568, CLK=>
      nx10123, R=>RST);
   ix7569 : mux21_ni port map ( Y=>nx7568, A0=>Q_273_EXMPLR, A1=>D(273), S0
      =>nx10245);
   reg_Q_274 : dffr port map ( Q=>Q_274_EXMPLR, QB=>OPEN, D=>nx7578, CLK=>
      nx10123, R=>RST);
   ix7579 : mux21_ni port map ( Y=>nx7578, A0=>Q_274_EXMPLR, A1=>D(274), S0
      =>nx10245);
   reg_Q_275 : dffr port map ( Q=>Q_275_EXMPLR, QB=>OPEN, D=>nx7588, CLK=>
      nx10123, R=>RST);
   ix7589 : mux21_ni port map ( Y=>nx7588, A0=>Q_275_EXMPLR, A1=>D(275), S0
      =>nx10245);
   reg_Q_276 : dffr port map ( Q=>Q_276_EXMPLR, QB=>OPEN, D=>nx7598, CLK=>
      nx10123, R=>RST);
   ix7599 : mux21_ni port map ( Y=>nx7598, A0=>Q_276_EXMPLR, A1=>D(276), S0
      =>nx10245);
   reg_Q_277 : dffr port map ( Q=>Q_277_EXMPLR, QB=>OPEN, D=>nx7608, CLK=>
      nx10123, R=>RST);
   ix7609 : mux21_ni port map ( Y=>nx7608, A0=>Q_277_EXMPLR, A1=>D(277), S0
      =>nx10245);
   reg_Q_278 : dffr port map ( Q=>Q_278_EXMPLR, QB=>OPEN, D=>nx7618, CLK=>
      nx10123, R=>RST);
   ix7619 : mux21_ni port map ( Y=>nx7618, A0=>Q_278_EXMPLR, A1=>D(278), S0
      =>nx10245);
   reg_Q_279 : dffr port map ( Q=>Q_279_EXMPLR, QB=>OPEN, D=>nx7628, CLK=>
      nx10123, R=>RST);
   ix7629 : mux21_ni port map ( Y=>nx7628, A0=>Q_279_EXMPLR, A1=>D(279), S0
      =>nx10245);
   reg_Q_280 : dffr port map ( Q=>Q_280_EXMPLR, QB=>OPEN, D=>nx7638, CLK=>
      nx10125, R=>RST);
   ix7639 : mux21_ni port map ( Y=>nx7638, A0=>Q_280_EXMPLR, A1=>D(280), S0
      =>nx10247);
   reg_Q_281 : dffr port map ( Q=>Q_281_EXMPLR, QB=>OPEN, D=>nx7648, CLK=>
      nx10125, R=>RST);
   ix7649 : mux21_ni port map ( Y=>nx7648, A0=>Q_281_EXMPLR, A1=>D(281), S0
      =>nx10247);
   reg_Q_282 : dffr port map ( Q=>Q_282_EXMPLR, QB=>OPEN, D=>nx7658, CLK=>
      nx10125, R=>RST);
   ix7659 : mux21_ni port map ( Y=>nx7658, A0=>Q_282_EXMPLR, A1=>D(282), S0
      =>nx10247);
   reg_Q_283 : dffr port map ( Q=>Q_283_EXMPLR, QB=>OPEN, D=>nx7668, CLK=>
      nx10125, R=>RST);
   ix7669 : mux21_ni port map ( Y=>nx7668, A0=>Q_283_EXMPLR, A1=>D(283), S0
      =>nx10247);
   reg_Q_284 : dffr port map ( Q=>Q_284_EXMPLR, QB=>OPEN, D=>nx7678, CLK=>
      nx10125, R=>RST);
   ix7679 : mux21_ni port map ( Y=>nx7678, A0=>Q_284_EXMPLR, A1=>D(284), S0
      =>nx10247);
   reg_Q_285 : dffr port map ( Q=>Q_285_EXMPLR, QB=>OPEN, D=>nx7688, CLK=>
      nx10125, R=>RST);
   ix7689 : mux21_ni port map ( Y=>nx7688, A0=>Q_285_EXMPLR, A1=>D(285), S0
      =>nx10247);
   reg_Q_286 : dffr port map ( Q=>Q_286_EXMPLR, QB=>OPEN, D=>nx7698, CLK=>
      nx10125, R=>RST);
   ix7699 : mux21_ni port map ( Y=>nx7698, A0=>Q_286_EXMPLR, A1=>D(286), S0
      =>nx10247);
   reg_Q_287 : dffr port map ( Q=>Q_287_EXMPLR, QB=>OPEN, D=>nx7708, CLK=>
      nx10127, R=>RST);
   ix7709 : mux21_ni port map ( Y=>nx7708, A0=>Q_287_EXMPLR, A1=>D(287), S0
      =>nx10249);
   reg_Q_288 : dffr port map ( Q=>Q_288_EXMPLR, QB=>OPEN, D=>nx7718, CLK=>
      nx10127, R=>RST);
   ix7719 : mux21_ni port map ( Y=>nx7718, A0=>Q_288_EXMPLR, A1=>D(288), S0
      =>nx10249);
   reg_Q_289 : dffr port map ( Q=>Q_289_EXMPLR, QB=>OPEN, D=>nx7728, CLK=>
      nx10127, R=>RST);
   ix7729 : mux21_ni port map ( Y=>nx7728, A0=>Q_289_EXMPLR, A1=>D(289), S0
      =>nx10249);
   reg_Q_290 : dffr port map ( Q=>Q_290_EXMPLR, QB=>OPEN, D=>nx7738, CLK=>
      nx10127, R=>RST);
   ix7739 : mux21_ni port map ( Y=>nx7738, A0=>Q_290_EXMPLR, A1=>D(290), S0
      =>nx10249);
   reg_Q_291 : dffr port map ( Q=>Q_291_EXMPLR, QB=>OPEN, D=>nx7748, CLK=>
      nx10127, R=>RST);
   ix7749 : mux21_ni port map ( Y=>nx7748, A0=>Q_291_EXMPLR, A1=>D(291), S0
      =>nx10249);
   reg_Q_292 : dffr port map ( Q=>Q_292_EXMPLR, QB=>OPEN, D=>nx7758, CLK=>
      nx10127, R=>RST);
   ix7759 : mux21_ni port map ( Y=>nx7758, A0=>Q_292_EXMPLR, A1=>D(292), S0
      =>nx10249);
   reg_Q_293 : dffr port map ( Q=>Q_293_EXMPLR, QB=>OPEN, D=>nx7768, CLK=>
      nx10127, R=>RST);
   ix7769 : mux21_ni port map ( Y=>nx7768, A0=>Q_293_EXMPLR, A1=>D(293), S0
      =>nx10249);
   reg_Q_294 : dffr port map ( Q=>Q_294_EXMPLR, QB=>OPEN, D=>nx7778, CLK=>
      nx10129, R=>RST);
   ix7779 : mux21_ni port map ( Y=>nx7778, A0=>Q_294_EXMPLR, A1=>D(294), S0
      =>nx10251);
   reg_Q_295 : dffr port map ( Q=>Q_295_EXMPLR, QB=>OPEN, D=>nx7788, CLK=>
      nx10129, R=>RST);
   ix7789 : mux21_ni port map ( Y=>nx7788, A0=>Q_295_EXMPLR, A1=>D(295), S0
      =>nx10251);
   reg_Q_296 : dffr port map ( Q=>Q_296_EXMPLR, QB=>OPEN, D=>nx7798, CLK=>
      nx10129, R=>RST);
   ix7799 : mux21_ni port map ( Y=>nx7798, A0=>Q_296_EXMPLR, A1=>D(296), S0
      =>nx10251);
   reg_Q_297 : dffr port map ( Q=>Q_297_EXMPLR, QB=>OPEN, D=>nx7808, CLK=>
      nx10129, R=>RST);
   ix7809 : mux21_ni port map ( Y=>nx7808, A0=>Q_297_EXMPLR, A1=>D(297), S0
      =>nx10251);
   reg_Q_298 : dffr port map ( Q=>Q_298_EXMPLR, QB=>OPEN, D=>nx7818, CLK=>
      nx10129, R=>RST);
   ix7819 : mux21_ni port map ( Y=>nx7818, A0=>Q_298_EXMPLR, A1=>D(298), S0
      =>nx10251);
   reg_Q_299 : dffr port map ( Q=>Q_299_EXMPLR, QB=>OPEN, D=>nx7828, CLK=>
      nx10129, R=>RST);
   ix7829 : mux21_ni port map ( Y=>nx7828, A0=>Q_299_EXMPLR, A1=>D(299), S0
      =>nx10251);
   reg_Q_300 : dffr port map ( Q=>Q_300_EXMPLR, QB=>OPEN, D=>nx7838, CLK=>
      nx10129, R=>RST);
   ix7839 : mux21_ni port map ( Y=>nx7838, A0=>Q_300_EXMPLR, A1=>D(300), S0
      =>nx10251);
   reg_Q_301 : dffr port map ( Q=>Q_301_EXMPLR, QB=>OPEN, D=>nx7848, CLK=>
      nx10131, R=>RST);
   ix7849 : mux21_ni port map ( Y=>nx7848, A0=>Q_301_EXMPLR, A1=>D(301), S0
      =>nx10253);
   reg_Q_302 : dffr port map ( Q=>Q_302_EXMPLR, QB=>OPEN, D=>nx7858, CLK=>
      nx10131, R=>RST);
   ix7859 : mux21_ni port map ( Y=>nx7858, A0=>Q_302_EXMPLR, A1=>D(302), S0
      =>nx10253);
   reg_Q_303 : dffr port map ( Q=>Q_303_EXMPLR, QB=>OPEN, D=>nx7868, CLK=>
      nx10131, R=>RST);
   ix7869 : mux21_ni port map ( Y=>nx7868, A0=>Q_303_EXMPLR, A1=>D(303), S0
      =>nx10253);
   reg_Q_304 : dffr port map ( Q=>Q_304_EXMPLR, QB=>OPEN, D=>nx7878, CLK=>
      nx10131, R=>RST);
   ix7879 : mux21_ni port map ( Y=>nx7878, A0=>Q_304_EXMPLR, A1=>D(304), S0
      =>nx10253);
   reg_Q_305 : dffr port map ( Q=>Q_305_EXMPLR, QB=>OPEN, D=>nx7888, CLK=>
      nx10131, R=>RST);
   ix7889 : mux21_ni port map ( Y=>nx7888, A0=>Q_305_EXMPLR, A1=>D(305), S0
      =>nx10253);
   reg_Q_306 : dffr port map ( Q=>Q_306_EXMPLR, QB=>OPEN, D=>nx7898, CLK=>
      nx10131, R=>RST);
   ix7899 : mux21_ni port map ( Y=>nx7898, A0=>Q_306_EXMPLR, A1=>D(306), S0
      =>nx10253);
   reg_Q_307 : dffr port map ( Q=>Q_307_EXMPLR, QB=>OPEN, D=>nx7908, CLK=>
      nx10131, R=>RST);
   ix7909 : mux21_ni port map ( Y=>nx7908, A0=>Q_307_EXMPLR, A1=>D(307), S0
      =>nx10253);
   reg_Q_308 : dffr port map ( Q=>Q_308_EXMPLR, QB=>OPEN, D=>nx7918, CLK=>
      nx10133, R=>RST);
   ix7919 : mux21_ni port map ( Y=>nx7918, A0=>Q_308_EXMPLR, A1=>D(308), S0
      =>nx10255);
   reg_Q_309 : dffr port map ( Q=>Q_309_EXMPLR, QB=>OPEN, D=>nx7928, CLK=>
      nx10133, R=>RST);
   ix7929 : mux21_ni port map ( Y=>nx7928, A0=>Q_309_EXMPLR, A1=>D(309), S0
      =>nx10255);
   reg_Q_310 : dffr port map ( Q=>Q_310_EXMPLR, QB=>OPEN, D=>nx7938, CLK=>
      nx10133, R=>RST);
   ix7939 : mux21_ni port map ( Y=>nx7938, A0=>Q_310_EXMPLR, A1=>D(310), S0
      =>nx10255);
   reg_Q_311 : dffr port map ( Q=>Q_311_EXMPLR, QB=>OPEN, D=>nx7948, CLK=>
      nx10133, R=>RST);
   ix7949 : mux21_ni port map ( Y=>nx7948, A0=>Q_311_EXMPLR, A1=>D(311), S0
      =>nx10255);
   reg_Q_312 : dffr port map ( Q=>Q_312_EXMPLR, QB=>OPEN, D=>nx7958, CLK=>
      nx10133, R=>RST);
   ix7959 : mux21_ni port map ( Y=>nx7958, A0=>Q_312_EXMPLR, A1=>D(312), S0
      =>nx10255);
   reg_Q_313 : dffr port map ( Q=>Q_313_EXMPLR, QB=>OPEN, D=>nx7968, CLK=>
      nx10133, R=>RST);
   ix7969 : mux21_ni port map ( Y=>nx7968, A0=>Q_313_EXMPLR, A1=>D(313), S0
      =>nx10255);
   reg_Q_314 : dffr port map ( Q=>Q_314_EXMPLR, QB=>OPEN, D=>nx7978, CLK=>
      nx10133, R=>RST);
   ix7979 : mux21_ni port map ( Y=>nx7978, A0=>Q_314_EXMPLR, A1=>D(314), S0
      =>nx10255);
   reg_Q_315 : dffr port map ( Q=>Q_315_EXMPLR, QB=>OPEN, D=>nx7988, CLK=>
      nx10135, R=>RST);
   ix7989 : mux21_ni port map ( Y=>nx7988, A0=>Q_315_EXMPLR, A1=>D(315), S0
      =>nx10257);
   reg_Q_316 : dffr port map ( Q=>Q_316_EXMPLR, QB=>OPEN, D=>nx7998, CLK=>
      nx10135, R=>RST);
   ix7999 : mux21_ni port map ( Y=>nx7998, A0=>Q_316_EXMPLR, A1=>D(316), S0
      =>nx10257);
   reg_Q_317 : dffr port map ( Q=>Q_317_EXMPLR, QB=>OPEN, D=>nx8008, CLK=>
      nx10135, R=>RST);
   ix8009 : mux21_ni port map ( Y=>nx8008, A0=>Q_317_EXMPLR, A1=>D(317), S0
      =>nx10257);
   reg_Q_318 : dffr port map ( Q=>Q_318_EXMPLR, QB=>OPEN, D=>nx8018, CLK=>
      nx10135, R=>RST);
   ix8019 : mux21_ni port map ( Y=>nx8018, A0=>Q_318_EXMPLR, A1=>D(318), S0
      =>nx10257);
   reg_Q_319 : dffr port map ( Q=>Q_319_EXMPLR, QB=>OPEN, D=>nx8028, CLK=>
      nx10135, R=>RST);
   ix8029 : mux21_ni port map ( Y=>nx8028, A0=>Q_319_EXMPLR, A1=>D(319), S0
      =>nx10257);
   reg_Q_320 : dffr port map ( Q=>Q_320_EXMPLR, QB=>OPEN, D=>nx8038, CLK=>
      nx10135, R=>RST);
   ix8039 : mux21_ni port map ( Y=>nx8038, A0=>Q_320_EXMPLR, A1=>D(320), S0
      =>nx10257);
   reg_Q_321 : dffr port map ( Q=>Q_321_EXMPLR, QB=>OPEN, D=>nx8048, CLK=>
      nx10135, R=>RST);
   ix8049 : mux21_ni port map ( Y=>nx8048, A0=>Q_321_EXMPLR, A1=>D(321), S0
      =>nx10257);
   reg_Q_322 : dffr port map ( Q=>Q_322_EXMPLR, QB=>OPEN, D=>nx8058, CLK=>
      nx10137, R=>RST);
   ix8059 : mux21_ni port map ( Y=>nx8058, A0=>Q_322_EXMPLR, A1=>D(322), S0
      =>nx10259);
   reg_Q_323 : dffr port map ( Q=>Q_323_EXMPLR, QB=>OPEN, D=>nx8068, CLK=>
      nx10137, R=>RST);
   ix8069 : mux21_ni port map ( Y=>nx8068, A0=>Q_323_EXMPLR, A1=>D(323), S0
      =>nx10259);
   reg_Q_324 : dffr port map ( Q=>Q_324_EXMPLR, QB=>OPEN, D=>nx8078, CLK=>
      nx10137, R=>RST);
   ix8079 : mux21_ni port map ( Y=>nx8078, A0=>Q_324_EXMPLR, A1=>D(324), S0
      =>nx10259);
   reg_Q_325 : dffr port map ( Q=>Q_325_EXMPLR, QB=>OPEN, D=>nx8088, CLK=>
      nx10137, R=>RST);
   ix8089 : mux21_ni port map ( Y=>nx8088, A0=>Q_325_EXMPLR, A1=>D(325), S0
      =>nx10259);
   reg_Q_326 : dffr port map ( Q=>Q_326_EXMPLR, QB=>OPEN, D=>nx8098, CLK=>
      nx10137, R=>RST);
   ix8099 : mux21_ni port map ( Y=>nx8098, A0=>Q_326_EXMPLR, A1=>D(326), S0
      =>nx10259);
   reg_Q_327 : dffr port map ( Q=>Q_327_EXMPLR, QB=>OPEN, D=>nx8108, CLK=>
      nx10137, R=>RST);
   ix8109 : mux21_ni port map ( Y=>nx8108, A0=>Q_327_EXMPLR, A1=>D(327), S0
      =>nx10259);
   reg_Q_328 : dffr port map ( Q=>Q_328_EXMPLR, QB=>OPEN, D=>nx8118, CLK=>
      nx10137, R=>RST);
   ix8119 : mux21_ni port map ( Y=>nx8118, A0=>Q_328_EXMPLR, A1=>D(328), S0
      =>nx10259);
   reg_Q_329 : dffr port map ( Q=>Q_329_EXMPLR, QB=>OPEN, D=>nx8128, CLK=>
      nx10139, R=>RST);
   ix8129 : mux21_ni port map ( Y=>nx8128, A0=>Q_329_EXMPLR, A1=>D(329), S0
      =>nx10261);
   reg_Q_330 : dffr port map ( Q=>Q_330_EXMPLR, QB=>OPEN, D=>nx8138, CLK=>
      nx10139, R=>RST);
   ix8139 : mux21_ni port map ( Y=>nx8138, A0=>Q_330_EXMPLR, A1=>D(330), S0
      =>nx10261);
   reg_Q_331 : dffr port map ( Q=>Q_331_EXMPLR, QB=>OPEN, D=>nx8148, CLK=>
      nx10139, R=>RST);
   ix8149 : mux21_ni port map ( Y=>nx8148, A0=>Q_331_EXMPLR, A1=>D(331), S0
      =>nx10261);
   reg_Q_332 : dffr port map ( Q=>Q_332_EXMPLR, QB=>OPEN, D=>nx8158, CLK=>
      nx10139, R=>RST);
   ix8159 : mux21_ni port map ( Y=>nx8158, A0=>Q_332_EXMPLR, A1=>D(332), S0
      =>nx10261);
   reg_Q_333 : dffr port map ( Q=>Q_333_EXMPLR, QB=>OPEN, D=>nx8168, CLK=>
      nx10139, R=>RST);
   ix8169 : mux21_ni port map ( Y=>nx8168, A0=>Q_333_EXMPLR, A1=>D(333), S0
      =>nx10261);
   reg_Q_334 : dffr port map ( Q=>Q_334_EXMPLR, QB=>OPEN, D=>nx8178, CLK=>
      nx10139, R=>RST);
   ix8179 : mux21_ni port map ( Y=>nx8178, A0=>Q_334_EXMPLR, A1=>D(334), S0
      =>nx10261);
   reg_Q_335 : dffr port map ( Q=>Q_335_EXMPLR, QB=>OPEN, D=>nx8188, CLK=>
      nx10139, R=>RST);
   ix8189 : mux21_ni port map ( Y=>nx8188, A0=>Q_335_EXMPLR, A1=>D(335), S0
      =>nx10261);
   reg_Q_336 : dffr port map ( Q=>Q_336_EXMPLR, QB=>OPEN, D=>nx8198, CLK=>
      nx10141, R=>RST);
   ix8199 : mux21_ni port map ( Y=>nx8198, A0=>Q_336_EXMPLR, A1=>D(336), S0
      =>nx10263);
   reg_Q_337 : dffr port map ( Q=>Q_337_EXMPLR, QB=>OPEN, D=>nx8208, CLK=>
      nx10141, R=>RST);
   ix8209 : mux21_ni port map ( Y=>nx8208, A0=>Q_337_EXMPLR, A1=>D(337), S0
      =>nx10263);
   reg_Q_338 : dffr port map ( Q=>Q_338_EXMPLR, QB=>OPEN, D=>nx8218, CLK=>
      nx10141, R=>RST);
   ix8219 : mux21_ni port map ( Y=>nx8218, A0=>Q_338_EXMPLR, A1=>D(338), S0
      =>nx10263);
   reg_Q_339 : dffr port map ( Q=>Q_339_EXMPLR, QB=>OPEN, D=>nx8228, CLK=>
      nx10141, R=>RST);
   ix8229 : mux21_ni port map ( Y=>nx8228, A0=>Q_339_EXMPLR, A1=>D(339), S0
      =>nx10263);
   reg_Q_340 : dffr port map ( Q=>Q_340_EXMPLR, QB=>OPEN, D=>nx8238, CLK=>
      nx10141, R=>RST);
   ix8239 : mux21_ni port map ( Y=>nx8238, A0=>Q_340_EXMPLR, A1=>D(340), S0
      =>nx10263);
   reg_Q_341 : dffr port map ( Q=>Q_341_EXMPLR, QB=>OPEN, D=>nx8248, CLK=>
      nx10141, R=>RST);
   ix8249 : mux21_ni port map ( Y=>nx8248, A0=>Q_341_EXMPLR, A1=>D(341), S0
      =>nx10263);
   reg_Q_342 : dffr port map ( Q=>Q_342_EXMPLR, QB=>OPEN, D=>nx8258, CLK=>
      nx10141, R=>RST);
   ix8259 : mux21_ni port map ( Y=>nx8258, A0=>Q_342_EXMPLR, A1=>D(342), S0
      =>nx10263);
   reg_Q_343 : dffr port map ( Q=>Q_343_EXMPLR, QB=>OPEN, D=>nx8268, CLK=>
      nx10143, R=>RST);
   ix8269 : mux21_ni port map ( Y=>nx8268, A0=>Q_343_EXMPLR, A1=>D(343), S0
      =>nx10265);
   reg_Q_344 : dffr port map ( Q=>Q_344_EXMPLR, QB=>OPEN, D=>nx8278, CLK=>
      nx10143, R=>RST);
   ix8279 : mux21_ni port map ( Y=>nx8278, A0=>Q_344_EXMPLR, A1=>D(344), S0
      =>nx10265);
   reg_Q_345 : dffr port map ( Q=>Q_345_EXMPLR, QB=>OPEN, D=>nx8288, CLK=>
      nx10143, R=>RST);
   ix8289 : mux21_ni port map ( Y=>nx8288, A0=>Q_345_EXMPLR, A1=>D(345), S0
      =>nx10265);
   reg_Q_346 : dffr port map ( Q=>Q_346_EXMPLR, QB=>OPEN, D=>nx8298, CLK=>
      nx10143, R=>RST);
   ix8299 : mux21_ni port map ( Y=>nx8298, A0=>Q_346_EXMPLR, A1=>D(346), S0
      =>nx10265);
   reg_Q_347 : dffr port map ( Q=>Q_347_EXMPLR, QB=>OPEN, D=>nx8308, CLK=>
      nx10143, R=>RST);
   ix8309 : mux21_ni port map ( Y=>nx8308, A0=>Q_347_EXMPLR, A1=>D(347), S0
      =>nx10265);
   reg_Q_348 : dffr port map ( Q=>Q_348_EXMPLR, QB=>OPEN, D=>nx8318, CLK=>
      nx10143, R=>RST);
   ix8319 : mux21_ni port map ( Y=>nx8318, A0=>Q_348_EXMPLR, A1=>D(348), S0
      =>nx10265);
   reg_Q_349 : dffr port map ( Q=>Q_349_EXMPLR, QB=>OPEN, D=>nx8328, CLK=>
      nx10143, R=>RST);
   ix8329 : mux21_ni port map ( Y=>nx8328, A0=>Q_349_EXMPLR, A1=>D(349), S0
      =>nx10265);
   reg_Q_350 : dffr port map ( Q=>Q_350_EXMPLR, QB=>OPEN, D=>nx8338, CLK=>
      nx10145, R=>RST);
   ix8339 : mux21_ni port map ( Y=>nx8338, A0=>Q_350_EXMPLR, A1=>D(350), S0
      =>nx10267);
   reg_Q_351 : dffr port map ( Q=>Q_351_EXMPLR, QB=>OPEN, D=>nx8348, CLK=>
      nx10145, R=>RST);
   ix8349 : mux21_ni port map ( Y=>nx8348, A0=>Q_351_EXMPLR, A1=>D(351), S0
      =>nx10267);
   reg_Q_352 : dffr port map ( Q=>Q_352_EXMPLR, QB=>OPEN, D=>nx8358, CLK=>
      nx10145, R=>RST);
   ix8359 : mux21_ni port map ( Y=>nx8358, A0=>Q_352_EXMPLR, A1=>D(352), S0
      =>nx10267);
   reg_Q_353 : dffr port map ( Q=>Q_353_EXMPLR, QB=>OPEN, D=>nx8368, CLK=>
      nx10145, R=>RST);
   ix8369 : mux21_ni port map ( Y=>nx8368, A0=>Q_353_EXMPLR, A1=>D(353), S0
      =>nx10267);
   reg_Q_354 : dffr port map ( Q=>Q_354_EXMPLR, QB=>OPEN, D=>nx8378, CLK=>
      nx10145, R=>RST);
   ix8379 : mux21_ni port map ( Y=>nx8378, A0=>Q_354_EXMPLR, A1=>D(354), S0
      =>nx10267);
   reg_Q_355 : dffr port map ( Q=>Q_355_EXMPLR, QB=>OPEN, D=>nx8388, CLK=>
      nx10145, R=>RST);
   ix8389 : mux21_ni port map ( Y=>nx8388, A0=>Q_355_EXMPLR, A1=>D(355), S0
      =>nx10267);
   reg_Q_356 : dffr port map ( Q=>Q_356_EXMPLR, QB=>OPEN, D=>nx8398, CLK=>
      nx10145, R=>RST);
   ix8399 : mux21_ni port map ( Y=>nx8398, A0=>Q_356_EXMPLR, A1=>D(356), S0
      =>nx10267);
   reg_Q_357 : dffr port map ( Q=>Q_357_EXMPLR, QB=>OPEN, D=>nx8408, CLK=>
      nx10147, R=>RST);
   ix8409 : mux21_ni port map ( Y=>nx8408, A0=>Q_357_EXMPLR, A1=>D(357), S0
      =>nx10269);
   reg_Q_358 : dffr port map ( Q=>Q_358_EXMPLR, QB=>OPEN, D=>nx8418, CLK=>
      nx10147, R=>RST);
   ix8419 : mux21_ni port map ( Y=>nx8418, A0=>Q_358_EXMPLR, A1=>D(358), S0
      =>nx10269);
   reg_Q_359 : dffr port map ( Q=>Q_359_EXMPLR, QB=>OPEN, D=>nx8428, CLK=>
      nx10147, R=>RST);
   ix8429 : mux21_ni port map ( Y=>nx8428, A0=>Q_359_EXMPLR, A1=>D(359), S0
      =>nx10269);
   reg_Q_360 : dffr port map ( Q=>Q_360_EXMPLR, QB=>OPEN, D=>nx8438, CLK=>
      nx10147, R=>RST);
   ix8439 : mux21_ni port map ( Y=>nx8438, A0=>Q_360_EXMPLR, A1=>D(360), S0
      =>nx10269);
   reg_Q_361 : dffr port map ( Q=>Q_361_EXMPLR, QB=>OPEN, D=>nx8448, CLK=>
      nx10147, R=>RST);
   ix8449 : mux21_ni port map ( Y=>nx8448, A0=>Q_361_EXMPLR, A1=>D(361), S0
      =>nx10269);
   reg_Q_362 : dffr port map ( Q=>Q_362_EXMPLR, QB=>OPEN, D=>nx8458, CLK=>
      nx10147, R=>RST);
   ix8459 : mux21_ni port map ( Y=>nx8458, A0=>Q_362_EXMPLR, A1=>D(362), S0
      =>nx10269);
   reg_Q_363 : dffr port map ( Q=>Q_363_EXMPLR, QB=>OPEN, D=>nx8468, CLK=>
      nx10147, R=>RST);
   ix8469 : mux21_ni port map ( Y=>nx8468, A0=>Q_363_EXMPLR, A1=>D(363), S0
      =>nx10269);
   reg_Q_364 : dffr port map ( Q=>Q_364_EXMPLR, QB=>OPEN, D=>nx8478, CLK=>
      nx10149, R=>RST);
   ix8479 : mux21_ni port map ( Y=>nx8478, A0=>Q_364_EXMPLR, A1=>D(364), S0
      =>nx10271);
   reg_Q_365 : dffr port map ( Q=>Q_365_EXMPLR, QB=>OPEN, D=>nx8488, CLK=>
      nx10149, R=>RST);
   ix8489 : mux21_ni port map ( Y=>nx8488, A0=>Q_365_EXMPLR, A1=>D(365), S0
      =>nx10271);
   reg_Q_366 : dffr port map ( Q=>Q_366_EXMPLR, QB=>OPEN, D=>nx8498, CLK=>
      nx10149, R=>RST);
   ix8499 : mux21_ni port map ( Y=>nx8498, A0=>Q_366_EXMPLR, A1=>D(366), S0
      =>nx10271);
   reg_Q_367 : dffr port map ( Q=>Q_367_EXMPLR, QB=>OPEN, D=>nx8508, CLK=>
      nx10149, R=>RST);
   ix8509 : mux21_ni port map ( Y=>nx8508, A0=>Q_367_EXMPLR, A1=>D(367), S0
      =>nx10271);
   reg_Q_368 : dffr port map ( Q=>Q_368_EXMPLR, QB=>OPEN, D=>nx8518, CLK=>
      nx10149, R=>RST);
   ix8519 : mux21_ni port map ( Y=>nx8518, A0=>Q_368_EXMPLR, A1=>D(368), S0
      =>nx10271);
   reg_Q_369 : dffr port map ( Q=>Q_369_EXMPLR, QB=>OPEN, D=>nx8528, CLK=>
      nx10149, R=>RST);
   ix8529 : mux21_ni port map ( Y=>nx8528, A0=>Q_369_EXMPLR, A1=>D(369), S0
      =>nx10271);
   reg_Q_370 : dffr port map ( Q=>Q_370_EXMPLR, QB=>OPEN, D=>nx8538, CLK=>
      nx10149, R=>RST);
   ix8539 : mux21_ni port map ( Y=>nx8538, A0=>Q_370_EXMPLR, A1=>D(370), S0
      =>nx10271);
   reg_Q_371 : dffr port map ( Q=>Q_371_EXMPLR, QB=>OPEN, D=>nx8548, CLK=>
      nx10151, R=>RST);
   ix8549 : mux21_ni port map ( Y=>nx8548, A0=>Q_371_EXMPLR, A1=>D(371), S0
      =>nx10273);
   reg_Q_372 : dffr port map ( Q=>Q_372_EXMPLR, QB=>OPEN, D=>nx8558, CLK=>
      nx10151, R=>RST);
   ix8559 : mux21_ni port map ( Y=>nx8558, A0=>Q_372_EXMPLR, A1=>D(372), S0
      =>nx10273);
   reg_Q_373 : dffr port map ( Q=>Q_373_EXMPLR, QB=>OPEN, D=>nx8568, CLK=>
      nx10151, R=>RST);
   ix8569 : mux21_ni port map ( Y=>nx8568, A0=>Q_373_EXMPLR, A1=>D(373), S0
      =>nx10273);
   reg_Q_374 : dffr port map ( Q=>Q_374_EXMPLR, QB=>OPEN, D=>nx8578, CLK=>
      nx10151, R=>RST);
   ix8579 : mux21_ni port map ( Y=>nx8578, A0=>Q_374_EXMPLR, A1=>D(374), S0
      =>nx10273);
   reg_Q_375 : dffr port map ( Q=>Q_375_EXMPLR, QB=>OPEN, D=>nx8588, CLK=>
      nx10151, R=>RST);
   ix8589 : mux21_ni port map ( Y=>nx8588, A0=>Q_375_EXMPLR, A1=>D(375), S0
      =>nx10273);
   reg_Q_376 : dffr port map ( Q=>Q_376_EXMPLR, QB=>OPEN, D=>nx8598, CLK=>
      nx10151, R=>RST);
   ix8599 : mux21_ni port map ( Y=>nx8598, A0=>Q_376_EXMPLR, A1=>D(376), S0
      =>nx10273);
   reg_Q_377 : dffr port map ( Q=>Q_377_EXMPLR, QB=>OPEN, D=>nx8608, CLK=>
      nx10151, R=>RST);
   ix8609 : mux21_ni port map ( Y=>nx8608, A0=>Q_377_EXMPLR, A1=>D(377), S0
      =>nx10273);
   reg_Q_378 : dffr port map ( Q=>Q_378_EXMPLR, QB=>OPEN, D=>nx8618, CLK=>
      nx10153, R=>RST);
   ix8619 : mux21_ni port map ( Y=>nx8618, A0=>Q_378_EXMPLR, A1=>D(378), S0
      =>nx10275);
   reg_Q_379 : dffr port map ( Q=>Q_379_EXMPLR, QB=>OPEN, D=>nx8628, CLK=>
      nx10153, R=>RST);
   ix8629 : mux21_ni port map ( Y=>nx8628, A0=>Q_379_EXMPLR, A1=>D(379), S0
      =>nx10275);
   reg_Q_380 : dffr port map ( Q=>Q_380_EXMPLR, QB=>OPEN, D=>nx8638, CLK=>
      nx10153, R=>RST);
   ix8639 : mux21_ni port map ( Y=>nx8638, A0=>Q_380_EXMPLR, A1=>D(380), S0
      =>nx10275);
   reg_Q_381 : dffr port map ( Q=>Q_381_EXMPLR, QB=>OPEN, D=>nx8648, CLK=>
      nx10153, R=>RST);
   ix8649 : mux21_ni port map ( Y=>nx8648, A0=>Q_381_EXMPLR, A1=>D(381), S0
      =>nx10275);
   reg_Q_382 : dffr port map ( Q=>Q_382_EXMPLR, QB=>OPEN, D=>nx8658, CLK=>
      nx10153, R=>RST);
   ix8659 : mux21_ni port map ( Y=>nx8658, A0=>Q_382_EXMPLR, A1=>D(382), S0
      =>nx10275);
   reg_Q_383 : dffr port map ( Q=>Q_383_EXMPLR, QB=>OPEN, D=>nx8668, CLK=>
      nx10153, R=>RST);
   ix8669 : mux21_ni port map ( Y=>nx8668, A0=>Q_383_EXMPLR, A1=>D(383), S0
      =>nx10275);
   reg_Q_384 : dffr port map ( Q=>Q_384_EXMPLR, QB=>OPEN, D=>nx8678, CLK=>
      nx10153, R=>RST);
   ix8679 : mux21_ni port map ( Y=>nx8678, A0=>Q_384_EXMPLR, A1=>D(384), S0
      =>nx10275);
   reg_Q_385 : dffr port map ( Q=>Q_385_EXMPLR, QB=>OPEN, D=>nx8688, CLK=>
      nx10155, R=>RST);
   ix8689 : mux21_ni port map ( Y=>nx8688, A0=>Q_385_EXMPLR, A1=>D(385), S0
      =>nx10277);
   reg_Q_386 : dffr port map ( Q=>Q_386_EXMPLR, QB=>OPEN, D=>nx8698, CLK=>
      nx10155, R=>RST);
   ix8699 : mux21_ni port map ( Y=>nx8698, A0=>Q_386_EXMPLR, A1=>D(386), S0
      =>nx10277);
   reg_Q_387 : dffr port map ( Q=>Q_387_EXMPLR, QB=>OPEN, D=>nx8708, CLK=>
      nx10155, R=>RST);
   ix8709 : mux21_ni port map ( Y=>nx8708, A0=>Q_387_EXMPLR, A1=>D(387), S0
      =>nx10277);
   reg_Q_388 : dffr port map ( Q=>Q_388_EXMPLR, QB=>OPEN, D=>nx8718, CLK=>
      nx10155, R=>RST);
   ix8719 : mux21_ni port map ( Y=>nx8718, A0=>Q_388_EXMPLR, A1=>D(388), S0
      =>nx10277);
   reg_Q_389 : dffr port map ( Q=>Q_389_EXMPLR, QB=>OPEN, D=>nx8728, CLK=>
      nx10155, R=>RST);
   ix8729 : mux21_ni port map ( Y=>nx8728, A0=>Q_389_EXMPLR, A1=>D(389), S0
      =>nx10277);
   reg_Q_390 : dffr port map ( Q=>Q_390_EXMPLR, QB=>OPEN, D=>nx8738, CLK=>
      nx10155, R=>RST);
   ix8739 : mux21_ni port map ( Y=>nx8738, A0=>Q_390_EXMPLR, A1=>D(390), S0
      =>nx10277);
   reg_Q_391 : dffr port map ( Q=>Q_391_EXMPLR, QB=>OPEN, D=>nx8748, CLK=>
      nx10155, R=>RST);
   ix8749 : mux21_ni port map ( Y=>nx8748, A0=>Q_391_EXMPLR, A1=>D(391), S0
      =>nx10277);
   reg_Q_392 : dffr port map ( Q=>Q_392_EXMPLR, QB=>OPEN, D=>nx8758, CLK=>
      nx10157, R=>RST);
   ix8759 : mux21_ni port map ( Y=>nx8758, A0=>Q_392_EXMPLR, A1=>D(392), S0
      =>nx10279);
   reg_Q_393 : dffr port map ( Q=>Q_393_EXMPLR, QB=>OPEN, D=>nx8768, CLK=>
      nx10157, R=>RST);
   ix8769 : mux21_ni port map ( Y=>nx8768, A0=>Q_393_EXMPLR, A1=>D(393), S0
      =>nx10279);
   reg_Q_394 : dffr port map ( Q=>Q_394_EXMPLR, QB=>OPEN, D=>nx8778, CLK=>
      nx10157, R=>RST);
   ix8779 : mux21_ni port map ( Y=>nx8778, A0=>Q_394_EXMPLR, A1=>D(394), S0
      =>nx10279);
   reg_Q_395 : dffr port map ( Q=>Q_395_EXMPLR, QB=>OPEN, D=>nx8788, CLK=>
      nx10157, R=>RST);
   ix8789 : mux21_ni port map ( Y=>nx8788, A0=>Q_395_EXMPLR, A1=>D(395), S0
      =>nx10279);
   reg_Q_396 : dffr port map ( Q=>Q_396_EXMPLR, QB=>OPEN, D=>nx8798, CLK=>
      nx10157, R=>RST);
   ix8799 : mux21_ni port map ( Y=>nx8798, A0=>Q_396_EXMPLR, A1=>D(396), S0
      =>nx10279);
   reg_Q_397 : dffr port map ( Q=>Q_397_EXMPLR, QB=>OPEN, D=>nx8808, CLK=>
      nx10157, R=>RST);
   ix8809 : mux21_ni port map ( Y=>nx8808, A0=>Q_397_EXMPLR, A1=>D(397), S0
      =>nx10279);
   reg_Q_398 : dffr port map ( Q=>Q_398_EXMPLR, QB=>OPEN, D=>nx8818, CLK=>
      nx10157, R=>RST);
   ix8819 : mux21_ni port map ( Y=>nx8818, A0=>Q_398_EXMPLR, A1=>D(398), S0
      =>nx10279);
   reg_Q_399 : dffr port map ( Q=>Q_399_EXMPLR, QB=>OPEN, D=>nx8828, CLK=>
      nx10159, R=>RST);
   ix8829 : mux21_ni port map ( Y=>nx8828, A0=>Q_399_EXMPLR, A1=>D(399), S0
      =>nx10281);
   ix10044 : inv02 port map ( Y=>nx10045, A=>CLK);
   ix10046 : inv02 port map ( Y=>nx10047, A=>nx10283);
   ix10048 : inv02 port map ( Y=>nx10049, A=>nx10283);
   ix10050 : inv02 port map ( Y=>nx10051, A=>nx10283);
   ix10052 : inv02 port map ( Y=>nx10053, A=>nx10283);
   ix10054 : inv02 port map ( Y=>nx10055, A=>nx10283);
   ix10056 : inv02 port map ( Y=>nx10057, A=>nx10283);
   ix10058 : inv02 port map ( Y=>nx10059, A=>nx10283);
   ix10060 : inv02 port map ( Y=>nx10061, A=>nx10285);
   ix10062 : inv02 port map ( Y=>nx10063, A=>nx10285);
   ix10064 : inv02 port map ( Y=>nx10065, A=>nx10285);
   ix10066 : inv02 port map ( Y=>nx10067, A=>nx10285);
   ix10068 : inv02 port map ( Y=>nx10069, A=>nx10285);
   ix10070 : inv02 port map ( Y=>nx10071, A=>nx10285);
   ix10072 : inv02 port map ( Y=>nx10073, A=>nx10285);
   ix10074 : inv02 port map ( Y=>nx10075, A=>nx10287);
   ix10076 : inv02 port map ( Y=>nx10077, A=>nx10287);
   ix10078 : inv02 port map ( Y=>nx10079, A=>nx10287);
   ix10080 : inv02 port map ( Y=>nx10081, A=>nx10287);
   ix10082 : inv02 port map ( Y=>nx10083, A=>nx10287);
   ix10084 : inv02 port map ( Y=>nx10085, A=>nx10287);
   ix10086 : inv02 port map ( Y=>nx10087, A=>nx10287);
   ix10088 : inv02 port map ( Y=>nx10089, A=>nx10289);
   ix10090 : inv02 port map ( Y=>nx10091, A=>nx10289);
   ix10092 : inv02 port map ( Y=>nx10093, A=>nx10289);
   ix10094 : inv02 port map ( Y=>nx10095, A=>nx10289);
   ix10096 : inv02 port map ( Y=>nx10097, A=>nx10289);
   ix10098 : inv02 port map ( Y=>nx10099, A=>nx10289);
   ix10100 : inv02 port map ( Y=>nx10101, A=>nx10289);
   ix10102 : inv02 port map ( Y=>nx10103, A=>nx10291);
   ix10104 : inv02 port map ( Y=>nx10105, A=>nx10291);
   ix10106 : inv02 port map ( Y=>nx10107, A=>nx10291);
   ix10108 : inv02 port map ( Y=>nx10109, A=>nx10291);
   ix10110 : inv02 port map ( Y=>nx10111, A=>nx10291);
   ix10112 : inv02 port map ( Y=>nx10113, A=>nx10291);
   ix10114 : inv02 port map ( Y=>nx10115, A=>nx10291);
   ix10116 : inv02 port map ( Y=>nx10117, A=>nx10293);
   ix10118 : inv02 port map ( Y=>nx10119, A=>nx10293);
   ix10120 : inv02 port map ( Y=>nx10121, A=>nx10293);
   ix10122 : inv02 port map ( Y=>nx10123, A=>nx10293);
   ix10124 : inv02 port map ( Y=>nx10125, A=>nx10293);
   ix10126 : inv02 port map ( Y=>nx10127, A=>nx10293);
   ix10128 : inv02 port map ( Y=>nx10129, A=>nx10293);
   ix10130 : inv02 port map ( Y=>nx10131, A=>nx10295);
   ix10132 : inv02 port map ( Y=>nx10133, A=>nx10295);
   ix10134 : inv02 port map ( Y=>nx10135, A=>nx10295);
   ix10136 : inv02 port map ( Y=>nx10137, A=>nx10295);
   ix10138 : inv02 port map ( Y=>nx10139, A=>nx10295);
   ix10140 : inv02 port map ( Y=>nx10141, A=>nx10295);
   ix10142 : inv02 port map ( Y=>nx10143, A=>nx10295);
   ix10144 : inv02 port map ( Y=>nx10145, A=>nx10297);
   ix10146 : inv02 port map ( Y=>nx10147, A=>nx10297);
   ix10148 : inv02 port map ( Y=>nx10149, A=>nx10297);
   ix10150 : inv02 port map ( Y=>nx10151, A=>nx10297);
   ix10152 : inv02 port map ( Y=>nx10153, A=>nx10297);
   ix10154 : inv02 port map ( Y=>nx10155, A=>nx10297);
   ix10156 : inv02 port map ( Y=>nx10157, A=>nx10297);
   ix10158 : inv02 port map ( Y=>nx10159, A=>nx10299);
   ix10166 : inv02 port map ( Y=>nx10167, A=>nx10305);
   ix10168 : inv02 port map ( Y=>nx10169, A=>nx10305);
   ix10170 : inv02 port map ( Y=>nx10171, A=>nx10305);
   ix10172 : inv02 port map ( Y=>nx10173, A=>nx10305);
   ix10174 : inv02 port map ( Y=>nx10175, A=>nx10305);
   ix10176 : inv02 port map ( Y=>nx10177, A=>nx10305);
   ix10178 : inv02 port map ( Y=>nx10179, A=>nx10305);
   ix10180 : inv02 port map ( Y=>nx10181, A=>nx10307);
   ix10182 : inv02 port map ( Y=>nx10183, A=>nx10307);
   ix10184 : inv02 port map ( Y=>nx10185, A=>nx10307);
   ix10186 : inv02 port map ( Y=>nx10187, A=>nx10307);
   ix10188 : inv02 port map ( Y=>nx10189, A=>nx10307);
   ix10190 : inv02 port map ( Y=>nx10191, A=>nx10307);
   ix10192 : inv02 port map ( Y=>nx10193, A=>nx10307);
   ix10194 : inv02 port map ( Y=>nx10195, A=>nx10309);
   ix10196 : inv02 port map ( Y=>nx10197, A=>nx10309);
   ix10198 : inv02 port map ( Y=>nx10199, A=>nx10309);
   ix10200 : inv02 port map ( Y=>nx10201, A=>nx10309);
   ix10202 : inv02 port map ( Y=>nx10203, A=>nx10309);
   ix10204 : inv02 port map ( Y=>nx10205, A=>nx10309);
   ix10206 : inv02 port map ( Y=>nx10207, A=>nx10309);
   ix10208 : inv02 port map ( Y=>nx10209, A=>nx10311);
   ix10210 : inv02 port map ( Y=>nx10211, A=>nx10311);
   ix10212 : inv02 port map ( Y=>nx10213, A=>nx10311);
   ix10214 : inv02 port map ( Y=>nx10215, A=>nx10311);
   ix10216 : inv02 port map ( Y=>nx10217, A=>nx10311);
   ix10218 : inv02 port map ( Y=>nx10219, A=>nx10311);
   ix10220 : inv02 port map ( Y=>nx10221, A=>nx10311);
   ix10222 : inv02 port map ( Y=>nx10223, A=>nx10313);
   ix10224 : inv02 port map ( Y=>nx10225, A=>nx10313);
   ix10226 : inv02 port map ( Y=>nx10227, A=>nx10313);
   ix10228 : inv02 port map ( Y=>nx10229, A=>nx10313);
   ix10230 : inv02 port map ( Y=>nx10231, A=>nx10313);
   ix10232 : inv02 port map ( Y=>nx10233, A=>nx10313);
   ix10234 : inv02 port map ( Y=>nx10235, A=>nx10313);
   ix10236 : inv02 port map ( Y=>nx10237, A=>nx10315);
   ix10238 : inv02 port map ( Y=>nx10239, A=>nx10315);
   ix10240 : inv02 port map ( Y=>nx10241, A=>nx10315);
   ix10242 : inv02 port map ( Y=>nx10243, A=>nx10315);
   ix10244 : inv02 port map ( Y=>nx10245, A=>nx10315);
   ix10246 : inv02 port map ( Y=>nx10247, A=>nx10315);
   ix10248 : inv02 port map ( Y=>nx10249, A=>nx10315);
   ix10250 : inv02 port map ( Y=>nx10251, A=>nx10317);
   ix10252 : inv02 port map ( Y=>nx10253, A=>nx10317);
   ix10254 : inv02 port map ( Y=>nx10255, A=>nx10317);
   ix10256 : inv02 port map ( Y=>nx10257, A=>nx10317);
   ix10258 : inv02 port map ( Y=>nx10259, A=>nx10317);
   ix10260 : inv02 port map ( Y=>nx10261, A=>nx10317);
   ix10262 : inv02 port map ( Y=>nx10263, A=>nx10317);
   ix10264 : inv02 port map ( Y=>nx10265, A=>nx10319);
   ix10266 : inv02 port map ( Y=>nx10267, A=>nx10319);
   ix10268 : inv02 port map ( Y=>nx10269, A=>nx10319);
   ix10270 : inv02 port map ( Y=>nx10271, A=>nx10319);
   ix10272 : inv02 port map ( Y=>nx10273, A=>nx10319);
   ix10274 : inv02 port map ( Y=>nx10275, A=>nx10319);
   ix10276 : inv02 port map ( Y=>nx10277, A=>nx10319);
   ix10278 : inv02 port map ( Y=>nx10279, A=>nx10321);
   ix10280 : inv02 port map ( Y=>nx10281, A=>nx10321);
   ix10282 : inv02 port map ( Y=>nx10283, A=>nx10303);
   ix10284 : inv02 port map ( Y=>nx10285, A=>nx10303);
   ix10286 : inv02 port map ( Y=>nx10287, A=>nx10303);
   ix10288 : inv02 port map ( Y=>nx10289, A=>nx10303);
   ix10290 : inv02 port map ( Y=>nx10291, A=>nx10303);
   ix10292 : inv02 port map ( Y=>nx10293, A=>nx10303);
   ix10294 : inv02 port map ( Y=>nx10295, A=>nx10303);
   ix10296 : inv02 port map ( Y=>nx10297, A=>nx10045);
   ix10298 : inv02 port map ( Y=>nx10299, A=>nx10045);
   ix10300 : inv02 port map ( Y=>nx10301, A=>CLK);
   ix10302 : inv02 port map ( Y=>nx10303, A=>CLK);
   ix10304 : inv02 port map ( Y=>nx10305, A=>EN);
   ix10306 : inv02 port map ( Y=>nx10307, A=>nx10327);
   ix10308 : inv02 port map ( Y=>nx10309, A=>nx10327);
   ix10310 : inv02 port map ( Y=>nx10311, A=>nx10327);
   ix10312 : inv02 port map ( Y=>nx10313, A=>nx10327);
   ix10314 : inv02 port map ( Y=>nx10315, A=>nx10327);
   ix10316 : inv02 port map ( Y=>nx10317, A=>nx10329);
   ix10318 : inv02 port map ( Y=>nx10319, A=>nx10329);
   ix10320 : inv02 port map ( Y=>nx10321, A=>nx10329);
   ix10326 : inv01 port map ( Y=>nx10327, A=>nx10305);
   ix10328 : inv01 port map ( Y=>nx10329, A=>nx10305);
end Data_flow ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity ReadFilter is
   port (
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
      depthcounter : IN std_logic_vector (3 DOWNTO 0) ;
      FilterCounter : IN std_logic_vector (3 DOWNTO 0) ;
      Heightcounter : IN std_logic_vector (4 DOWNTO 0) ;
      FILTER : IN std_logic_vector (399 DOWNTO 0) ;
      FilterAddress : IN std_logic_vector (12 DOWNTO 0) ;
      msbNoOfFilters : IN std_logic ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      QImgStat : IN std_logic ;
      ACKF : IN std_logic ;
      IndicatorFilter : OUT std_logic_vector (0 DOWNTO 0) ;
      DMAAddress : OUT std_logic_vector (12 DOWNTO 0) ;
      UpdatedAddress : OUT std_logic_vector (12 DOWNTO 0) ;
      outFilter0 : OUT std_logic_vector (399 DOWNTO 0) ;
      outFilter1 : OUT std_logic_vector (399 DOWNTO 0) ;
      donttrust : OUT std_logic ;
      LastFilterIND : OUT std_logic ;
      LastHeightOut : OUT std_logic ;
      lastDepthOut : OUT std_logic) ;
end ReadFilter ;

architecture DATA_FLOW of ReadFilter is
   component my_nadder_4
      port (
         a : IN std_logic_vector (3 DOWNTO 0) ;
         b : IN std_logic_vector (3 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (3 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component my_nadder_5
      port (
         a : IN std_logic_vector (4 DOWNTO 0) ;
         b : IN std_logic_vector (4 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (4 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component nBitRegister_400
      port (
         D : IN std_logic_vector (399 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (399 DOWNTO 0)) ;
   end component ;
   component nBitRegister_1
      port (
         D : IN std_logic_vector (0 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (0 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component my_nadder_13
      port (
         a : IN std_logic_vector (12 DOWNTO 0) ;
         b : IN std_logic_vector (12 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (12 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal IndicatorFilter_0_EXMPLR, DFFCLK, newAddress_12, newAddress_11, 
      newAddress_10, newAddress_9, newAddress_8, newAddress_7, newAddress_6, 
      newAddress_5, newAddress_4, newAddress_3, newAddress_2, newAddress_1, 
      newAddress_0, depthminus_3, depthminus_2, depthminus_1, depthminus_0, 
      FilterMinus_3, FilterMinus_2, FilterMinus_1, FilterMinus_0, 
      Heightminus_4, Heightminus_3, Heightminus_2, Heightminus_1, 
      Heightminus_0, donttrust_EXMPLR, LastFilterIND_EXMPLR, filter1EN, 
      filter2EN, lastDepthOut_EXMPLR, IndRst, tristateAddEn, secOperand_12, 
      secOperand_3, NOT_IndicatorFilter_0, nx2, nx22, nx24, nx96, nx108, 
      nx120, nx130, nx1466, nx1469, nx1471, nx1473, nx1475, nx1477, nx1479, 
      nx1482, nx1484, nx1486, nx1488, nx1491, nx1493, nx1495, nx1497: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (3 downto 0 );

begin
   IndicatorFilter(0) <= IndicatorFilter_0_EXMPLR ;
   donttrust <= donttrust_EXMPLR ;
   LastFilterIND <= LastFilterIND_EXMPLR ;
   LastHeightOut <= donttrust_EXMPLR ;
   lastDepthOut <= lastDepthOut_EXMPLR ;
   adder2 : my_nadder_4 port map ( a(3)=>LayerInfo(12), a(2)=>LayerInfo(11), 
      a(1)=>LayerInfo(10), a(0)=>LayerInfo(9), b(3)=>secOperand_3, b(2)=>
      secOperand_3, b(1)=>secOperand_3, b(0)=>secOperand_3, cin=>
      secOperand_12, s(3)=>depthminus_3, s(2)=>depthminus_2, s(1)=>
      depthminus_1, s(0)=>depthminus_0, cout=>DANGLING(0));
   adder3 : my_nadder_5 port map ( a(4)=>LayerInfo(8), a(3)=>LayerInfo(7), 
      a(2)=>LayerInfo(6), a(1)=>LayerInfo(5), a(0)=>LayerInfo(4), b(4)=>
      secOperand_3, b(3)=>secOperand_3, b(2)=>secOperand_3, b(1)=>
      secOperand_3, b(0)=>secOperand_3, cin=>secOperand_12, s(4)=>
      Heightminus_4, s(3)=>Heightminus_3, s(2)=>Heightminus_2, s(1)=>
      Heightminus_1, s(0)=>Heightminus_0, cout=>DANGLING(1));
   adder4 : my_nadder_4 port map ( a(3)=>LayerInfo(3), a(2)=>LayerInfo(2), 
      a(1)=>LayerInfo(1), a(0)=>LayerInfo(0), b(3)=>secOperand_3, b(2)=>
      secOperand_3, b(1)=>secOperand_3, b(0)=>secOperand_3, cin=>
      secOperand_12, s(3)=>FilterMinus_3, s(2)=>FilterMinus_2, s(1)=>
      FilterMinus_1, s(0)=>FilterMinus_0, cout=>DANGLING(2));
   F0 : nBitRegister_400 port map ( D(399)=>FILTER(399), D(398)=>FILTER(398), 
      D(397)=>FILTER(397), D(396)=>FILTER(396), D(395)=>FILTER(395), D(394)
      =>FILTER(394), D(393)=>FILTER(393), D(392)=>FILTER(392), D(391)=>
      FILTER(391), D(390)=>FILTER(390), D(389)=>FILTER(389), D(388)=>
      FILTER(388), D(387)=>FILTER(387), D(386)=>FILTER(386), D(385)=>
      FILTER(385), D(384)=>FILTER(384), D(383)=>FILTER(383), D(382)=>
      FILTER(382), D(381)=>FILTER(381), D(380)=>FILTER(380), D(379)=>
      FILTER(379), D(378)=>FILTER(378), D(377)=>FILTER(377), D(376)=>
      FILTER(376), D(375)=>FILTER(375), D(374)=>FILTER(374), D(373)=>
      FILTER(373), D(372)=>FILTER(372), D(371)=>FILTER(371), D(370)=>
      FILTER(370), D(369)=>FILTER(369), D(368)=>FILTER(368), D(367)=>
      FILTER(367), D(366)=>FILTER(366), D(365)=>FILTER(365), D(364)=>
      FILTER(364), D(363)=>FILTER(363), D(362)=>FILTER(362), D(361)=>
      FILTER(361), D(360)=>FILTER(360), D(359)=>FILTER(359), D(358)=>
      FILTER(358), D(357)=>FILTER(357), D(356)=>FILTER(356), D(355)=>
      FILTER(355), D(354)=>FILTER(354), D(353)=>FILTER(353), D(352)=>
      FILTER(352), D(351)=>FILTER(351), D(350)=>FILTER(350), D(349)=>
      FILTER(349), D(348)=>FILTER(348), D(347)=>FILTER(347), D(346)=>
      FILTER(346), D(345)=>FILTER(345), D(344)=>FILTER(344), D(343)=>
      FILTER(343), D(342)=>FILTER(342), D(341)=>FILTER(341), D(340)=>
      FILTER(340), D(339)=>FILTER(339), D(338)=>FILTER(338), D(337)=>
      FILTER(337), D(336)=>FILTER(336), D(335)=>FILTER(335), D(334)=>
      FILTER(334), D(333)=>FILTER(333), D(332)=>FILTER(332), D(331)=>
      FILTER(331), D(330)=>FILTER(330), D(329)=>FILTER(329), D(328)=>
      FILTER(328), D(327)=>FILTER(327), D(326)=>FILTER(326), D(325)=>
      FILTER(325), D(324)=>FILTER(324), D(323)=>FILTER(323), D(322)=>
      FILTER(322), D(321)=>FILTER(321), D(320)=>FILTER(320), D(319)=>
      FILTER(319), D(318)=>FILTER(318), D(317)=>FILTER(317), D(316)=>
      FILTER(316), D(315)=>FILTER(315), D(314)=>FILTER(314), D(313)=>
      FILTER(313), D(312)=>FILTER(312), D(311)=>FILTER(311), D(310)=>
      FILTER(310), D(309)=>FILTER(309), D(308)=>FILTER(308), D(307)=>
      FILTER(307), D(306)=>FILTER(306), D(305)=>FILTER(305), D(304)=>
      FILTER(304), D(303)=>FILTER(303), D(302)=>FILTER(302), D(301)=>
      FILTER(301), D(300)=>FILTER(300), D(299)=>FILTER(299), D(298)=>
      FILTER(298), D(297)=>FILTER(297), D(296)=>FILTER(296), D(295)=>
      FILTER(295), D(294)=>FILTER(294), D(293)=>FILTER(293), D(292)=>
      FILTER(292), D(291)=>FILTER(291), D(290)=>FILTER(290), D(289)=>
      FILTER(289), D(288)=>FILTER(288), D(287)=>FILTER(287), D(286)=>
      FILTER(286), D(285)=>FILTER(285), D(284)=>FILTER(284), D(283)=>
      FILTER(283), D(282)=>FILTER(282), D(281)=>FILTER(281), D(280)=>
      FILTER(280), D(279)=>FILTER(279), D(278)=>FILTER(278), D(277)=>
      FILTER(277), D(276)=>FILTER(276), D(275)=>FILTER(275), D(274)=>
      FILTER(274), D(273)=>FILTER(273), D(272)=>FILTER(272), D(271)=>
      FILTER(271), D(270)=>FILTER(270), D(269)=>FILTER(269), D(268)=>
      FILTER(268), D(267)=>FILTER(267), D(266)=>FILTER(266), D(265)=>
      FILTER(265), D(264)=>FILTER(264), D(263)=>FILTER(263), D(262)=>
      FILTER(262), D(261)=>FILTER(261), D(260)=>FILTER(260), D(259)=>
      FILTER(259), D(258)=>FILTER(258), D(257)=>FILTER(257), D(256)=>
      FILTER(256), D(255)=>FILTER(255), D(254)=>FILTER(254), D(253)=>
      FILTER(253), D(252)=>FILTER(252), D(251)=>FILTER(251), D(250)=>
      FILTER(250), D(249)=>FILTER(249), D(248)=>FILTER(248), D(247)=>
      FILTER(247), D(246)=>FILTER(246), D(245)=>FILTER(245), D(244)=>
      FILTER(244), D(243)=>FILTER(243), D(242)=>FILTER(242), D(241)=>
      FILTER(241), D(240)=>FILTER(240), D(239)=>FILTER(239), D(238)=>
      FILTER(238), D(237)=>FILTER(237), D(236)=>FILTER(236), D(235)=>
      FILTER(235), D(234)=>FILTER(234), D(233)=>FILTER(233), D(232)=>
      FILTER(232), D(231)=>FILTER(231), D(230)=>FILTER(230), D(229)=>
      FILTER(229), D(228)=>FILTER(228), D(227)=>FILTER(227), D(226)=>
      FILTER(226), D(225)=>FILTER(225), D(224)=>FILTER(224), D(223)=>
      FILTER(223), D(222)=>FILTER(222), D(221)=>FILTER(221), D(220)=>
      FILTER(220), D(219)=>FILTER(219), D(218)=>FILTER(218), D(217)=>
      FILTER(217), D(216)=>FILTER(216), D(215)=>FILTER(215), D(214)=>
      FILTER(214), D(213)=>FILTER(213), D(212)=>FILTER(212), D(211)=>
      FILTER(211), D(210)=>FILTER(210), D(209)=>FILTER(209), D(208)=>
      FILTER(208), D(207)=>FILTER(207), D(206)=>FILTER(206), D(205)=>
      FILTER(205), D(204)=>FILTER(204), D(203)=>FILTER(203), D(202)=>
      FILTER(202), D(201)=>FILTER(201), D(200)=>FILTER(200), D(199)=>
      FILTER(199), D(198)=>FILTER(198), D(197)=>FILTER(197), D(196)=>
      FILTER(196), D(195)=>FILTER(195), D(194)=>FILTER(194), D(193)=>
      FILTER(193), D(192)=>FILTER(192), D(191)=>FILTER(191), D(190)=>
      FILTER(190), D(189)=>FILTER(189), D(188)=>FILTER(188), D(187)=>
      FILTER(187), D(186)=>FILTER(186), D(185)=>FILTER(185), D(184)=>
      FILTER(184), D(183)=>FILTER(183), D(182)=>FILTER(182), D(181)=>
      FILTER(181), D(180)=>FILTER(180), D(179)=>FILTER(179), D(178)=>
      FILTER(178), D(177)=>FILTER(177), D(176)=>FILTER(176), D(175)=>
      FILTER(175), D(174)=>FILTER(174), D(173)=>FILTER(173), D(172)=>
      FILTER(172), D(171)=>FILTER(171), D(170)=>FILTER(170), D(169)=>
      FILTER(169), D(168)=>FILTER(168), D(167)=>FILTER(167), D(166)=>
      FILTER(166), D(165)=>FILTER(165), D(164)=>FILTER(164), D(163)=>
      FILTER(163), D(162)=>FILTER(162), D(161)=>FILTER(161), D(160)=>
      FILTER(160), D(159)=>FILTER(159), D(158)=>FILTER(158), D(157)=>
      FILTER(157), D(156)=>FILTER(156), D(155)=>FILTER(155), D(154)=>
      FILTER(154), D(153)=>FILTER(153), D(152)=>FILTER(152), D(151)=>
      FILTER(151), D(150)=>FILTER(150), D(149)=>FILTER(149), D(148)=>
      FILTER(148), D(147)=>FILTER(147), D(146)=>FILTER(146), D(145)=>
      FILTER(145), D(144)=>FILTER(144), D(143)=>FILTER(143), D(142)=>
      FILTER(142), D(141)=>FILTER(141), D(140)=>FILTER(140), D(139)=>
      FILTER(139), D(138)=>FILTER(138), D(137)=>FILTER(137), D(136)=>
      FILTER(136), D(135)=>FILTER(135), D(134)=>FILTER(134), D(133)=>
      FILTER(133), D(132)=>FILTER(132), D(131)=>FILTER(131), D(130)=>
      FILTER(130), D(129)=>FILTER(129), D(128)=>FILTER(128), D(127)=>
      FILTER(127), D(126)=>FILTER(126), D(125)=>FILTER(125), D(124)=>
      FILTER(124), D(123)=>FILTER(123), D(122)=>FILTER(122), D(121)=>
      FILTER(121), D(120)=>FILTER(120), D(119)=>FILTER(119), D(118)=>
      FILTER(118), D(117)=>FILTER(117), D(116)=>FILTER(116), D(115)=>
      FILTER(115), D(114)=>FILTER(114), D(113)=>FILTER(113), D(112)=>
      FILTER(112), D(111)=>FILTER(111), D(110)=>FILTER(110), D(109)=>
      FILTER(109), D(108)=>FILTER(108), D(107)=>FILTER(107), D(106)=>
      FILTER(106), D(105)=>FILTER(105), D(104)=>FILTER(104), D(103)=>
      FILTER(103), D(102)=>FILTER(102), D(101)=>FILTER(101), D(100)=>
      FILTER(100), D(99)=>FILTER(99), D(98)=>FILTER(98), D(97)=>FILTER(97), 
      D(96)=>FILTER(96), D(95)=>FILTER(95), D(94)=>FILTER(94), D(93)=>
      FILTER(93), D(92)=>FILTER(92), D(91)=>FILTER(91), D(90)=>FILTER(90), 
      D(89)=>FILTER(89), D(88)=>FILTER(88), D(87)=>FILTER(87), D(86)=>
      FILTER(86), D(85)=>FILTER(85), D(84)=>FILTER(84), D(83)=>FILTER(83), 
      D(82)=>FILTER(82), D(81)=>FILTER(81), D(80)=>FILTER(80), D(79)=>
      FILTER(79), D(78)=>FILTER(78), D(77)=>FILTER(77), D(76)=>FILTER(76), 
      D(75)=>FILTER(75), D(74)=>FILTER(74), D(73)=>FILTER(73), D(72)=>
      FILTER(72), D(71)=>FILTER(71), D(70)=>FILTER(70), D(69)=>FILTER(69), 
      D(68)=>FILTER(68), D(67)=>FILTER(67), D(66)=>FILTER(66), D(65)=>
      FILTER(65), D(64)=>FILTER(64), D(63)=>FILTER(63), D(62)=>FILTER(62), 
      D(61)=>FILTER(61), D(60)=>FILTER(60), D(59)=>FILTER(59), D(58)=>
      FILTER(58), D(57)=>FILTER(57), D(56)=>FILTER(56), D(55)=>FILTER(55), 
      D(54)=>FILTER(54), D(53)=>FILTER(53), D(52)=>FILTER(52), D(51)=>
      FILTER(51), D(50)=>FILTER(50), D(49)=>FILTER(49), D(48)=>FILTER(48), 
      D(47)=>FILTER(47), D(46)=>FILTER(46), D(45)=>FILTER(45), D(44)=>
      FILTER(44), D(43)=>FILTER(43), D(42)=>FILTER(42), D(41)=>FILTER(41), 
      D(40)=>FILTER(40), D(39)=>FILTER(39), D(38)=>FILTER(38), D(37)=>
      FILTER(37), D(36)=>FILTER(36), D(35)=>FILTER(35), D(34)=>FILTER(34), 
      D(33)=>FILTER(33), D(32)=>FILTER(32), D(31)=>FILTER(31), D(30)=>
      FILTER(30), D(29)=>FILTER(29), D(28)=>FILTER(28), D(27)=>FILTER(27), 
      D(26)=>FILTER(26), D(25)=>FILTER(25), D(24)=>FILTER(24), D(23)=>
      FILTER(23), D(22)=>FILTER(22), D(21)=>FILTER(21), D(20)=>FILTER(20), 
      D(19)=>FILTER(19), D(18)=>FILTER(18), D(17)=>FILTER(17), D(16)=>
      FILTER(16), D(15)=>FILTER(15), D(14)=>FILTER(14), D(13)=>FILTER(13), 
      D(12)=>FILTER(12), D(11)=>FILTER(11), D(10)=>FILTER(10), D(9)=>
      FILTER(9), D(8)=>FILTER(8), D(7)=>FILTER(7), D(6)=>FILTER(6), D(5)=>
      FILTER(5), D(4)=>FILTER(4), D(3)=>FILTER(3), D(2)=>FILTER(2), D(1)=>
      FILTER(1), D(0)=>FILTER(0), CLK=>CLK, RST=>RST, EN=>filter1EN, Q(399)
      =>outFilter0(399), Q(398)=>outFilter0(398), Q(397)=>outFilter0(397), 
      Q(396)=>outFilter0(396), Q(395)=>outFilter0(395), Q(394)=>
      outFilter0(394), Q(393)=>outFilter0(393), Q(392)=>outFilter0(392), 
      Q(391)=>outFilter0(391), Q(390)=>outFilter0(390), Q(389)=>
      outFilter0(389), Q(388)=>outFilter0(388), Q(387)=>outFilter0(387), 
      Q(386)=>outFilter0(386), Q(385)=>outFilter0(385), Q(384)=>
      outFilter0(384), Q(383)=>outFilter0(383), Q(382)=>outFilter0(382), 
      Q(381)=>outFilter0(381), Q(380)=>outFilter0(380), Q(379)=>
      outFilter0(379), Q(378)=>outFilter0(378), Q(377)=>outFilter0(377), 
      Q(376)=>outFilter0(376), Q(375)=>outFilter0(375), Q(374)=>
      outFilter0(374), Q(373)=>outFilter0(373), Q(372)=>outFilter0(372), 
      Q(371)=>outFilter0(371), Q(370)=>outFilter0(370), Q(369)=>
      outFilter0(369), Q(368)=>outFilter0(368), Q(367)=>outFilter0(367), 
      Q(366)=>outFilter0(366), Q(365)=>outFilter0(365), Q(364)=>
      outFilter0(364), Q(363)=>outFilter0(363), Q(362)=>outFilter0(362), 
      Q(361)=>outFilter0(361), Q(360)=>outFilter0(360), Q(359)=>
      outFilter0(359), Q(358)=>outFilter0(358), Q(357)=>outFilter0(357), 
      Q(356)=>outFilter0(356), Q(355)=>outFilter0(355), Q(354)=>
      outFilter0(354), Q(353)=>outFilter0(353), Q(352)=>outFilter0(352), 
      Q(351)=>outFilter0(351), Q(350)=>outFilter0(350), Q(349)=>
      outFilter0(349), Q(348)=>outFilter0(348), Q(347)=>outFilter0(347), 
      Q(346)=>outFilter0(346), Q(345)=>outFilter0(345), Q(344)=>
      outFilter0(344), Q(343)=>outFilter0(343), Q(342)=>outFilter0(342), 
      Q(341)=>outFilter0(341), Q(340)=>outFilter0(340), Q(339)=>
      outFilter0(339), Q(338)=>outFilter0(338), Q(337)=>outFilter0(337), 
      Q(336)=>outFilter0(336), Q(335)=>outFilter0(335), Q(334)=>
      outFilter0(334), Q(333)=>outFilter0(333), Q(332)=>outFilter0(332), 
      Q(331)=>outFilter0(331), Q(330)=>outFilter0(330), Q(329)=>
      outFilter0(329), Q(328)=>outFilter0(328), Q(327)=>outFilter0(327), 
      Q(326)=>outFilter0(326), Q(325)=>outFilter0(325), Q(324)=>
      outFilter0(324), Q(323)=>outFilter0(323), Q(322)=>outFilter0(322), 
      Q(321)=>outFilter0(321), Q(320)=>outFilter0(320), Q(319)=>
      outFilter0(319), Q(318)=>outFilter0(318), Q(317)=>outFilter0(317), 
      Q(316)=>outFilter0(316), Q(315)=>outFilter0(315), Q(314)=>
      outFilter0(314), Q(313)=>outFilter0(313), Q(312)=>outFilter0(312), 
      Q(311)=>outFilter0(311), Q(310)=>outFilter0(310), Q(309)=>
      outFilter0(309), Q(308)=>outFilter0(308), Q(307)=>outFilter0(307), 
      Q(306)=>outFilter0(306), Q(305)=>outFilter0(305), Q(304)=>
      outFilter0(304), Q(303)=>outFilter0(303), Q(302)=>outFilter0(302), 
      Q(301)=>outFilter0(301), Q(300)=>outFilter0(300), Q(299)=>
      outFilter0(299), Q(298)=>outFilter0(298), Q(297)=>outFilter0(297), 
      Q(296)=>outFilter0(296), Q(295)=>outFilter0(295), Q(294)=>
      outFilter0(294), Q(293)=>outFilter0(293), Q(292)=>outFilter0(292), 
      Q(291)=>outFilter0(291), Q(290)=>outFilter0(290), Q(289)=>
      outFilter0(289), Q(288)=>outFilter0(288), Q(287)=>outFilter0(287), 
      Q(286)=>outFilter0(286), Q(285)=>outFilter0(285), Q(284)=>
      outFilter0(284), Q(283)=>outFilter0(283), Q(282)=>outFilter0(282), 
      Q(281)=>outFilter0(281), Q(280)=>outFilter0(280), Q(279)=>
      outFilter0(279), Q(278)=>outFilter0(278), Q(277)=>outFilter0(277), 
      Q(276)=>outFilter0(276), Q(275)=>outFilter0(275), Q(274)=>
      outFilter0(274), Q(273)=>outFilter0(273), Q(272)=>outFilter0(272), 
      Q(271)=>outFilter0(271), Q(270)=>outFilter0(270), Q(269)=>
      outFilter0(269), Q(268)=>outFilter0(268), Q(267)=>outFilter0(267), 
      Q(266)=>outFilter0(266), Q(265)=>outFilter0(265), Q(264)=>
      outFilter0(264), Q(263)=>outFilter0(263), Q(262)=>outFilter0(262), 
      Q(261)=>outFilter0(261), Q(260)=>outFilter0(260), Q(259)=>
      outFilter0(259), Q(258)=>outFilter0(258), Q(257)=>outFilter0(257), 
      Q(256)=>outFilter0(256), Q(255)=>outFilter0(255), Q(254)=>
      outFilter0(254), Q(253)=>outFilter0(253), Q(252)=>outFilter0(252), 
      Q(251)=>outFilter0(251), Q(250)=>outFilter0(250), Q(249)=>
      outFilter0(249), Q(248)=>outFilter0(248), Q(247)=>outFilter0(247), 
      Q(246)=>outFilter0(246), Q(245)=>outFilter0(245), Q(244)=>
      outFilter0(244), Q(243)=>outFilter0(243), Q(242)=>outFilter0(242), 
      Q(241)=>outFilter0(241), Q(240)=>outFilter0(240), Q(239)=>
      outFilter0(239), Q(238)=>outFilter0(238), Q(237)=>outFilter0(237), 
      Q(236)=>outFilter0(236), Q(235)=>outFilter0(235), Q(234)=>
      outFilter0(234), Q(233)=>outFilter0(233), Q(232)=>outFilter0(232), 
      Q(231)=>outFilter0(231), Q(230)=>outFilter0(230), Q(229)=>
      outFilter0(229), Q(228)=>outFilter0(228), Q(227)=>outFilter0(227), 
      Q(226)=>outFilter0(226), Q(225)=>outFilter0(225), Q(224)=>
      outFilter0(224), Q(223)=>outFilter0(223), Q(222)=>outFilter0(222), 
      Q(221)=>outFilter0(221), Q(220)=>outFilter0(220), Q(219)=>
      outFilter0(219), Q(218)=>outFilter0(218), Q(217)=>outFilter0(217), 
      Q(216)=>outFilter0(216), Q(215)=>outFilter0(215), Q(214)=>
      outFilter0(214), Q(213)=>outFilter0(213), Q(212)=>outFilter0(212), 
      Q(211)=>outFilter0(211), Q(210)=>outFilter0(210), Q(209)=>
      outFilter0(209), Q(208)=>outFilter0(208), Q(207)=>outFilter0(207), 
      Q(206)=>outFilter0(206), Q(205)=>outFilter0(205), Q(204)=>
      outFilter0(204), Q(203)=>outFilter0(203), Q(202)=>outFilter0(202), 
      Q(201)=>outFilter0(201), Q(200)=>outFilter0(200), Q(199)=>
      outFilter0(199), Q(198)=>outFilter0(198), Q(197)=>outFilter0(197), 
      Q(196)=>outFilter0(196), Q(195)=>outFilter0(195), Q(194)=>
      outFilter0(194), Q(193)=>outFilter0(193), Q(192)=>outFilter0(192), 
      Q(191)=>outFilter0(191), Q(190)=>outFilter0(190), Q(189)=>
      outFilter0(189), Q(188)=>outFilter0(188), Q(187)=>outFilter0(187), 
      Q(186)=>outFilter0(186), Q(185)=>outFilter0(185), Q(184)=>
      outFilter0(184), Q(183)=>outFilter0(183), Q(182)=>outFilter0(182), 
      Q(181)=>outFilter0(181), Q(180)=>outFilter0(180), Q(179)=>
      outFilter0(179), Q(178)=>outFilter0(178), Q(177)=>outFilter0(177), 
      Q(176)=>outFilter0(176), Q(175)=>outFilter0(175), Q(174)=>
      outFilter0(174), Q(173)=>outFilter0(173), Q(172)=>outFilter0(172), 
      Q(171)=>outFilter0(171), Q(170)=>outFilter0(170), Q(169)=>
      outFilter0(169), Q(168)=>outFilter0(168), Q(167)=>outFilter0(167), 
      Q(166)=>outFilter0(166), Q(165)=>outFilter0(165), Q(164)=>
      outFilter0(164), Q(163)=>outFilter0(163), Q(162)=>outFilter0(162), 
      Q(161)=>outFilter0(161), Q(160)=>outFilter0(160), Q(159)=>
      outFilter0(159), Q(158)=>outFilter0(158), Q(157)=>outFilter0(157), 
      Q(156)=>outFilter0(156), Q(155)=>outFilter0(155), Q(154)=>
      outFilter0(154), Q(153)=>outFilter0(153), Q(152)=>outFilter0(152), 
      Q(151)=>outFilter0(151), Q(150)=>outFilter0(150), Q(149)=>
      outFilter0(149), Q(148)=>outFilter0(148), Q(147)=>outFilter0(147), 
      Q(146)=>outFilter0(146), Q(145)=>outFilter0(145), Q(144)=>
      outFilter0(144), Q(143)=>outFilter0(143), Q(142)=>outFilter0(142), 
      Q(141)=>outFilter0(141), Q(140)=>outFilter0(140), Q(139)=>
      outFilter0(139), Q(138)=>outFilter0(138), Q(137)=>outFilter0(137), 
      Q(136)=>outFilter0(136), Q(135)=>outFilter0(135), Q(134)=>
      outFilter0(134), Q(133)=>outFilter0(133), Q(132)=>outFilter0(132), 
      Q(131)=>outFilter0(131), Q(130)=>outFilter0(130), Q(129)=>
      outFilter0(129), Q(128)=>outFilter0(128), Q(127)=>outFilter0(127), 
      Q(126)=>outFilter0(126), Q(125)=>outFilter0(125), Q(124)=>
      outFilter0(124), Q(123)=>outFilter0(123), Q(122)=>outFilter0(122), 
      Q(121)=>outFilter0(121), Q(120)=>outFilter0(120), Q(119)=>
      outFilter0(119), Q(118)=>outFilter0(118), Q(117)=>outFilter0(117), 
      Q(116)=>outFilter0(116), Q(115)=>outFilter0(115), Q(114)=>
      outFilter0(114), Q(113)=>outFilter0(113), Q(112)=>outFilter0(112), 
      Q(111)=>outFilter0(111), Q(110)=>outFilter0(110), Q(109)=>
      outFilter0(109), Q(108)=>outFilter0(108), Q(107)=>outFilter0(107), 
      Q(106)=>outFilter0(106), Q(105)=>outFilter0(105), Q(104)=>
      outFilter0(104), Q(103)=>outFilter0(103), Q(102)=>outFilter0(102), 
      Q(101)=>outFilter0(101), Q(100)=>outFilter0(100), Q(99)=>
      outFilter0(99), Q(98)=>outFilter0(98), Q(97)=>outFilter0(97), Q(96)=>
      outFilter0(96), Q(95)=>outFilter0(95), Q(94)=>outFilter0(94), Q(93)=>
      outFilter0(93), Q(92)=>outFilter0(92), Q(91)=>outFilter0(91), Q(90)=>
      outFilter0(90), Q(89)=>outFilter0(89), Q(88)=>outFilter0(88), Q(87)=>
      outFilter0(87), Q(86)=>outFilter0(86), Q(85)=>outFilter0(85), Q(84)=>
      outFilter0(84), Q(83)=>outFilter0(83), Q(82)=>outFilter0(82), Q(81)=>
      outFilter0(81), Q(80)=>outFilter0(80), Q(79)=>outFilter0(79), Q(78)=>
      outFilter0(78), Q(77)=>outFilter0(77), Q(76)=>outFilter0(76), Q(75)=>
      outFilter0(75), Q(74)=>outFilter0(74), Q(73)=>outFilter0(73), Q(72)=>
      outFilter0(72), Q(71)=>outFilter0(71), Q(70)=>outFilter0(70), Q(69)=>
      outFilter0(69), Q(68)=>outFilter0(68), Q(67)=>outFilter0(67), Q(66)=>
      outFilter0(66), Q(65)=>outFilter0(65), Q(64)=>outFilter0(64), Q(63)=>
      outFilter0(63), Q(62)=>outFilter0(62), Q(61)=>outFilter0(61), Q(60)=>
      outFilter0(60), Q(59)=>outFilter0(59), Q(58)=>outFilter0(58), Q(57)=>
      outFilter0(57), Q(56)=>outFilter0(56), Q(55)=>outFilter0(55), Q(54)=>
      outFilter0(54), Q(53)=>outFilter0(53), Q(52)=>outFilter0(52), Q(51)=>
      outFilter0(51), Q(50)=>outFilter0(50), Q(49)=>outFilter0(49), Q(48)=>
      outFilter0(48), Q(47)=>outFilter0(47), Q(46)=>outFilter0(46), Q(45)=>
      outFilter0(45), Q(44)=>outFilter0(44), Q(43)=>outFilter0(43), Q(42)=>
      outFilter0(42), Q(41)=>outFilter0(41), Q(40)=>outFilter0(40), Q(39)=>
      outFilter0(39), Q(38)=>outFilter0(38), Q(37)=>outFilter0(37), Q(36)=>
      outFilter0(36), Q(35)=>outFilter0(35), Q(34)=>outFilter0(34), Q(33)=>
      outFilter0(33), Q(32)=>outFilter0(32), Q(31)=>outFilter0(31), Q(30)=>
      outFilter0(30), Q(29)=>outFilter0(29), Q(28)=>outFilter0(28), Q(27)=>
      outFilter0(27), Q(26)=>outFilter0(26), Q(25)=>outFilter0(25), Q(24)=>
      outFilter0(24), Q(23)=>outFilter0(23), Q(22)=>outFilter0(22), Q(21)=>
      outFilter0(21), Q(20)=>outFilter0(20), Q(19)=>outFilter0(19), Q(18)=>
      outFilter0(18), Q(17)=>outFilter0(17), Q(16)=>outFilter0(16), Q(15)=>
      outFilter0(15), Q(14)=>outFilter0(14), Q(13)=>outFilter0(13), Q(12)=>
      outFilter0(12), Q(11)=>outFilter0(11), Q(10)=>outFilter0(10), Q(9)=>
      outFilter0(9), Q(8)=>outFilter0(8), Q(7)=>outFilter0(7), Q(6)=>
      outFilter0(6), Q(5)=>outFilter0(5), Q(4)=>outFilter0(4), Q(3)=>
      outFilter0(3), Q(2)=>outFilter0(2), Q(1)=>outFilter0(1), Q(0)=>
      outFilter0(0));
   F1 : nBitRegister_400 port map ( D(399)=>FILTER(399), D(398)=>FILTER(398), 
      D(397)=>FILTER(397), D(396)=>FILTER(396), D(395)=>FILTER(395), D(394)
      =>FILTER(394), D(393)=>FILTER(393), D(392)=>FILTER(392), D(391)=>
      FILTER(391), D(390)=>FILTER(390), D(389)=>FILTER(389), D(388)=>
      FILTER(388), D(387)=>FILTER(387), D(386)=>FILTER(386), D(385)=>
      FILTER(385), D(384)=>FILTER(384), D(383)=>FILTER(383), D(382)=>
      FILTER(382), D(381)=>FILTER(381), D(380)=>FILTER(380), D(379)=>
      FILTER(379), D(378)=>FILTER(378), D(377)=>FILTER(377), D(376)=>
      FILTER(376), D(375)=>FILTER(375), D(374)=>FILTER(374), D(373)=>
      FILTER(373), D(372)=>FILTER(372), D(371)=>FILTER(371), D(370)=>
      FILTER(370), D(369)=>FILTER(369), D(368)=>FILTER(368), D(367)=>
      FILTER(367), D(366)=>FILTER(366), D(365)=>FILTER(365), D(364)=>
      FILTER(364), D(363)=>FILTER(363), D(362)=>FILTER(362), D(361)=>
      FILTER(361), D(360)=>FILTER(360), D(359)=>FILTER(359), D(358)=>
      FILTER(358), D(357)=>FILTER(357), D(356)=>FILTER(356), D(355)=>
      FILTER(355), D(354)=>FILTER(354), D(353)=>FILTER(353), D(352)=>
      FILTER(352), D(351)=>FILTER(351), D(350)=>FILTER(350), D(349)=>
      FILTER(349), D(348)=>FILTER(348), D(347)=>FILTER(347), D(346)=>
      FILTER(346), D(345)=>FILTER(345), D(344)=>FILTER(344), D(343)=>
      FILTER(343), D(342)=>FILTER(342), D(341)=>FILTER(341), D(340)=>
      FILTER(340), D(339)=>FILTER(339), D(338)=>FILTER(338), D(337)=>
      FILTER(337), D(336)=>FILTER(336), D(335)=>FILTER(335), D(334)=>
      FILTER(334), D(333)=>FILTER(333), D(332)=>FILTER(332), D(331)=>
      FILTER(331), D(330)=>FILTER(330), D(329)=>FILTER(329), D(328)=>
      FILTER(328), D(327)=>FILTER(327), D(326)=>FILTER(326), D(325)=>
      FILTER(325), D(324)=>FILTER(324), D(323)=>FILTER(323), D(322)=>
      FILTER(322), D(321)=>FILTER(321), D(320)=>FILTER(320), D(319)=>
      FILTER(319), D(318)=>FILTER(318), D(317)=>FILTER(317), D(316)=>
      FILTER(316), D(315)=>FILTER(315), D(314)=>FILTER(314), D(313)=>
      FILTER(313), D(312)=>FILTER(312), D(311)=>FILTER(311), D(310)=>
      FILTER(310), D(309)=>FILTER(309), D(308)=>FILTER(308), D(307)=>
      FILTER(307), D(306)=>FILTER(306), D(305)=>FILTER(305), D(304)=>
      FILTER(304), D(303)=>FILTER(303), D(302)=>FILTER(302), D(301)=>
      FILTER(301), D(300)=>FILTER(300), D(299)=>FILTER(299), D(298)=>
      FILTER(298), D(297)=>FILTER(297), D(296)=>FILTER(296), D(295)=>
      FILTER(295), D(294)=>FILTER(294), D(293)=>FILTER(293), D(292)=>
      FILTER(292), D(291)=>FILTER(291), D(290)=>FILTER(290), D(289)=>
      FILTER(289), D(288)=>FILTER(288), D(287)=>FILTER(287), D(286)=>
      FILTER(286), D(285)=>FILTER(285), D(284)=>FILTER(284), D(283)=>
      FILTER(283), D(282)=>FILTER(282), D(281)=>FILTER(281), D(280)=>
      FILTER(280), D(279)=>FILTER(279), D(278)=>FILTER(278), D(277)=>
      FILTER(277), D(276)=>FILTER(276), D(275)=>FILTER(275), D(274)=>
      FILTER(274), D(273)=>FILTER(273), D(272)=>FILTER(272), D(271)=>
      FILTER(271), D(270)=>FILTER(270), D(269)=>FILTER(269), D(268)=>
      FILTER(268), D(267)=>FILTER(267), D(266)=>FILTER(266), D(265)=>
      FILTER(265), D(264)=>FILTER(264), D(263)=>FILTER(263), D(262)=>
      FILTER(262), D(261)=>FILTER(261), D(260)=>FILTER(260), D(259)=>
      FILTER(259), D(258)=>FILTER(258), D(257)=>FILTER(257), D(256)=>
      FILTER(256), D(255)=>FILTER(255), D(254)=>FILTER(254), D(253)=>
      FILTER(253), D(252)=>FILTER(252), D(251)=>FILTER(251), D(250)=>
      FILTER(250), D(249)=>FILTER(249), D(248)=>FILTER(248), D(247)=>
      FILTER(247), D(246)=>FILTER(246), D(245)=>FILTER(245), D(244)=>
      FILTER(244), D(243)=>FILTER(243), D(242)=>FILTER(242), D(241)=>
      FILTER(241), D(240)=>FILTER(240), D(239)=>FILTER(239), D(238)=>
      FILTER(238), D(237)=>FILTER(237), D(236)=>FILTER(236), D(235)=>
      FILTER(235), D(234)=>FILTER(234), D(233)=>FILTER(233), D(232)=>
      FILTER(232), D(231)=>FILTER(231), D(230)=>FILTER(230), D(229)=>
      FILTER(229), D(228)=>FILTER(228), D(227)=>FILTER(227), D(226)=>
      FILTER(226), D(225)=>FILTER(225), D(224)=>FILTER(224), D(223)=>
      FILTER(223), D(222)=>FILTER(222), D(221)=>FILTER(221), D(220)=>
      FILTER(220), D(219)=>FILTER(219), D(218)=>FILTER(218), D(217)=>
      FILTER(217), D(216)=>FILTER(216), D(215)=>FILTER(215), D(214)=>
      FILTER(214), D(213)=>FILTER(213), D(212)=>FILTER(212), D(211)=>
      FILTER(211), D(210)=>FILTER(210), D(209)=>FILTER(209), D(208)=>
      FILTER(208), D(207)=>FILTER(207), D(206)=>FILTER(206), D(205)=>
      FILTER(205), D(204)=>FILTER(204), D(203)=>FILTER(203), D(202)=>
      FILTER(202), D(201)=>FILTER(201), D(200)=>FILTER(200), D(199)=>
      FILTER(199), D(198)=>FILTER(198), D(197)=>FILTER(197), D(196)=>
      FILTER(196), D(195)=>FILTER(195), D(194)=>FILTER(194), D(193)=>
      FILTER(193), D(192)=>FILTER(192), D(191)=>FILTER(191), D(190)=>
      FILTER(190), D(189)=>FILTER(189), D(188)=>FILTER(188), D(187)=>
      FILTER(187), D(186)=>FILTER(186), D(185)=>FILTER(185), D(184)=>
      FILTER(184), D(183)=>FILTER(183), D(182)=>FILTER(182), D(181)=>
      FILTER(181), D(180)=>FILTER(180), D(179)=>FILTER(179), D(178)=>
      FILTER(178), D(177)=>FILTER(177), D(176)=>FILTER(176), D(175)=>
      FILTER(175), D(174)=>FILTER(174), D(173)=>FILTER(173), D(172)=>
      FILTER(172), D(171)=>FILTER(171), D(170)=>FILTER(170), D(169)=>
      FILTER(169), D(168)=>FILTER(168), D(167)=>FILTER(167), D(166)=>
      FILTER(166), D(165)=>FILTER(165), D(164)=>FILTER(164), D(163)=>
      FILTER(163), D(162)=>FILTER(162), D(161)=>FILTER(161), D(160)=>
      FILTER(160), D(159)=>FILTER(159), D(158)=>FILTER(158), D(157)=>
      FILTER(157), D(156)=>FILTER(156), D(155)=>FILTER(155), D(154)=>
      FILTER(154), D(153)=>FILTER(153), D(152)=>FILTER(152), D(151)=>
      FILTER(151), D(150)=>FILTER(150), D(149)=>FILTER(149), D(148)=>
      FILTER(148), D(147)=>FILTER(147), D(146)=>FILTER(146), D(145)=>
      FILTER(145), D(144)=>FILTER(144), D(143)=>FILTER(143), D(142)=>
      FILTER(142), D(141)=>FILTER(141), D(140)=>FILTER(140), D(139)=>
      FILTER(139), D(138)=>FILTER(138), D(137)=>FILTER(137), D(136)=>
      FILTER(136), D(135)=>FILTER(135), D(134)=>FILTER(134), D(133)=>
      FILTER(133), D(132)=>FILTER(132), D(131)=>FILTER(131), D(130)=>
      FILTER(130), D(129)=>FILTER(129), D(128)=>FILTER(128), D(127)=>
      FILTER(127), D(126)=>FILTER(126), D(125)=>FILTER(125), D(124)=>
      FILTER(124), D(123)=>FILTER(123), D(122)=>FILTER(122), D(121)=>
      FILTER(121), D(120)=>FILTER(120), D(119)=>FILTER(119), D(118)=>
      FILTER(118), D(117)=>FILTER(117), D(116)=>FILTER(116), D(115)=>
      FILTER(115), D(114)=>FILTER(114), D(113)=>FILTER(113), D(112)=>
      FILTER(112), D(111)=>FILTER(111), D(110)=>FILTER(110), D(109)=>
      FILTER(109), D(108)=>FILTER(108), D(107)=>FILTER(107), D(106)=>
      FILTER(106), D(105)=>FILTER(105), D(104)=>FILTER(104), D(103)=>
      FILTER(103), D(102)=>FILTER(102), D(101)=>FILTER(101), D(100)=>
      FILTER(100), D(99)=>FILTER(99), D(98)=>FILTER(98), D(97)=>FILTER(97), 
      D(96)=>FILTER(96), D(95)=>FILTER(95), D(94)=>FILTER(94), D(93)=>
      FILTER(93), D(92)=>FILTER(92), D(91)=>FILTER(91), D(90)=>FILTER(90), 
      D(89)=>FILTER(89), D(88)=>FILTER(88), D(87)=>FILTER(87), D(86)=>
      FILTER(86), D(85)=>FILTER(85), D(84)=>FILTER(84), D(83)=>FILTER(83), 
      D(82)=>FILTER(82), D(81)=>FILTER(81), D(80)=>FILTER(80), D(79)=>
      FILTER(79), D(78)=>FILTER(78), D(77)=>FILTER(77), D(76)=>FILTER(76), 
      D(75)=>FILTER(75), D(74)=>FILTER(74), D(73)=>FILTER(73), D(72)=>
      FILTER(72), D(71)=>FILTER(71), D(70)=>FILTER(70), D(69)=>FILTER(69), 
      D(68)=>FILTER(68), D(67)=>FILTER(67), D(66)=>FILTER(66), D(65)=>
      FILTER(65), D(64)=>FILTER(64), D(63)=>FILTER(63), D(62)=>FILTER(62), 
      D(61)=>FILTER(61), D(60)=>FILTER(60), D(59)=>FILTER(59), D(58)=>
      FILTER(58), D(57)=>FILTER(57), D(56)=>FILTER(56), D(55)=>FILTER(55), 
      D(54)=>FILTER(54), D(53)=>FILTER(53), D(52)=>FILTER(52), D(51)=>
      FILTER(51), D(50)=>FILTER(50), D(49)=>FILTER(49), D(48)=>FILTER(48), 
      D(47)=>FILTER(47), D(46)=>FILTER(46), D(45)=>FILTER(45), D(44)=>
      FILTER(44), D(43)=>FILTER(43), D(42)=>FILTER(42), D(41)=>FILTER(41), 
      D(40)=>FILTER(40), D(39)=>FILTER(39), D(38)=>FILTER(38), D(37)=>
      FILTER(37), D(36)=>FILTER(36), D(35)=>FILTER(35), D(34)=>FILTER(34), 
      D(33)=>FILTER(33), D(32)=>FILTER(32), D(31)=>FILTER(31), D(30)=>
      FILTER(30), D(29)=>FILTER(29), D(28)=>FILTER(28), D(27)=>FILTER(27), 
      D(26)=>FILTER(26), D(25)=>FILTER(25), D(24)=>FILTER(24), D(23)=>
      FILTER(23), D(22)=>FILTER(22), D(21)=>FILTER(21), D(20)=>FILTER(20), 
      D(19)=>FILTER(19), D(18)=>FILTER(18), D(17)=>FILTER(17), D(16)=>
      FILTER(16), D(15)=>FILTER(15), D(14)=>FILTER(14), D(13)=>FILTER(13), 
      D(12)=>FILTER(12), D(11)=>FILTER(11), D(10)=>FILTER(10), D(9)=>
      FILTER(9), D(8)=>FILTER(8), D(7)=>FILTER(7), D(6)=>FILTER(6), D(5)=>
      FILTER(5), D(4)=>FILTER(4), D(3)=>FILTER(3), D(2)=>FILTER(2), D(1)=>
      FILTER(1), D(0)=>FILTER(0), CLK=>CLK, RST=>RST, EN=>filter2EN, Q(399)
      =>outFilter1(399), Q(398)=>outFilter1(398), Q(397)=>outFilter1(397), 
      Q(396)=>outFilter1(396), Q(395)=>outFilter1(395), Q(394)=>
      outFilter1(394), Q(393)=>outFilter1(393), Q(392)=>outFilter1(392), 
      Q(391)=>outFilter1(391), Q(390)=>outFilter1(390), Q(389)=>
      outFilter1(389), Q(388)=>outFilter1(388), Q(387)=>outFilter1(387), 
      Q(386)=>outFilter1(386), Q(385)=>outFilter1(385), Q(384)=>
      outFilter1(384), Q(383)=>outFilter1(383), Q(382)=>outFilter1(382), 
      Q(381)=>outFilter1(381), Q(380)=>outFilter1(380), Q(379)=>
      outFilter1(379), Q(378)=>outFilter1(378), Q(377)=>outFilter1(377), 
      Q(376)=>outFilter1(376), Q(375)=>outFilter1(375), Q(374)=>
      outFilter1(374), Q(373)=>outFilter1(373), Q(372)=>outFilter1(372), 
      Q(371)=>outFilter1(371), Q(370)=>outFilter1(370), Q(369)=>
      outFilter1(369), Q(368)=>outFilter1(368), Q(367)=>outFilter1(367), 
      Q(366)=>outFilter1(366), Q(365)=>outFilter1(365), Q(364)=>
      outFilter1(364), Q(363)=>outFilter1(363), Q(362)=>outFilter1(362), 
      Q(361)=>outFilter1(361), Q(360)=>outFilter1(360), Q(359)=>
      outFilter1(359), Q(358)=>outFilter1(358), Q(357)=>outFilter1(357), 
      Q(356)=>outFilter1(356), Q(355)=>outFilter1(355), Q(354)=>
      outFilter1(354), Q(353)=>outFilter1(353), Q(352)=>outFilter1(352), 
      Q(351)=>outFilter1(351), Q(350)=>outFilter1(350), Q(349)=>
      outFilter1(349), Q(348)=>outFilter1(348), Q(347)=>outFilter1(347), 
      Q(346)=>outFilter1(346), Q(345)=>outFilter1(345), Q(344)=>
      outFilter1(344), Q(343)=>outFilter1(343), Q(342)=>outFilter1(342), 
      Q(341)=>outFilter1(341), Q(340)=>outFilter1(340), Q(339)=>
      outFilter1(339), Q(338)=>outFilter1(338), Q(337)=>outFilter1(337), 
      Q(336)=>outFilter1(336), Q(335)=>outFilter1(335), Q(334)=>
      outFilter1(334), Q(333)=>outFilter1(333), Q(332)=>outFilter1(332), 
      Q(331)=>outFilter1(331), Q(330)=>outFilter1(330), Q(329)=>
      outFilter1(329), Q(328)=>outFilter1(328), Q(327)=>outFilter1(327), 
      Q(326)=>outFilter1(326), Q(325)=>outFilter1(325), Q(324)=>
      outFilter1(324), Q(323)=>outFilter1(323), Q(322)=>outFilter1(322), 
      Q(321)=>outFilter1(321), Q(320)=>outFilter1(320), Q(319)=>
      outFilter1(319), Q(318)=>outFilter1(318), Q(317)=>outFilter1(317), 
      Q(316)=>outFilter1(316), Q(315)=>outFilter1(315), Q(314)=>
      outFilter1(314), Q(313)=>outFilter1(313), Q(312)=>outFilter1(312), 
      Q(311)=>outFilter1(311), Q(310)=>outFilter1(310), Q(309)=>
      outFilter1(309), Q(308)=>outFilter1(308), Q(307)=>outFilter1(307), 
      Q(306)=>outFilter1(306), Q(305)=>outFilter1(305), Q(304)=>
      outFilter1(304), Q(303)=>outFilter1(303), Q(302)=>outFilter1(302), 
      Q(301)=>outFilter1(301), Q(300)=>outFilter1(300), Q(299)=>
      outFilter1(299), Q(298)=>outFilter1(298), Q(297)=>outFilter1(297), 
      Q(296)=>outFilter1(296), Q(295)=>outFilter1(295), Q(294)=>
      outFilter1(294), Q(293)=>outFilter1(293), Q(292)=>outFilter1(292), 
      Q(291)=>outFilter1(291), Q(290)=>outFilter1(290), Q(289)=>
      outFilter1(289), Q(288)=>outFilter1(288), Q(287)=>outFilter1(287), 
      Q(286)=>outFilter1(286), Q(285)=>outFilter1(285), Q(284)=>
      outFilter1(284), Q(283)=>outFilter1(283), Q(282)=>outFilter1(282), 
      Q(281)=>outFilter1(281), Q(280)=>outFilter1(280), Q(279)=>
      outFilter1(279), Q(278)=>outFilter1(278), Q(277)=>outFilter1(277), 
      Q(276)=>outFilter1(276), Q(275)=>outFilter1(275), Q(274)=>
      outFilter1(274), Q(273)=>outFilter1(273), Q(272)=>outFilter1(272), 
      Q(271)=>outFilter1(271), Q(270)=>outFilter1(270), Q(269)=>
      outFilter1(269), Q(268)=>outFilter1(268), Q(267)=>outFilter1(267), 
      Q(266)=>outFilter1(266), Q(265)=>outFilter1(265), Q(264)=>
      outFilter1(264), Q(263)=>outFilter1(263), Q(262)=>outFilter1(262), 
      Q(261)=>outFilter1(261), Q(260)=>outFilter1(260), Q(259)=>
      outFilter1(259), Q(258)=>outFilter1(258), Q(257)=>outFilter1(257), 
      Q(256)=>outFilter1(256), Q(255)=>outFilter1(255), Q(254)=>
      outFilter1(254), Q(253)=>outFilter1(253), Q(252)=>outFilter1(252), 
      Q(251)=>outFilter1(251), Q(250)=>outFilter1(250), Q(249)=>
      outFilter1(249), Q(248)=>outFilter1(248), Q(247)=>outFilter1(247), 
      Q(246)=>outFilter1(246), Q(245)=>outFilter1(245), Q(244)=>
      outFilter1(244), Q(243)=>outFilter1(243), Q(242)=>outFilter1(242), 
      Q(241)=>outFilter1(241), Q(240)=>outFilter1(240), Q(239)=>
      outFilter1(239), Q(238)=>outFilter1(238), Q(237)=>outFilter1(237), 
      Q(236)=>outFilter1(236), Q(235)=>outFilter1(235), Q(234)=>
      outFilter1(234), Q(233)=>outFilter1(233), Q(232)=>outFilter1(232), 
      Q(231)=>outFilter1(231), Q(230)=>outFilter1(230), Q(229)=>
      outFilter1(229), Q(228)=>outFilter1(228), Q(227)=>outFilter1(227), 
      Q(226)=>outFilter1(226), Q(225)=>outFilter1(225), Q(224)=>
      outFilter1(224), Q(223)=>outFilter1(223), Q(222)=>outFilter1(222), 
      Q(221)=>outFilter1(221), Q(220)=>outFilter1(220), Q(219)=>
      outFilter1(219), Q(218)=>outFilter1(218), Q(217)=>outFilter1(217), 
      Q(216)=>outFilter1(216), Q(215)=>outFilter1(215), Q(214)=>
      outFilter1(214), Q(213)=>outFilter1(213), Q(212)=>outFilter1(212), 
      Q(211)=>outFilter1(211), Q(210)=>outFilter1(210), Q(209)=>
      outFilter1(209), Q(208)=>outFilter1(208), Q(207)=>outFilter1(207), 
      Q(206)=>outFilter1(206), Q(205)=>outFilter1(205), Q(204)=>
      outFilter1(204), Q(203)=>outFilter1(203), Q(202)=>outFilter1(202), 
      Q(201)=>outFilter1(201), Q(200)=>outFilter1(200), Q(199)=>
      outFilter1(199), Q(198)=>outFilter1(198), Q(197)=>outFilter1(197), 
      Q(196)=>outFilter1(196), Q(195)=>outFilter1(195), Q(194)=>
      outFilter1(194), Q(193)=>outFilter1(193), Q(192)=>outFilter1(192), 
      Q(191)=>outFilter1(191), Q(190)=>outFilter1(190), Q(189)=>
      outFilter1(189), Q(188)=>outFilter1(188), Q(187)=>outFilter1(187), 
      Q(186)=>outFilter1(186), Q(185)=>outFilter1(185), Q(184)=>
      outFilter1(184), Q(183)=>outFilter1(183), Q(182)=>outFilter1(182), 
      Q(181)=>outFilter1(181), Q(180)=>outFilter1(180), Q(179)=>
      outFilter1(179), Q(178)=>outFilter1(178), Q(177)=>outFilter1(177), 
      Q(176)=>outFilter1(176), Q(175)=>outFilter1(175), Q(174)=>
      outFilter1(174), Q(173)=>outFilter1(173), Q(172)=>outFilter1(172), 
      Q(171)=>outFilter1(171), Q(170)=>outFilter1(170), Q(169)=>
      outFilter1(169), Q(168)=>outFilter1(168), Q(167)=>outFilter1(167), 
      Q(166)=>outFilter1(166), Q(165)=>outFilter1(165), Q(164)=>
      outFilter1(164), Q(163)=>outFilter1(163), Q(162)=>outFilter1(162), 
      Q(161)=>outFilter1(161), Q(160)=>outFilter1(160), Q(159)=>
      outFilter1(159), Q(158)=>outFilter1(158), Q(157)=>outFilter1(157), 
      Q(156)=>outFilter1(156), Q(155)=>outFilter1(155), Q(154)=>
      outFilter1(154), Q(153)=>outFilter1(153), Q(152)=>outFilter1(152), 
      Q(151)=>outFilter1(151), Q(150)=>outFilter1(150), Q(149)=>
      outFilter1(149), Q(148)=>outFilter1(148), Q(147)=>outFilter1(147), 
      Q(146)=>outFilter1(146), Q(145)=>outFilter1(145), Q(144)=>
      outFilter1(144), Q(143)=>outFilter1(143), Q(142)=>outFilter1(142), 
      Q(141)=>outFilter1(141), Q(140)=>outFilter1(140), Q(139)=>
      outFilter1(139), Q(138)=>outFilter1(138), Q(137)=>outFilter1(137), 
      Q(136)=>outFilter1(136), Q(135)=>outFilter1(135), Q(134)=>
      outFilter1(134), Q(133)=>outFilter1(133), Q(132)=>outFilter1(132), 
      Q(131)=>outFilter1(131), Q(130)=>outFilter1(130), Q(129)=>
      outFilter1(129), Q(128)=>outFilter1(128), Q(127)=>outFilter1(127), 
      Q(126)=>outFilter1(126), Q(125)=>outFilter1(125), Q(124)=>
      outFilter1(124), Q(123)=>outFilter1(123), Q(122)=>outFilter1(122), 
      Q(121)=>outFilter1(121), Q(120)=>outFilter1(120), Q(119)=>
      outFilter1(119), Q(118)=>outFilter1(118), Q(117)=>outFilter1(117), 
      Q(116)=>outFilter1(116), Q(115)=>outFilter1(115), Q(114)=>
      outFilter1(114), Q(113)=>outFilter1(113), Q(112)=>outFilter1(112), 
      Q(111)=>outFilter1(111), Q(110)=>outFilter1(110), Q(109)=>
      outFilter1(109), Q(108)=>outFilter1(108), Q(107)=>outFilter1(107), 
      Q(106)=>outFilter1(106), Q(105)=>outFilter1(105), Q(104)=>
      outFilter1(104), Q(103)=>outFilter1(103), Q(102)=>outFilter1(102), 
      Q(101)=>outFilter1(101), Q(100)=>outFilter1(100), Q(99)=>
      outFilter1(99), Q(98)=>outFilter1(98), Q(97)=>outFilter1(97), Q(96)=>
      outFilter1(96), Q(95)=>outFilter1(95), Q(94)=>outFilter1(94), Q(93)=>
      outFilter1(93), Q(92)=>outFilter1(92), Q(91)=>outFilter1(91), Q(90)=>
      outFilter1(90), Q(89)=>outFilter1(89), Q(88)=>outFilter1(88), Q(87)=>
      outFilter1(87), Q(86)=>outFilter1(86), Q(85)=>outFilter1(85), Q(84)=>
      outFilter1(84), Q(83)=>outFilter1(83), Q(82)=>outFilter1(82), Q(81)=>
      outFilter1(81), Q(80)=>outFilter1(80), Q(79)=>outFilter1(79), Q(78)=>
      outFilter1(78), Q(77)=>outFilter1(77), Q(76)=>outFilter1(76), Q(75)=>
      outFilter1(75), Q(74)=>outFilter1(74), Q(73)=>outFilter1(73), Q(72)=>
      outFilter1(72), Q(71)=>outFilter1(71), Q(70)=>outFilter1(70), Q(69)=>
      outFilter1(69), Q(68)=>outFilter1(68), Q(67)=>outFilter1(67), Q(66)=>
      outFilter1(66), Q(65)=>outFilter1(65), Q(64)=>outFilter1(64), Q(63)=>
      outFilter1(63), Q(62)=>outFilter1(62), Q(61)=>outFilter1(61), Q(60)=>
      outFilter1(60), Q(59)=>outFilter1(59), Q(58)=>outFilter1(58), Q(57)=>
      outFilter1(57), Q(56)=>outFilter1(56), Q(55)=>outFilter1(55), Q(54)=>
      outFilter1(54), Q(53)=>outFilter1(53), Q(52)=>outFilter1(52), Q(51)=>
      outFilter1(51), Q(50)=>outFilter1(50), Q(49)=>outFilter1(49), Q(48)=>
      outFilter1(48), Q(47)=>outFilter1(47), Q(46)=>outFilter1(46), Q(45)=>
      outFilter1(45), Q(44)=>outFilter1(44), Q(43)=>outFilter1(43), Q(42)=>
      outFilter1(42), Q(41)=>outFilter1(41), Q(40)=>outFilter1(40), Q(39)=>
      outFilter1(39), Q(38)=>outFilter1(38), Q(37)=>outFilter1(37), Q(36)=>
      outFilter1(36), Q(35)=>outFilter1(35), Q(34)=>outFilter1(34), Q(33)=>
      outFilter1(33), Q(32)=>outFilter1(32), Q(31)=>outFilter1(31), Q(30)=>
      outFilter1(30), Q(29)=>outFilter1(29), Q(28)=>outFilter1(28), Q(27)=>
      outFilter1(27), Q(26)=>outFilter1(26), Q(25)=>outFilter1(25), Q(24)=>
      outFilter1(24), Q(23)=>outFilter1(23), Q(22)=>outFilter1(22), Q(21)=>
      outFilter1(21), Q(20)=>outFilter1(20), Q(19)=>outFilter1(19), Q(18)=>
      outFilter1(18), Q(17)=>outFilter1(17), Q(16)=>outFilter1(16), Q(15)=>
      outFilter1(15), Q(14)=>outFilter1(14), Q(13)=>outFilter1(13), Q(12)=>
      outFilter1(12), Q(11)=>outFilter1(11), Q(10)=>outFilter1(10), Q(9)=>
      outFilter1(9), Q(8)=>outFilter1(8), Q(7)=>outFilter1(7), Q(6)=>
      outFilter1(6), Q(5)=>outFilter1(5), Q(4)=>outFilter1(4), Q(3)=>
      outFilter1(3), Q(2)=>outFilter1(2), Q(1)=>outFilter1(1), Q(0)=>
      outFilter1(0));
   DDF0 : nBitRegister_1 port map ( D(0)=>NOT_IndicatorFilter_0, CLK=>DFFCLK, 
      RST=>IndRst, EN=>secOperand_3, Q(0)=>IndicatorFilter_0_EXMPLR);
   tsb0 : triStateBuffer_13 port map ( D(12)=>FilterAddress(12), D(11)=>
      FilterAddress(11), D(10)=>FilterAddress(10), D(9)=>FilterAddress(9), 
      D(8)=>FilterAddress(8), D(7)=>FilterAddress(7), D(6)=>FilterAddress(6), 
      D(5)=>FilterAddress(5), D(4)=>FilterAddress(4), D(3)=>FilterAddress(3), 
      D(2)=>FilterAddress(2), D(1)=>FilterAddress(1), D(0)=>FilterAddress(0), 
      EN=>tristateAddEn, F(12)=>DMAAddress(12), F(11)=>DMAAddress(11), F(10)
      =>DMAAddress(10), F(9)=>DMAAddress(9), F(8)=>DMAAddress(8), F(7)=>
      DMAAddress(7), F(6)=>DMAAddress(6), F(5)=>DMAAddress(5), F(4)=>
      DMAAddress(4), F(3)=>DMAAddress(3), F(2)=>DMAAddress(2), F(1)=>
      DMAAddress(1), F(0)=>DMAAddress(0));
   adder0 : my_nadder_13 port map ( a(12)=>FilterAddress(12), a(11)=>
      FilterAddress(11), a(10)=>FilterAddress(10), a(9)=>FilterAddress(9), 
      a(8)=>FilterAddress(8), a(7)=>FilterAddress(7), a(6)=>FilterAddress(6), 
      a(5)=>FilterAddress(5), a(4)=>FilterAddress(4), a(3)=>FilterAddress(3), 
      a(2)=>FilterAddress(2), a(1)=>FilterAddress(1), a(0)=>FilterAddress(0), 
      b(12)=>secOperand_12, b(11)=>secOperand_12, b(10)=>secOperand_12, b(9)
      =>secOperand_12, b(8)=>secOperand_12, b(7)=>secOperand_12, b(6)=>
      secOperand_12, b(5)=>secOperand_12, b(4)=>msbNoOfFilters, b(3)=>
      secOperand_3, b(2)=>secOperand_12, b(1)=>secOperand_12, b(0)=>
      secOperand_3, cin=>secOperand_12, s(12)=>newAddress_12, s(11)=>
      newAddress_11, s(10)=>newAddress_10, s(9)=>newAddress_9, s(8)=>
      newAddress_8, s(7)=>newAddress_7, s(6)=>newAddress_6, s(5)=>
      newAddress_5, s(4)=>newAddress_4, s(3)=>newAddress_3, s(2)=>
      newAddress_2, s(1)=>newAddress_1, s(0)=>newAddress_0, cout=>DANGLING(3
      ));
   tsb2 : triStateBuffer_13 port map ( D(12)=>newAddress_12, D(11)=>
      newAddress_11, D(10)=>newAddress_10, D(9)=>newAddress_9, D(8)=>
      newAddress_8, D(7)=>newAddress_7, D(6)=>newAddress_6, D(5)=>
      newAddress_5, D(4)=>newAddress_4, D(3)=>newAddress_3, D(2)=>
      newAddress_2, D(1)=>newAddress_1, D(0)=>newAddress_0, EN=>
      tristateAddEn, F(12)=>UpdatedAddress(12), F(11)=>UpdatedAddress(11), 
      F(10)=>UpdatedAddress(10), F(9)=>UpdatedAddress(9), F(8)=>
      UpdatedAddress(8), F(7)=>UpdatedAddress(7), F(6)=>UpdatedAddress(6), 
      F(5)=>UpdatedAddress(5), F(4)=>UpdatedAddress(4), F(3)=>
      UpdatedAddress(3), F(2)=>UpdatedAddress(2), F(1)=>UpdatedAddress(1), 
      F(0)=>UpdatedAddress(0));
   ix1459 : inv01 port map ( Y=>NOT_IndicatorFilter_0, A=>
      IndicatorFilter_0_EXMPLR);
   ix1418 : fake_vcc port map ( Y=>secOperand_3);
   ix1416 : fake_gnd port map ( Y=>secOperand_12);
   ix5 : or02 port map ( Y=>tristateAddEn, A0=>nx2, A1=>current_state(5));
   ix3 : nor02ii port map ( Y=>nx2, A0=>IndicatorFilter_0_EXMPLR, A1=>
      current_state(7));
   ix101 : ao21 port map ( Y=>IndRst, A0=>current_state(10), A1=>nx96, B0=>
      RST);
   ix97 : nand03 port map ( Y=>nx96, A0=>nx1466, A1=>lastDepthOut_EXMPLR, A2
      =>donttrust_EXMPLR);
   ix1467 : or02 port map ( Y=>nx1466, A0=>LastFilterIND_EXMPLR, A1=>nx1477
   );
   ix77 : and04 port map ( Y=>LastFilterIND_EXMPLR, A0=>nx1469, A1=>nx1471, 
      A2=>nx1473, A3=>nx1475);
   ix1470 : xnor2 port map ( Y=>nx1469, A0=>FilterMinus_0, A1=>
      FilterCounter(0));
   ix1472 : xnor2 port map ( Y=>nx1471, A0=>FilterMinus_1, A1=>
      FilterCounter(1));
   ix1474 : xnor2 port map ( Y=>nx1473, A0=>FilterMinus_2, A1=>
      FilterCounter(2));
   ix1476 : xnor2 port map ( Y=>nx1475, A0=>FilterMinus_3, A1=>
      FilterCounter(3));
   ix1478 : nor04 port map ( Y=>nx1477, A0=>LayerInfo(1), A1=>LayerInfo(2), 
      A2=>LayerInfo(3), A3=>nx1479);
   ix1480 : inv01 port map ( Y=>nx1479, A=>LayerInfo(0));
   ix55 : and04 port map ( Y=>lastDepthOut_EXMPLR, A0=>nx1482, A1=>nx1484, 
      A2=>nx1486, A3=>nx1488);
   ix1483 : xnor2 port map ( Y=>nx1482, A0=>depthcounter(0), A1=>
      depthminus_0);
   ix1485 : xnor2 port map ( Y=>nx1484, A0=>depthcounter(1), A1=>
      depthminus_1);
   ix1487 : xnor2 port map ( Y=>nx1486, A0=>depthcounter(2), A1=>
      depthminus_2);
   ix1489 : xnor2 port map ( Y=>nx1488, A0=>depthcounter(3), A1=>
      depthminus_3);
   ix33 : nor03_2x port map ( Y=>donttrust_EXMPLR, A0=>nx1491, A1=>nx22, A2
      =>nx24);
   ix1492 : nand03 port map ( Y=>nx1491, A0=>nx1493, A1=>nx1495, A2=>nx1497
   );
   ix1494 : xnor2 port map ( Y=>nx1493, A0=>Heightminus_1, A1=>
      Heightcounter(1));
   ix1496 : xnor2 port map ( Y=>nx1495, A0=>Heightminus_4, A1=>
      Heightcounter(4));
   ix1498 : xnor2 port map ( Y=>nx1497, A0=>Heightminus_0, A1=>
      Heightcounter(0));
   ix23 : xor2 port map ( Y=>nx22, A0=>Heightminus_2, A1=>Heightcounter(2));
   ix25 : xor2 port map ( Y=>nx24, A0=>Heightminus_3, A1=>Heightcounter(3));
   ix123 : and02 port map ( Y=>filter2EN, A0=>ACKF, A1=>nx120);
   ix121 : mux21_ni port map ( Y=>nx120, A0=>nx2, A1=>current_state(5), S0=>
      QImgStat);
   ix133 : and02 port map ( Y=>filter1EN, A0=>ACKF, A1=>nx130);
   ix131 : mux21_ni port map ( Y=>nx130, A0=>current_state(5), A1=>nx2, S0=>
      QImgStat);
   reg_DFFCLK_dup_0 : dffr port map ( Q=>DFFCLK, QB=>OPEN, D=>secOperand_3, 
      CLK=>CLK, R=>nx108);
   ix109 : nand02 port map ( Y=>nx108, A0=>ACKF, A1=>current_state(7));
end DATA_FLOW ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity my_nadder_16 is
   port (
      a : IN std_logic_vector (15 DOWNTO 0) ;
      b : IN std_logic_vector (15 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (15 DOWNTO 0) ;
      cout : OUT std_logic) ;
end my_nadder_16 ;

architecture a_my_nadder of my_nadder_16 is
   component my_adder
      port (
         a : IN std_logic ;
         b : IN std_logic ;
         cin : IN std_logic ;
         s : OUT std_logic ;
         cout : OUT std_logic) ;
   end component ;
   signal temp_14, temp_13, temp_12, temp_11, temp_10, temp_9, temp_8, 
      temp_7, temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0: 
   std_logic ;

begin
   f0 : my_adder port map ( a=>a(0), b=>b(0), cin=>cin, s=>s(0), cout=>
      temp_0);
   loop1_1_fx : my_adder port map ( a=>a(1), b=>b(1), cin=>temp_0, s=>s(1), 
      cout=>temp_1);
   loop1_2_fx : my_adder port map ( a=>a(2), b=>b(2), cin=>temp_1, s=>s(2), 
      cout=>temp_2);
   loop1_3_fx : my_adder port map ( a=>a(3), b=>b(3), cin=>temp_2, s=>s(3), 
      cout=>temp_3);
   loop1_4_fx : my_adder port map ( a=>a(4), b=>b(4), cin=>temp_3, s=>s(4), 
      cout=>temp_4);
   loop1_5_fx : my_adder port map ( a=>a(5), b=>b(5), cin=>temp_4, s=>s(5), 
      cout=>temp_5);
   loop1_6_fx : my_adder port map ( a=>a(6), b=>b(6), cin=>temp_5, s=>s(6), 
      cout=>temp_6);
   loop1_7_fx : my_adder port map ( a=>a(7), b=>b(7), cin=>temp_6, s=>s(7), 
      cout=>temp_7);
   loop1_8_fx : my_adder port map ( a=>a(8), b=>b(8), cin=>temp_7, s=>s(8), 
      cout=>temp_8);
   loop1_9_fx : my_adder port map ( a=>a(9), b=>b(9), cin=>temp_8, s=>s(9), 
      cout=>temp_9);
   loop1_10_fx : my_adder port map ( a=>a(10), b=>b(10), cin=>temp_9, s=>
      s(10), cout=>temp_10);
   loop1_11_fx : my_adder port map ( a=>a(11), b=>b(11), cin=>temp_10, s=>
      s(11), cout=>temp_11);
   loop1_12_fx : my_adder port map ( a=>a(12), b=>b(12), cin=>temp_11, s=>
      s(12), cout=>temp_12);
   loop1_13_fx : my_adder port map ( a=>a(13), b=>b(13), cin=>temp_12, s=>
      s(13), cout=>temp_13);
   loop1_14_fx : my_adder port map ( a=>a(14), b=>b(14), cin=>temp_13, s=>
      s(14), cout=>temp_14);
   loop1_15_fx : my_adder port map ( a=>a(15), b=>b(15), cin=>temp_14, s=>
      s(15), cout=>cout);
end a_my_nadder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity my_nadder_3 is
   port (
      a : IN std_logic_vector (2 DOWNTO 0) ;
      b : IN std_logic_vector (2 DOWNTO 0) ;
      cin : IN std_logic ;
      s : OUT std_logic_vector (2 DOWNTO 0) ;
      cout : OUT std_logic) ;
end my_nadder_3 ;

architecture a_my_nadder of my_nadder_3 is
   component my_adder
      port (
         a : IN std_logic ;
         b : IN std_logic ;
         cin : IN std_logic ;
         s : OUT std_logic ;
         cout : OUT std_logic) ;
   end component ;
   signal temp_1, temp_0: std_logic ;

begin
   f0 : my_adder port map ( a=>a(0), b=>b(0), cin=>cin, s=>s(0), cout=>
      temp_0);
   loop1_1_fx : my_adder port map ( a=>a(1), b=>b(1), cin=>temp_0, s=>s(1), 
      cout=>temp_1);
   loop1_2_fx : my_adder port map ( a=>a(2), b=>b(2), cin=>temp_1, s=>s(2), 
      cout=>cout);
end a_my_nadder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Counter_3 is
   port (
      enable : IN std_logic ;
      reset : IN std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      output : OUT std_logic_vector (2 DOWNTO 0) ;
      input : IN std_logic_vector (2 DOWNTO 0)) ;
end Counter_3 ;

architecture CounterImplementation of Counter_3 is
   component my_nadder_3
      port (
         a : IN std_logic_vector (2 DOWNTO 0) ;
         b : IN std_logic_vector (2 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (2 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal output_2_EXMPLR, output_1_EXMPLR, output_0_EXMPLR, addResult_2, 
      addResult_1, addResult_0, one_0, one_2, nx40, NOT_clk, nx8, nx12, nx34, 
      nx20, nx24, nx28, nx33, nx37, nx114, nx124, nx134, nx143: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   output(2) <= output_2_EXMPLR ;
   output(1) <= output_1_EXMPLR ;
   output(0) <= output_0_EXMPLR ;
   A1 : my_nadder_3 port map ( a(2)=>output_2_EXMPLR, a(1)=>output_1_EXMPLR, 
      a(0)=>output_0_EXMPLR, b(2)=>one_2, b(1)=>one_2, b(0)=>one_0, cin=>
      one_2, s(2)=>addResult_2, s(1)=>addResult_1, s(0)=>addResult_0, cout=>
      DANGLING(0));
   ix94 : fake_gnd port map ( Y=>one_2);
   ix92 : fake_vcc port map ( Y=>one_0);
   reg_toOutput_0_dup_1 : dffsr_ni port map ( Q=>output_0_EXMPLR, QB=>OPEN, 
      D=>nx114, CLK=>clk, S=>nx8, R=>nx12);
   ix115 : mux21_ni port map ( Y=>nx114, A0=>output_0_EXMPLR, A1=>
      addResult_0, S0=>enable);
   ix9 : nor02ii port map ( Y=>nx8, A0=>nx143, A1=>nx40);
   ix144 : nor02_2x port map ( Y=>nx143, A0=>reset, A1=>load);
   ix41 : dffr port map ( Q=>nx40, QB=>OPEN, D=>input(0), CLK=>NOT_clk, R=>
      reset);
   ix147 : inv01 port map ( Y=>NOT_clk, A=>clk);
   ix13 : nor02_2x port map ( Y=>nx12, A0=>nx40, A1=>nx143);
   reg_toOutput_1_dup_1 : dffsr_ni port map ( Q=>output_1_EXMPLR, QB=>OPEN, 
      D=>nx124, CLK=>clk, S=>nx20, R=>nx24);
   ix125 : mux21_ni port map ( Y=>nx124, A0=>output_1_EXMPLR, A1=>
      addResult_1, S0=>enable);
   ix21 : nor02ii port map ( Y=>nx20, A0=>nx143, A1=>nx34);
   ix35 : dffr port map ( Q=>nx34, QB=>OPEN, D=>input(1), CLK=>NOT_clk, R=>
      reset);
   ix25 : nor02_2x port map ( Y=>nx24, A0=>nx34, A1=>nx143);
   reg_toOutput_2_dup_1 : dffsr_ni port map ( Q=>output_2_EXMPLR, QB=>OPEN, 
      D=>nx134, CLK=>clk, S=>nx33, R=>nx37);
   ix135 : mux21_ni port map ( Y=>nx134, A0=>output_2_EXMPLR, A1=>
      addResult_2, S0=>enable);
   ix34 : nor02ii port map ( Y=>nx33, A0=>nx143, A1=>nx28);
   ix29 : dffr port map ( Q=>nx28, QB=>OPEN, D=>input(2), CLK=>NOT_clk, R=>
      reset);
   ix38 : nor02_2x port map ( Y=>nx37, A0=>nx28, A1=>nx143);
end CounterImplementation ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Decoder is
   port (
      input : IN std_logic_vector (2 DOWNTO 0) ;
      output : OUT std_logic_vector (5 DOWNTO 0)) ;
end Decoder ;

architecture dec of Decoder is
   signal nx4, nx14, nx28, nx42, nx54, nx68, nx80, nx145, nx149, nx155, 
      nx164, nx166: std_logic ;

begin
   lat_output_0 : latch port map ( Q=>output(0), D=>nx14, CLK=>nx4);
   ix15 : nor03_2x port map ( Y=>nx14, A0=>nx164, A1=>nx166, A2=>input(0));
   ix5 : nand02 port map ( Y=>nx4, A0=>nx164, A1=>nx166);
   lat_output_1 : latch port map ( Q=>output(1), D=>nx28, CLK=>nx4);
   ix29 : nor03_2x port map ( Y=>nx28, A0=>nx164, A1=>nx166, A2=>nx145);
   ix146 : inv01 port map ( Y=>nx145, A=>input(0));
   lat_output_2 : latch port map ( Q=>output(2), D=>nx42, CLK=>nx4);
   ix43 : nor03_2x port map ( Y=>nx42, A0=>nx164, A1=>nx149, A2=>input(0));
   ix150 : inv01 port map ( Y=>nx149, A=>input(1));
   lat_output_3 : latch port map ( Q=>output(3), D=>nx54, CLK=>nx4);
   ix55 : nor03_2x port map ( Y=>nx54, A0=>nx164, A1=>nx149, A2=>nx145);
   lat_output_4 : latch port map ( Q=>output(4), D=>nx68, CLK=>nx4);
   ix69 : nor03_2x port map ( Y=>nx68, A0=>nx155, A1=>nx166, A2=>input(0));
   ix156 : inv01 port map ( Y=>nx155, A=>input(2));
   lat_output_5 : latch port map ( Q=>output(5), D=>nx80, CLK=>nx4);
   ix81 : nor03_2x port map ( Y=>nx80, A0=>nx155, A1=>nx166, A2=>nx145);
   ix163 : inv02 port map ( Y=>nx164, A=>nx155);
   ix165 : inv02 port map ( Y=>nx166, A=>nx149);
end dec ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity triStateBuffer_6 is
   port (
      D : IN std_logic_vector (5 DOWNTO 0) ;
      EN : IN std_logic ;
      F : OUT std_logic_vector (5 DOWNTO 0)) ;
end triStateBuffer_6 ;

architecture triBuffer of triStateBuffer_6 is
   signal nx115, nx118, nx121, nx124, nx127, nx130: std_logic ;

begin
   tri_F_0 : tri01 port map ( Y=>F(0), A=>nx115, E=>EN);
   ix116 : inv01 port map ( Y=>nx115, A=>D(0));
   tri_F_1 : tri01 port map ( Y=>F(1), A=>nx118, E=>EN);
   ix119 : inv01 port map ( Y=>nx118, A=>D(1));
   tri_F_2 : tri01 port map ( Y=>F(2), A=>nx121, E=>EN);
   ix122 : inv01 port map ( Y=>nx121, A=>D(2));
   tri_F_3 : tri01 port map ( Y=>F(3), A=>nx124, E=>EN);
   ix125 : inv01 port map ( Y=>nx124, A=>D(3));
   tri_F_4 : tri01 port map ( Y=>F(4), A=>nx127, E=>EN);
   ix128 : inv01 port map ( Y=>nx127, A=>D(4));
   tri_F_5 : tri01 port map ( Y=>F(5), A=>nx130, E=>EN);
   ix131 : inv01 port map ( Y=>nx130, A=>D(5));
end triBuffer ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity ReadImage is
   port (
      WI : IN std_logic ;
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      ACK : IN std_logic ;
      ImgAddress : IN std_logic_vector (12 DOWNTO 0) ;
      ImgWidth : IN std_logic_vector (15 DOWNTO 0) ;
      DATA : IN std_logic_vector (447 DOWNTO 0) ;
      OutputImg0 : OUT std_logic_vector (447 DOWNTO 0) ;
      OutputImg1 : OUT std_logic_vector (447 DOWNTO 0) ;
      OutputImg2 : OUT std_logic_vector (447 DOWNTO 0) ;
      OutputImg3 : OUT std_logic_vector (447 DOWNTO 0) ;
      OutputImg4 : OUT std_logic_vector (447 DOWNTO 0) ;
      OutputImg5 : OUT std_logic_vector (447 DOWNTO 0) ;
      ImgCounterOuput : OUT std_logic_vector (2 DOWNTO 0) ;
      ImgAddToDma : OUT std_logic_vector (12 DOWNTO 0) ;
      UpdatedAddress : OUT std_logic_vector (12 DOWNTO 0) ;
      ImgIndic : OUT std_logic_vector (0 DOWNTO 0) ;
      ImgEn : OUT std_logic_vector (5 DOWNTO 0) ;
      dontTrust : IN std_logic) ;
end ReadImage ;

architecture archRI of ReadImage is
   component my_nadder_16
      port (
         a : IN std_logic_vector (15 DOWNTO 0) ;
         b : IN std_logic_vector (15 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (15 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component nBitRegister_1
      port (
         D : IN std_logic_vector (0 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (0 DOWNTO 0)) ;
   end component ;
   component Counter_3
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (2 DOWNTO 0) ;
         input : IN std_logic_vector (2 DOWNTO 0)) ;
   end component ;
   component Decoder
      port (
         input : IN std_logic_vector (2 DOWNTO 0) ;
         output : OUT std_logic_vector (5 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_6
      port (
         D : IN std_logic_vector (5 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (5 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component nBitRegister_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal OutputImg0_447_EXMPLR, OutputImg0_446_EXMPLR, 
      OutputImg0_445_EXMPLR, OutputImg0_444_EXMPLR, OutputImg0_443_EXMPLR, 
      OutputImg0_442_EXMPLR, OutputImg0_441_EXMPLR, OutputImg0_440_EXMPLR, 
      OutputImg0_439_EXMPLR, OutputImg0_438_EXMPLR, OutputImg0_437_EXMPLR, 
      OutputImg0_436_EXMPLR, OutputImg0_435_EXMPLR, OutputImg0_434_EXMPLR, 
      OutputImg0_433_EXMPLR, OutputImg0_432_EXMPLR, OutputImg0_431_EXMPLR, 
      OutputImg0_430_EXMPLR, OutputImg0_429_EXMPLR, OutputImg0_428_EXMPLR, 
      OutputImg0_427_EXMPLR, OutputImg0_426_EXMPLR, OutputImg0_425_EXMPLR, 
      OutputImg0_424_EXMPLR, OutputImg0_423_EXMPLR, OutputImg0_422_EXMPLR, 
      OutputImg0_421_EXMPLR, OutputImg0_420_EXMPLR, OutputImg0_419_EXMPLR, 
      OutputImg0_418_EXMPLR, OutputImg0_417_EXMPLR, OutputImg0_416_EXMPLR, 
      OutputImg0_415_EXMPLR, OutputImg0_414_EXMPLR, OutputImg0_413_EXMPLR, 
      OutputImg0_412_EXMPLR, OutputImg0_411_EXMPLR, OutputImg0_410_EXMPLR, 
      OutputImg0_409_EXMPLR, OutputImg0_408_EXMPLR, OutputImg0_407_EXMPLR, 
      OutputImg0_406_EXMPLR, OutputImg0_405_EXMPLR, OutputImg0_404_EXMPLR, 
      OutputImg0_403_EXMPLR, OutputImg0_402_EXMPLR, OutputImg0_401_EXMPLR, 
      OutputImg0_400_EXMPLR, OutputImg0_399_EXMPLR, OutputImg0_398_EXMPLR, 
      OutputImg0_397_EXMPLR, OutputImg0_396_EXMPLR, OutputImg0_395_EXMPLR, 
      OutputImg0_394_EXMPLR, OutputImg0_393_EXMPLR, OutputImg0_392_EXMPLR, 
      OutputImg0_391_EXMPLR, OutputImg0_390_EXMPLR, OutputImg0_389_EXMPLR, 
      OutputImg0_388_EXMPLR, OutputImg0_387_EXMPLR, OutputImg0_386_EXMPLR, 
      OutputImg0_385_EXMPLR, OutputImg0_384_EXMPLR, OutputImg0_383_EXMPLR, 
      OutputImg0_382_EXMPLR, OutputImg0_381_EXMPLR, OutputImg0_380_EXMPLR, 
      OutputImg0_379_EXMPLR, OutputImg0_378_EXMPLR, OutputImg0_377_EXMPLR, 
      OutputImg0_376_EXMPLR, OutputImg0_375_EXMPLR, OutputImg0_374_EXMPLR, 
      OutputImg0_373_EXMPLR, OutputImg0_372_EXMPLR, OutputImg0_371_EXMPLR, 
      OutputImg0_370_EXMPLR, OutputImg0_369_EXMPLR, OutputImg0_368_EXMPLR, 
      OutputImg0_367_EXMPLR, OutputImg0_366_EXMPLR, OutputImg0_365_EXMPLR, 
      OutputImg0_364_EXMPLR, OutputImg0_363_EXMPLR, OutputImg0_362_EXMPLR, 
      OutputImg0_361_EXMPLR, OutputImg0_360_EXMPLR, OutputImg0_359_EXMPLR, 
      OutputImg0_358_EXMPLR, OutputImg0_357_EXMPLR, OutputImg0_356_EXMPLR, 
      OutputImg0_355_EXMPLR, OutputImg0_354_EXMPLR, OutputImg0_353_EXMPLR, 
      OutputImg0_352_EXMPLR, OutputImg0_351_EXMPLR, OutputImg0_350_EXMPLR, 
      OutputImg0_349_EXMPLR, OutputImg0_348_EXMPLR, OutputImg0_347_EXMPLR, 
      OutputImg0_346_EXMPLR, OutputImg0_345_EXMPLR, OutputImg0_344_EXMPLR, 
      OutputImg0_343_EXMPLR, OutputImg0_342_EXMPLR, OutputImg0_341_EXMPLR, 
      OutputImg0_340_EXMPLR, OutputImg0_339_EXMPLR, OutputImg0_338_EXMPLR, 
      OutputImg0_337_EXMPLR, OutputImg0_336_EXMPLR, OutputImg0_335_EXMPLR, 
      OutputImg0_334_EXMPLR, OutputImg0_333_EXMPLR, OutputImg0_332_EXMPLR, 
      OutputImg0_331_EXMPLR, OutputImg0_330_EXMPLR, OutputImg0_329_EXMPLR, 
      OutputImg0_328_EXMPLR, OutputImg0_327_EXMPLR, OutputImg0_326_EXMPLR, 
      OutputImg0_325_EXMPLR, OutputImg0_324_EXMPLR, OutputImg0_323_EXMPLR, 
      OutputImg0_322_EXMPLR, OutputImg0_321_EXMPLR, OutputImg0_320_EXMPLR, 
      OutputImg0_319_EXMPLR, OutputImg0_318_EXMPLR, OutputImg0_317_EXMPLR, 
      OutputImg0_316_EXMPLR, OutputImg0_315_EXMPLR, OutputImg0_314_EXMPLR, 
      OutputImg0_313_EXMPLR, OutputImg0_312_EXMPLR, OutputImg0_311_EXMPLR, 
      OutputImg0_310_EXMPLR, OutputImg0_309_EXMPLR, OutputImg0_308_EXMPLR, 
      OutputImg0_307_EXMPLR, OutputImg0_306_EXMPLR, OutputImg0_305_EXMPLR, 
      OutputImg0_304_EXMPLR, OutputImg0_303_EXMPLR, OutputImg0_302_EXMPLR, 
      OutputImg0_301_EXMPLR, OutputImg0_300_EXMPLR, OutputImg0_299_EXMPLR, 
      OutputImg0_298_EXMPLR, OutputImg0_297_EXMPLR, OutputImg0_296_EXMPLR, 
      OutputImg0_295_EXMPLR, OutputImg0_294_EXMPLR, OutputImg0_293_EXMPLR, 
      OutputImg0_292_EXMPLR, OutputImg0_291_EXMPLR, OutputImg0_290_EXMPLR, 
      OutputImg0_289_EXMPLR, OutputImg0_288_EXMPLR, OutputImg0_287_EXMPLR, 
      OutputImg0_286_EXMPLR, OutputImg0_285_EXMPLR, OutputImg0_284_EXMPLR, 
      OutputImg0_283_EXMPLR, OutputImg0_282_EXMPLR, OutputImg0_281_EXMPLR, 
      OutputImg0_280_EXMPLR, OutputImg0_279_EXMPLR, OutputImg0_278_EXMPLR, 
      OutputImg0_277_EXMPLR, OutputImg0_276_EXMPLR, OutputImg0_275_EXMPLR, 
      OutputImg0_274_EXMPLR, OutputImg0_273_EXMPLR, OutputImg0_272_EXMPLR, 
      OutputImg0_271_EXMPLR, OutputImg0_270_EXMPLR, OutputImg0_269_EXMPLR, 
      OutputImg0_268_EXMPLR, OutputImg0_267_EXMPLR, OutputImg0_266_EXMPLR, 
      OutputImg0_265_EXMPLR, OutputImg0_264_EXMPLR, OutputImg0_263_EXMPLR, 
      OutputImg0_262_EXMPLR, OutputImg0_261_EXMPLR, OutputImg0_260_EXMPLR, 
      OutputImg0_259_EXMPLR, OutputImg0_258_EXMPLR, OutputImg0_257_EXMPLR, 
      OutputImg0_256_EXMPLR, OutputImg0_255_EXMPLR, OutputImg0_254_EXMPLR, 
      OutputImg0_253_EXMPLR, OutputImg0_252_EXMPLR, OutputImg0_251_EXMPLR, 
      OutputImg0_250_EXMPLR, OutputImg0_249_EXMPLR, OutputImg0_248_EXMPLR, 
      OutputImg0_247_EXMPLR, OutputImg0_246_EXMPLR, OutputImg0_245_EXMPLR, 
      OutputImg0_244_EXMPLR, OutputImg0_243_EXMPLR, OutputImg0_242_EXMPLR, 
      OutputImg0_241_EXMPLR, OutputImg0_240_EXMPLR, OutputImg0_239_EXMPLR, 
      OutputImg0_238_EXMPLR, OutputImg0_237_EXMPLR, OutputImg0_236_EXMPLR, 
      OutputImg0_235_EXMPLR, OutputImg0_234_EXMPLR, OutputImg0_233_EXMPLR, 
      OutputImg0_232_EXMPLR, OutputImg0_231_EXMPLR, OutputImg0_230_EXMPLR, 
      OutputImg0_229_EXMPLR, OutputImg0_228_EXMPLR, OutputImg0_227_EXMPLR, 
      OutputImg0_226_EXMPLR, OutputImg0_225_EXMPLR, OutputImg0_224_EXMPLR, 
      OutputImg0_223_EXMPLR, OutputImg0_222_EXMPLR, OutputImg0_221_EXMPLR, 
      OutputImg0_220_EXMPLR, OutputImg0_219_EXMPLR, OutputImg0_218_EXMPLR, 
      OutputImg0_217_EXMPLR, OutputImg0_216_EXMPLR, OutputImg0_215_EXMPLR, 
      OutputImg0_214_EXMPLR, OutputImg0_213_EXMPLR, OutputImg0_212_EXMPLR, 
      OutputImg0_211_EXMPLR, OutputImg0_210_EXMPLR, OutputImg0_209_EXMPLR, 
      OutputImg0_208_EXMPLR, OutputImg0_207_EXMPLR, OutputImg0_206_EXMPLR, 
      OutputImg0_205_EXMPLR, OutputImg0_204_EXMPLR, OutputImg0_203_EXMPLR, 
      OutputImg0_202_EXMPLR, OutputImg0_201_EXMPLR, OutputImg0_200_EXMPLR, 
      OutputImg0_199_EXMPLR, OutputImg0_198_EXMPLR, OutputImg0_197_EXMPLR, 
      OutputImg0_196_EXMPLR, OutputImg0_195_EXMPLR, OutputImg0_194_EXMPLR, 
      OutputImg0_193_EXMPLR, OutputImg0_192_EXMPLR, OutputImg0_191_EXMPLR, 
      OutputImg0_190_EXMPLR, OutputImg0_189_EXMPLR, OutputImg0_188_EXMPLR, 
      OutputImg0_187_EXMPLR, OutputImg0_186_EXMPLR, OutputImg0_185_EXMPLR, 
      OutputImg0_184_EXMPLR, OutputImg0_183_EXMPLR, OutputImg0_182_EXMPLR, 
      OutputImg0_181_EXMPLR, OutputImg0_180_EXMPLR, OutputImg0_179_EXMPLR, 
      OutputImg0_178_EXMPLR, OutputImg0_177_EXMPLR, OutputImg0_176_EXMPLR, 
      OutputImg0_175_EXMPLR, OutputImg0_174_EXMPLR, OutputImg0_173_EXMPLR, 
      OutputImg0_172_EXMPLR, OutputImg0_171_EXMPLR, OutputImg0_170_EXMPLR, 
      OutputImg0_169_EXMPLR, OutputImg0_168_EXMPLR, OutputImg0_167_EXMPLR, 
      OutputImg0_166_EXMPLR, OutputImg0_165_EXMPLR, OutputImg0_164_EXMPLR, 
      OutputImg0_163_EXMPLR, OutputImg0_162_EXMPLR, OutputImg0_161_EXMPLR, 
      OutputImg0_160_EXMPLR, OutputImg0_159_EXMPLR, OutputImg0_158_EXMPLR, 
      OutputImg0_157_EXMPLR, OutputImg0_156_EXMPLR, OutputImg0_155_EXMPLR, 
      OutputImg0_154_EXMPLR, OutputImg0_153_EXMPLR, OutputImg0_152_EXMPLR, 
      OutputImg0_151_EXMPLR, OutputImg0_150_EXMPLR, OutputImg0_149_EXMPLR, 
      OutputImg0_148_EXMPLR, OutputImg0_147_EXMPLR, OutputImg0_146_EXMPLR, 
      OutputImg0_145_EXMPLR, OutputImg0_144_EXMPLR, OutputImg0_143_EXMPLR, 
      OutputImg0_142_EXMPLR, OutputImg0_141_EXMPLR, OutputImg0_140_EXMPLR, 
      OutputImg0_139_EXMPLR, OutputImg0_138_EXMPLR, OutputImg0_137_EXMPLR, 
      OutputImg0_136_EXMPLR, OutputImg0_135_EXMPLR, OutputImg0_134_EXMPLR, 
      OutputImg0_133_EXMPLR, OutputImg0_132_EXMPLR, OutputImg0_131_EXMPLR, 
      OutputImg0_130_EXMPLR, OutputImg0_129_EXMPLR, OutputImg0_128_EXMPLR, 
      OutputImg0_127_EXMPLR, OutputImg0_126_EXMPLR, OutputImg0_125_EXMPLR, 
      OutputImg0_124_EXMPLR, OutputImg0_123_EXMPLR, OutputImg0_122_EXMPLR, 
      OutputImg0_121_EXMPLR, OutputImg0_120_EXMPLR, OutputImg0_119_EXMPLR, 
      OutputImg0_118_EXMPLR, OutputImg0_117_EXMPLR, OutputImg0_116_EXMPLR, 
      OutputImg0_115_EXMPLR, OutputImg0_114_EXMPLR, OutputImg0_113_EXMPLR, 
      OutputImg0_112_EXMPLR, OutputImg0_111_EXMPLR, OutputImg0_110_EXMPLR, 
      OutputImg0_109_EXMPLR, OutputImg0_108_EXMPLR, OutputImg0_107_EXMPLR, 
      OutputImg0_106_EXMPLR, OutputImg0_105_EXMPLR, OutputImg0_104_EXMPLR, 
      OutputImg0_103_EXMPLR, OutputImg0_102_EXMPLR, OutputImg0_101_EXMPLR, 
      OutputImg0_100_EXMPLR, OutputImg0_99_EXMPLR, OutputImg0_98_EXMPLR, 
      OutputImg0_97_EXMPLR, OutputImg0_96_EXMPLR, OutputImg0_95_EXMPLR, 
      OutputImg0_94_EXMPLR, OutputImg0_93_EXMPLR, OutputImg0_92_EXMPLR, 
      OutputImg0_91_EXMPLR, OutputImg0_90_EXMPLR, OutputImg0_89_EXMPLR, 
      OutputImg0_88_EXMPLR, OutputImg0_87_EXMPLR, OutputImg0_86_EXMPLR, 
      OutputImg0_85_EXMPLR, OutputImg0_84_EXMPLR, OutputImg0_83_EXMPLR, 
      OutputImg0_82_EXMPLR, OutputImg0_81_EXMPLR, OutputImg0_80_EXMPLR, 
      OutputImg0_79_EXMPLR, OutputImg0_78_EXMPLR, OutputImg0_77_EXMPLR, 
      OutputImg0_76_EXMPLR, OutputImg0_75_EXMPLR, OutputImg0_74_EXMPLR, 
      OutputImg0_73_EXMPLR, OutputImg0_72_EXMPLR, OutputImg0_71_EXMPLR, 
      OutputImg0_70_EXMPLR, OutputImg0_69_EXMPLR, OutputImg0_68_EXMPLR, 
      OutputImg0_67_EXMPLR, OutputImg0_66_EXMPLR, OutputImg0_65_EXMPLR, 
      OutputImg0_64_EXMPLR, OutputImg0_63_EXMPLR, OutputImg0_62_EXMPLR, 
      OutputImg0_61_EXMPLR, OutputImg0_60_EXMPLR, OutputImg0_59_EXMPLR, 
      OutputImg0_58_EXMPLR, OutputImg0_57_EXMPLR, OutputImg0_56_EXMPLR, 
      OutputImg0_55_EXMPLR, OutputImg0_54_EXMPLR, OutputImg0_53_EXMPLR, 
      OutputImg0_52_EXMPLR, OutputImg0_51_EXMPLR, OutputImg0_50_EXMPLR, 
      OutputImg0_49_EXMPLR, OutputImg0_48_EXMPLR, OutputImg0_47_EXMPLR, 
      OutputImg0_46_EXMPLR, OutputImg0_45_EXMPLR, OutputImg0_44_EXMPLR, 
      OutputImg0_43_EXMPLR, OutputImg0_42_EXMPLR, OutputImg0_41_EXMPLR, 
      OutputImg0_40_EXMPLR, OutputImg0_39_EXMPLR, OutputImg0_38_EXMPLR, 
      OutputImg0_37_EXMPLR, OutputImg0_36_EXMPLR, OutputImg0_35_EXMPLR, 
      OutputImg0_34_EXMPLR, OutputImg0_33_EXMPLR, OutputImg0_32_EXMPLR, 
      OutputImg0_31_EXMPLR, OutputImg0_30_EXMPLR, OutputImg0_29_EXMPLR, 
      OutputImg0_28_EXMPLR, OutputImg0_27_EXMPLR, OutputImg0_26_EXMPLR, 
      OutputImg0_25_EXMPLR, OutputImg0_24_EXMPLR, OutputImg0_23_EXMPLR, 
      OutputImg0_22_EXMPLR, OutputImg0_21_EXMPLR, OutputImg0_20_EXMPLR, 
      OutputImg0_19_EXMPLR, OutputImg0_18_EXMPLR, OutputImg0_17_EXMPLR, 
      OutputImg0_16_EXMPLR, OutputImg0_15_EXMPLR, OutputImg0_14_EXMPLR, 
      OutputImg0_13_EXMPLR, OutputImg0_12_EXMPLR, OutputImg0_11_EXMPLR, 
      OutputImg0_10_EXMPLR, OutputImg0_9_EXMPLR, OutputImg0_8_EXMPLR, 
      OutputImg0_7_EXMPLR, OutputImg0_6_EXMPLR, OutputImg0_5_EXMPLR, 
      OutputImg0_4_EXMPLR, OutputImg0_3_EXMPLR, OutputImg0_2_EXMPLR, 
      OutputImg0_1_EXMPLR, OutputImg0_0_EXMPLR, OutputImg1_447_EXMPLR, 
      OutputImg1_446_EXMPLR, OutputImg1_445_EXMPLR, OutputImg1_444_EXMPLR, 
      OutputImg1_443_EXMPLR, OutputImg1_442_EXMPLR, OutputImg1_441_EXMPLR, 
      OutputImg1_440_EXMPLR, OutputImg1_439_EXMPLR, OutputImg1_438_EXMPLR, 
      OutputImg1_437_EXMPLR, OutputImg1_436_EXMPLR, OutputImg1_435_EXMPLR, 
      OutputImg1_434_EXMPLR, OutputImg1_433_EXMPLR, OutputImg1_432_EXMPLR, 
      OutputImg1_431_EXMPLR, OutputImg1_430_EXMPLR, OutputImg1_429_EXMPLR, 
      OutputImg1_428_EXMPLR, OutputImg1_427_EXMPLR, OutputImg1_426_EXMPLR, 
      OutputImg1_425_EXMPLR, OutputImg1_424_EXMPLR, OutputImg1_423_EXMPLR, 
      OutputImg1_422_EXMPLR, OutputImg1_421_EXMPLR, OutputImg1_420_EXMPLR, 
      OutputImg1_419_EXMPLR, OutputImg1_418_EXMPLR, OutputImg1_417_EXMPLR, 
      OutputImg1_416_EXMPLR, OutputImg1_415_EXMPLR, OutputImg1_414_EXMPLR, 
      OutputImg1_413_EXMPLR, OutputImg1_412_EXMPLR, OutputImg1_411_EXMPLR, 
      OutputImg1_410_EXMPLR, OutputImg1_409_EXMPLR, OutputImg1_408_EXMPLR, 
      OutputImg1_407_EXMPLR, OutputImg1_406_EXMPLR, OutputImg1_405_EXMPLR, 
      OutputImg1_404_EXMPLR, OutputImg1_403_EXMPLR, OutputImg1_402_EXMPLR, 
      OutputImg1_401_EXMPLR, OutputImg1_400_EXMPLR, OutputImg1_399_EXMPLR, 
      OutputImg1_398_EXMPLR, OutputImg1_397_EXMPLR, OutputImg1_396_EXMPLR, 
      OutputImg1_395_EXMPLR, OutputImg1_394_EXMPLR, OutputImg1_393_EXMPLR, 
      OutputImg1_392_EXMPLR, OutputImg1_391_EXMPLR, OutputImg1_390_EXMPLR, 
      OutputImg1_389_EXMPLR, OutputImg1_388_EXMPLR, OutputImg1_387_EXMPLR, 
      OutputImg1_386_EXMPLR, OutputImg1_385_EXMPLR, OutputImg1_384_EXMPLR, 
      OutputImg1_383_EXMPLR, OutputImg1_382_EXMPLR, OutputImg1_381_EXMPLR, 
      OutputImg1_380_EXMPLR, OutputImg1_379_EXMPLR, OutputImg1_378_EXMPLR, 
      OutputImg1_377_EXMPLR, OutputImg1_376_EXMPLR, OutputImg1_375_EXMPLR, 
      OutputImg1_374_EXMPLR, OutputImg1_373_EXMPLR, OutputImg1_372_EXMPLR, 
      OutputImg1_371_EXMPLR, OutputImg1_370_EXMPLR, OutputImg1_369_EXMPLR, 
      OutputImg1_368_EXMPLR, OutputImg1_367_EXMPLR, OutputImg1_366_EXMPLR, 
      OutputImg1_365_EXMPLR, OutputImg1_364_EXMPLR, OutputImg1_363_EXMPLR, 
      OutputImg1_362_EXMPLR, OutputImg1_361_EXMPLR, OutputImg1_360_EXMPLR, 
      OutputImg1_359_EXMPLR, OutputImg1_358_EXMPLR, OutputImg1_357_EXMPLR, 
      OutputImg1_356_EXMPLR, OutputImg1_355_EXMPLR, OutputImg1_354_EXMPLR, 
      OutputImg1_353_EXMPLR, OutputImg1_352_EXMPLR, OutputImg1_351_EXMPLR, 
      OutputImg1_350_EXMPLR, OutputImg1_349_EXMPLR, OutputImg1_348_EXMPLR, 
      OutputImg1_347_EXMPLR, OutputImg1_346_EXMPLR, OutputImg1_345_EXMPLR, 
      OutputImg1_344_EXMPLR, OutputImg1_343_EXMPLR, OutputImg1_342_EXMPLR, 
      OutputImg1_341_EXMPLR, OutputImg1_340_EXMPLR, OutputImg1_339_EXMPLR, 
      OutputImg1_338_EXMPLR, OutputImg1_337_EXMPLR, OutputImg1_336_EXMPLR, 
      OutputImg1_335_EXMPLR, OutputImg1_334_EXMPLR, OutputImg1_333_EXMPLR, 
      OutputImg1_332_EXMPLR, OutputImg1_331_EXMPLR, OutputImg1_330_EXMPLR, 
      OutputImg1_329_EXMPLR, OutputImg1_328_EXMPLR, OutputImg1_327_EXMPLR, 
      OutputImg1_326_EXMPLR, OutputImg1_325_EXMPLR, OutputImg1_324_EXMPLR, 
      OutputImg1_323_EXMPLR, OutputImg1_322_EXMPLR, OutputImg1_321_EXMPLR, 
      OutputImg1_320_EXMPLR, OutputImg1_319_EXMPLR, OutputImg1_318_EXMPLR, 
      OutputImg1_317_EXMPLR, OutputImg1_316_EXMPLR, OutputImg1_315_EXMPLR, 
      OutputImg1_314_EXMPLR, OutputImg1_313_EXMPLR, OutputImg1_312_EXMPLR, 
      OutputImg1_311_EXMPLR, OutputImg1_310_EXMPLR, OutputImg1_309_EXMPLR, 
      OutputImg1_308_EXMPLR, OutputImg1_307_EXMPLR, OutputImg1_306_EXMPLR, 
      OutputImg1_305_EXMPLR, OutputImg1_304_EXMPLR, OutputImg1_303_EXMPLR, 
      OutputImg1_302_EXMPLR, OutputImg1_301_EXMPLR, OutputImg1_300_EXMPLR, 
      OutputImg1_299_EXMPLR, OutputImg1_298_EXMPLR, OutputImg1_297_EXMPLR, 
      OutputImg1_296_EXMPLR, OutputImg1_295_EXMPLR, OutputImg1_294_EXMPLR, 
      OutputImg1_293_EXMPLR, OutputImg1_292_EXMPLR, OutputImg1_291_EXMPLR, 
      OutputImg1_290_EXMPLR, OutputImg1_289_EXMPLR, OutputImg1_288_EXMPLR, 
      OutputImg1_287_EXMPLR, OutputImg1_286_EXMPLR, OutputImg1_285_EXMPLR, 
      OutputImg1_284_EXMPLR, OutputImg1_283_EXMPLR, OutputImg1_282_EXMPLR, 
      OutputImg1_281_EXMPLR, OutputImg1_280_EXMPLR, OutputImg1_279_EXMPLR, 
      OutputImg1_278_EXMPLR, OutputImg1_277_EXMPLR, OutputImg1_276_EXMPLR, 
      OutputImg1_275_EXMPLR, OutputImg1_274_EXMPLR, OutputImg1_273_EXMPLR, 
      OutputImg1_272_EXMPLR, OutputImg1_271_EXMPLR, OutputImg1_270_EXMPLR, 
      OutputImg1_269_EXMPLR, OutputImg1_268_EXMPLR, OutputImg1_267_EXMPLR, 
      OutputImg1_266_EXMPLR, OutputImg1_265_EXMPLR, OutputImg1_264_EXMPLR, 
      OutputImg1_263_EXMPLR, OutputImg1_262_EXMPLR, OutputImg1_261_EXMPLR, 
      OutputImg1_260_EXMPLR, OutputImg1_259_EXMPLR, OutputImg1_258_EXMPLR, 
      OutputImg1_257_EXMPLR, OutputImg1_256_EXMPLR, OutputImg1_255_EXMPLR, 
      OutputImg1_254_EXMPLR, OutputImg1_253_EXMPLR, OutputImg1_252_EXMPLR, 
      OutputImg1_251_EXMPLR, OutputImg1_250_EXMPLR, OutputImg1_249_EXMPLR, 
      OutputImg1_248_EXMPLR, OutputImg1_247_EXMPLR, OutputImg1_246_EXMPLR, 
      OutputImg1_245_EXMPLR, OutputImg1_244_EXMPLR, OutputImg1_243_EXMPLR, 
      OutputImg1_242_EXMPLR, OutputImg1_241_EXMPLR, OutputImg1_240_EXMPLR, 
      OutputImg1_239_EXMPLR, OutputImg1_238_EXMPLR, OutputImg1_237_EXMPLR, 
      OutputImg1_236_EXMPLR, OutputImg1_235_EXMPLR, OutputImg1_234_EXMPLR, 
      OutputImg1_233_EXMPLR, OutputImg1_232_EXMPLR, OutputImg1_231_EXMPLR, 
      OutputImg1_230_EXMPLR, OutputImg1_229_EXMPLR, OutputImg1_228_EXMPLR, 
      OutputImg1_227_EXMPLR, OutputImg1_226_EXMPLR, OutputImg1_225_EXMPLR, 
      OutputImg1_224_EXMPLR, OutputImg1_223_EXMPLR, OutputImg1_222_EXMPLR, 
      OutputImg1_221_EXMPLR, OutputImg1_220_EXMPLR, OutputImg1_219_EXMPLR, 
      OutputImg1_218_EXMPLR, OutputImg1_217_EXMPLR, OutputImg1_216_EXMPLR, 
      OutputImg1_215_EXMPLR, OutputImg1_214_EXMPLR, OutputImg1_213_EXMPLR, 
      OutputImg1_212_EXMPLR, OutputImg1_211_EXMPLR, OutputImg1_210_EXMPLR, 
      OutputImg1_209_EXMPLR, OutputImg1_208_EXMPLR, OutputImg1_207_EXMPLR, 
      OutputImg1_206_EXMPLR, OutputImg1_205_EXMPLR, OutputImg1_204_EXMPLR, 
      OutputImg1_203_EXMPLR, OutputImg1_202_EXMPLR, OutputImg1_201_EXMPLR, 
      OutputImg1_200_EXMPLR, OutputImg1_199_EXMPLR, OutputImg1_198_EXMPLR, 
      OutputImg1_197_EXMPLR, OutputImg1_196_EXMPLR, OutputImg1_195_EXMPLR, 
      OutputImg1_194_EXMPLR, OutputImg1_193_EXMPLR, OutputImg1_192_EXMPLR, 
      OutputImg1_191_EXMPLR, OutputImg1_190_EXMPLR, OutputImg1_189_EXMPLR, 
      OutputImg1_188_EXMPLR, OutputImg1_187_EXMPLR, OutputImg1_186_EXMPLR, 
      OutputImg1_185_EXMPLR, OutputImg1_184_EXMPLR, OutputImg1_183_EXMPLR, 
      OutputImg1_182_EXMPLR, OutputImg1_181_EXMPLR, OutputImg1_180_EXMPLR, 
      OutputImg1_179_EXMPLR, OutputImg1_178_EXMPLR, OutputImg1_177_EXMPLR, 
      OutputImg1_176_EXMPLR, OutputImg1_175_EXMPLR, OutputImg1_174_EXMPLR, 
      OutputImg1_173_EXMPLR, OutputImg1_172_EXMPLR, OutputImg1_171_EXMPLR, 
      OutputImg1_170_EXMPLR, OutputImg1_169_EXMPLR, OutputImg1_168_EXMPLR, 
      OutputImg1_167_EXMPLR, OutputImg1_166_EXMPLR, OutputImg1_165_EXMPLR, 
      OutputImg1_164_EXMPLR, OutputImg1_163_EXMPLR, OutputImg1_162_EXMPLR, 
      OutputImg1_161_EXMPLR, OutputImg1_160_EXMPLR, OutputImg1_159_EXMPLR, 
      OutputImg1_158_EXMPLR, OutputImg1_157_EXMPLR, OutputImg1_156_EXMPLR, 
      OutputImg1_155_EXMPLR, OutputImg1_154_EXMPLR, OutputImg1_153_EXMPLR, 
      OutputImg1_152_EXMPLR, OutputImg1_151_EXMPLR, OutputImg1_150_EXMPLR, 
      OutputImg1_149_EXMPLR, OutputImg1_148_EXMPLR, OutputImg1_147_EXMPLR, 
      OutputImg1_146_EXMPLR, OutputImg1_145_EXMPLR, OutputImg1_144_EXMPLR, 
      OutputImg1_143_EXMPLR, OutputImg1_142_EXMPLR, OutputImg1_141_EXMPLR, 
      OutputImg1_140_EXMPLR, OutputImg1_139_EXMPLR, OutputImg1_138_EXMPLR, 
      OutputImg1_137_EXMPLR, OutputImg1_136_EXMPLR, OutputImg1_135_EXMPLR, 
      OutputImg1_134_EXMPLR, OutputImg1_133_EXMPLR, OutputImg1_132_EXMPLR, 
      OutputImg1_131_EXMPLR, OutputImg1_130_EXMPLR, OutputImg1_129_EXMPLR, 
      OutputImg1_128_EXMPLR, OutputImg1_127_EXMPLR, OutputImg1_126_EXMPLR, 
      OutputImg1_125_EXMPLR, OutputImg1_124_EXMPLR, OutputImg1_123_EXMPLR, 
      OutputImg1_122_EXMPLR, OutputImg1_121_EXMPLR, OutputImg1_120_EXMPLR, 
      OutputImg1_119_EXMPLR, OutputImg1_118_EXMPLR, OutputImg1_117_EXMPLR, 
      OutputImg1_116_EXMPLR, OutputImg1_115_EXMPLR, OutputImg1_114_EXMPLR, 
      OutputImg1_113_EXMPLR, OutputImg1_112_EXMPLR, OutputImg1_111_EXMPLR, 
      OutputImg1_110_EXMPLR, OutputImg1_109_EXMPLR, OutputImg1_108_EXMPLR, 
      OutputImg1_107_EXMPLR, OutputImg1_106_EXMPLR, OutputImg1_105_EXMPLR, 
      OutputImg1_104_EXMPLR, OutputImg1_103_EXMPLR, OutputImg1_102_EXMPLR, 
      OutputImg1_101_EXMPLR, OutputImg1_100_EXMPLR, OutputImg1_99_EXMPLR, 
      OutputImg1_98_EXMPLR, OutputImg1_97_EXMPLR, OutputImg1_96_EXMPLR, 
      OutputImg1_95_EXMPLR, OutputImg1_94_EXMPLR, OutputImg1_93_EXMPLR, 
      OutputImg1_92_EXMPLR, OutputImg1_91_EXMPLR, OutputImg1_90_EXMPLR, 
      OutputImg1_89_EXMPLR, OutputImg1_88_EXMPLR, OutputImg1_87_EXMPLR, 
      OutputImg1_86_EXMPLR, OutputImg1_85_EXMPLR, OutputImg1_84_EXMPLR, 
      OutputImg1_83_EXMPLR, OutputImg1_82_EXMPLR, OutputImg1_81_EXMPLR, 
      OutputImg1_80_EXMPLR, OutputImg1_79_EXMPLR, OutputImg1_78_EXMPLR, 
      OutputImg1_77_EXMPLR, OutputImg1_76_EXMPLR, OutputImg1_75_EXMPLR, 
      OutputImg1_74_EXMPLR, OutputImg1_73_EXMPLR, OutputImg1_72_EXMPLR, 
      OutputImg1_71_EXMPLR, OutputImg1_70_EXMPLR, OutputImg1_69_EXMPLR, 
      OutputImg1_68_EXMPLR, OutputImg1_67_EXMPLR, OutputImg1_66_EXMPLR, 
      OutputImg1_65_EXMPLR, OutputImg1_64_EXMPLR, OutputImg1_63_EXMPLR, 
      OutputImg1_62_EXMPLR, OutputImg1_61_EXMPLR, OutputImg1_60_EXMPLR, 
      OutputImg1_59_EXMPLR, OutputImg1_58_EXMPLR, OutputImg1_57_EXMPLR, 
      OutputImg1_56_EXMPLR, OutputImg1_55_EXMPLR, OutputImg1_54_EXMPLR, 
      OutputImg1_53_EXMPLR, OutputImg1_52_EXMPLR, OutputImg1_51_EXMPLR, 
      OutputImg1_50_EXMPLR, OutputImg1_49_EXMPLR, OutputImg1_48_EXMPLR, 
      OutputImg1_47_EXMPLR, OutputImg1_46_EXMPLR, OutputImg1_45_EXMPLR, 
      OutputImg1_44_EXMPLR, OutputImg1_43_EXMPLR, OutputImg1_42_EXMPLR, 
      OutputImg1_41_EXMPLR, OutputImg1_40_EXMPLR, OutputImg1_39_EXMPLR, 
      OutputImg1_38_EXMPLR, OutputImg1_37_EXMPLR, OutputImg1_36_EXMPLR, 
      OutputImg1_35_EXMPLR, OutputImg1_34_EXMPLR, OutputImg1_33_EXMPLR, 
      OutputImg1_32_EXMPLR, OutputImg1_31_EXMPLR, OutputImg1_30_EXMPLR, 
      OutputImg1_29_EXMPLR, OutputImg1_28_EXMPLR, OutputImg1_27_EXMPLR, 
      OutputImg1_26_EXMPLR, OutputImg1_25_EXMPLR, OutputImg1_24_EXMPLR, 
      OutputImg1_23_EXMPLR, OutputImg1_22_EXMPLR, OutputImg1_21_EXMPLR, 
      OutputImg1_20_EXMPLR, OutputImg1_19_EXMPLR, OutputImg1_18_EXMPLR, 
      OutputImg1_17_EXMPLR, OutputImg1_16_EXMPLR, OutputImg1_15_EXMPLR, 
      OutputImg1_14_EXMPLR, OutputImg1_13_EXMPLR, OutputImg1_12_EXMPLR, 
      OutputImg1_11_EXMPLR, OutputImg1_10_EXMPLR, OutputImg1_9_EXMPLR, 
      OutputImg1_8_EXMPLR, OutputImg1_7_EXMPLR, OutputImg1_6_EXMPLR, 
      OutputImg1_5_EXMPLR, OutputImg1_4_EXMPLR, OutputImg1_3_EXMPLR, 
      OutputImg1_2_EXMPLR, OutputImg1_1_EXMPLR, OutputImg1_0_EXMPLR, 
      OutputImg2_447_EXMPLR, OutputImg2_446_EXMPLR, OutputImg2_445_EXMPLR, 
      OutputImg2_444_EXMPLR, OutputImg2_443_EXMPLR, OutputImg2_442_EXMPLR, 
      OutputImg2_441_EXMPLR, OutputImg2_440_EXMPLR, OutputImg2_439_EXMPLR, 
      OutputImg2_438_EXMPLR, OutputImg2_437_EXMPLR, OutputImg2_436_EXMPLR, 
      OutputImg2_435_EXMPLR, OutputImg2_434_EXMPLR, OutputImg2_433_EXMPLR, 
      OutputImg2_432_EXMPLR, OutputImg2_431_EXMPLR, OutputImg2_430_EXMPLR, 
      OutputImg2_429_EXMPLR, OutputImg2_428_EXMPLR, OutputImg2_427_EXMPLR, 
      OutputImg2_426_EXMPLR, OutputImg2_425_EXMPLR, OutputImg2_424_EXMPLR, 
      OutputImg2_423_EXMPLR, OutputImg2_422_EXMPLR, OutputImg2_421_EXMPLR, 
      OutputImg2_420_EXMPLR, OutputImg2_419_EXMPLR, OutputImg2_418_EXMPLR, 
      OutputImg2_417_EXMPLR, OutputImg2_416_EXMPLR, OutputImg2_415_EXMPLR, 
      OutputImg2_414_EXMPLR, OutputImg2_413_EXMPLR, OutputImg2_412_EXMPLR, 
      OutputImg2_411_EXMPLR, OutputImg2_410_EXMPLR, OutputImg2_409_EXMPLR, 
      OutputImg2_408_EXMPLR, OutputImg2_407_EXMPLR, OutputImg2_406_EXMPLR, 
      OutputImg2_405_EXMPLR, OutputImg2_404_EXMPLR, OutputImg2_403_EXMPLR, 
      OutputImg2_402_EXMPLR, OutputImg2_401_EXMPLR, OutputImg2_400_EXMPLR, 
      OutputImg2_399_EXMPLR, OutputImg2_398_EXMPLR, OutputImg2_397_EXMPLR, 
      OutputImg2_396_EXMPLR, OutputImg2_395_EXMPLR, OutputImg2_394_EXMPLR, 
      OutputImg2_393_EXMPLR, OutputImg2_392_EXMPLR, OutputImg2_391_EXMPLR, 
      OutputImg2_390_EXMPLR, OutputImg2_389_EXMPLR, OutputImg2_388_EXMPLR, 
      OutputImg2_387_EXMPLR, OutputImg2_386_EXMPLR, OutputImg2_385_EXMPLR, 
      OutputImg2_384_EXMPLR, OutputImg2_383_EXMPLR, OutputImg2_382_EXMPLR, 
      OutputImg2_381_EXMPLR, OutputImg2_380_EXMPLR, OutputImg2_379_EXMPLR, 
      OutputImg2_378_EXMPLR, OutputImg2_377_EXMPLR, OutputImg2_376_EXMPLR, 
      OutputImg2_375_EXMPLR, OutputImg2_374_EXMPLR, OutputImg2_373_EXMPLR, 
      OutputImg2_372_EXMPLR, OutputImg2_371_EXMPLR, OutputImg2_370_EXMPLR, 
      OutputImg2_369_EXMPLR, OutputImg2_368_EXMPLR, OutputImg2_367_EXMPLR, 
      OutputImg2_366_EXMPLR, OutputImg2_365_EXMPLR, OutputImg2_364_EXMPLR, 
      OutputImg2_363_EXMPLR, OutputImg2_362_EXMPLR, OutputImg2_361_EXMPLR, 
      OutputImg2_360_EXMPLR, OutputImg2_359_EXMPLR, OutputImg2_358_EXMPLR, 
      OutputImg2_357_EXMPLR, OutputImg2_356_EXMPLR, OutputImg2_355_EXMPLR, 
      OutputImg2_354_EXMPLR, OutputImg2_353_EXMPLR, OutputImg2_352_EXMPLR, 
      OutputImg2_351_EXMPLR, OutputImg2_350_EXMPLR, OutputImg2_349_EXMPLR, 
      OutputImg2_348_EXMPLR, OutputImg2_347_EXMPLR, OutputImg2_346_EXMPLR, 
      OutputImg2_345_EXMPLR, OutputImg2_344_EXMPLR, OutputImg2_343_EXMPLR, 
      OutputImg2_342_EXMPLR, OutputImg2_341_EXMPLR, OutputImg2_340_EXMPLR, 
      OutputImg2_339_EXMPLR, OutputImg2_338_EXMPLR, OutputImg2_337_EXMPLR, 
      OutputImg2_336_EXMPLR, OutputImg2_335_EXMPLR, OutputImg2_334_EXMPLR, 
      OutputImg2_333_EXMPLR, OutputImg2_332_EXMPLR, OutputImg2_331_EXMPLR, 
      OutputImg2_330_EXMPLR, OutputImg2_329_EXMPLR, OutputImg2_328_EXMPLR, 
      OutputImg2_327_EXMPLR, OutputImg2_326_EXMPLR, OutputImg2_325_EXMPLR, 
      OutputImg2_324_EXMPLR, OutputImg2_323_EXMPLR, OutputImg2_322_EXMPLR, 
      OutputImg2_321_EXMPLR, OutputImg2_320_EXMPLR, OutputImg2_319_EXMPLR, 
      OutputImg2_318_EXMPLR, OutputImg2_317_EXMPLR, OutputImg2_316_EXMPLR, 
      OutputImg2_315_EXMPLR, OutputImg2_314_EXMPLR, OutputImg2_313_EXMPLR, 
      OutputImg2_312_EXMPLR, OutputImg2_311_EXMPLR, OutputImg2_310_EXMPLR, 
      OutputImg2_309_EXMPLR, OutputImg2_308_EXMPLR, OutputImg2_307_EXMPLR, 
      OutputImg2_306_EXMPLR, OutputImg2_305_EXMPLR, OutputImg2_304_EXMPLR, 
      OutputImg2_303_EXMPLR, OutputImg2_302_EXMPLR, OutputImg2_301_EXMPLR, 
      OutputImg2_300_EXMPLR, OutputImg2_299_EXMPLR, OutputImg2_298_EXMPLR, 
      OutputImg2_297_EXMPLR, OutputImg2_296_EXMPLR, OutputImg2_295_EXMPLR, 
      OutputImg2_294_EXMPLR, OutputImg2_293_EXMPLR, OutputImg2_292_EXMPLR, 
      OutputImg2_291_EXMPLR, OutputImg2_290_EXMPLR, OutputImg2_289_EXMPLR, 
      OutputImg2_288_EXMPLR, OutputImg2_287_EXMPLR, OutputImg2_286_EXMPLR, 
      OutputImg2_285_EXMPLR, OutputImg2_284_EXMPLR, OutputImg2_283_EXMPLR, 
      OutputImg2_282_EXMPLR, OutputImg2_281_EXMPLR, OutputImg2_280_EXMPLR, 
      OutputImg2_279_EXMPLR, OutputImg2_278_EXMPLR, OutputImg2_277_EXMPLR, 
      OutputImg2_276_EXMPLR, OutputImg2_275_EXMPLR, OutputImg2_274_EXMPLR, 
      OutputImg2_273_EXMPLR, OutputImg2_272_EXMPLR, OutputImg2_271_EXMPLR, 
      OutputImg2_270_EXMPLR, OutputImg2_269_EXMPLR, OutputImg2_268_EXMPLR, 
      OutputImg2_267_EXMPLR, OutputImg2_266_EXMPLR, OutputImg2_265_EXMPLR, 
      OutputImg2_264_EXMPLR, OutputImg2_263_EXMPLR, OutputImg2_262_EXMPLR, 
      OutputImg2_261_EXMPLR, OutputImg2_260_EXMPLR, OutputImg2_259_EXMPLR, 
      OutputImg2_258_EXMPLR, OutputImg2_257_EXMPLR, OutputImg2_256_EXMPLR, 
      OutputImg2_255_EXMPLR, OutputImg2_254_EXMPLR, OutputImg2_253_EXMPLR, 
      OutputImg2_252_EXMPLR, OutputImg2_251_EXMPLR, OutputImg2_250_EXMPLR, 
      OutputImg2_249_EXMPLR, OutputImg2_248_EXMPLR, OutputImg2_247_EXMPLR, 
      OutputImg2_246_EXMPLR, OutputImg2_245_EXMPLR, OutputImg2_244_EXMPLR, 
      OutputImg2_243_EXMPLR, OutputImg2_242_EXMPLR, OutputImg2_241_EXMPLR, 
      OutputImg2_240_EXMPLR, OutputImg2_239_EXMPLR, OutputImg2_238_EXMPLR, 
      OutputImg2_237_EXMPLR, OutputImg2_236_EXMPLR, OutputImg2_235_EXMPLR, 
      OutputImg2_234_EXMPLR, OutputImg2_233_EXMPLR, OutputImg2_232_EXMPLR, 
      OutputImg2_231_EXMPLR, OutputImg2_230_EXMPLR, OutputImg2_229_EXMPLR, 
      OutputImg2_228_EXMPLR, OutputImg2_227_EXMPLR, OutputImg2_226_EXMPLR, 
      OutputImg2_225_EXMPLR, OutputImg2_224_EXMPLR, OutputImg2_223_EXMPLR, 
      OutputImg2_222_EXMPLR, OutputImg2_221_EXMPLR, OutputImg2_220_EXMPLR, 
      OutputImg2_219_EXMPLR, OutputImg2_218_EXMPLR, OutputImg2_217_EXMPLR, 
      OutputImg2_216_EXMPLR, OutputImg2_215_EXMPLR, OutputImg2_214_EXMPLR, 
      OutputImg2_213_EXMPLR, OutputImg2_212_EXMPLR, OutputImg2_211_EXMPLR, 
      OutputImg2_210_EXMPLR, OutputImg2_209_EXMPLR, OutputImg2_208_EXMPLR, 
      OutputImg2_207_EXMPLR, OutputImg2_206_EXMPLR, OutputImg2_205_EXMPLR, 
      OutputImg2_204_EXMPLR, OutputImg2_203_EXMPLR, OutputImg2_202_EXMPLR, 
      OutputImg2_201_EXMPLR, OutputImg2_200_EXMPLR, OutputImg2_199_EXMPLR, 
      OutputImg2_198_EXMPLR, OutputImg2_197_EXMPLR, OutputImg2_196_EXMPLR, 
      OutputImg2_195_EXMPLR, OutputImg2_194_EXMPLR, OutputImg2_193_EXMPLR, 
      OutputImg2_192_EXMPLR, OutputImg2_191_EXMPLR, OutputImg2_190_EXMPLR, 
      OutputImg2_189_EXMPLR, OutputImg2_188_EXMPLR, OutputImg2_187_EXMPLR, 
      OutputImg2_186_EXMPLR, OutputImg2_185_EXMPLR, OutputImg2_184_EXMPLR, 
      OutputImg2_183_EXMPLR, OutputImg2_182_EXMPLR, OutputImg2_181_EXMPLR, 
      OutputImg2_180_EXMPLR, OutputImg2_179_EXMPLR, OutputImg2_178_EXMPLR, 
      OutputImg2_177_EXMPLR, OutputImg2_176_EXMPLR, OutputImg2_175_EXMPLR, 
      OutputImg2_174_EXMPLR, OutputImg2_173_EXMPLR, OutputImg2_172_EXMPLR, 
      OutputImg2_171_EXMPLR, OutputImg2_170_EXMPLR, OutputImg2_169_EXMPLR, 
      OutputImg2_168_EXMPLR, OutputImg2_167_EXMPLR, OutputImg2_166_EXMPLR, 
      OutputImg2_165_EXMPLR, OutputImg2_164_EXMPLR, OutputImg2_163_EXMPLR, 
      OutputImg2_162_EXMPLR, OutputImg2_161_EXMPLR, OutputImg2_160_EXMPLR, 
      OutputImg2_159_EXMPLR, OutputImg2_158_EXMPLR, OutputImg2_157_EXMPLR, 
      OutputImg2_156_EXMPLR, OutputImg2_155_EXMPLR, OutputImg2_154_EXMPLR, 
      OutputImg2_153_EXMPLR, OutputImg2_152_EXMPLR, OutputImg2_151_EXMPLR, 
      OutputImg2_150_EXMPLR, OutputImg2_149_EXMPLR, OutputImg2_148_EXMPLR, 
      OutputImg2_147_EXMPLR, OutputImg2_146_EXMPLR, OutputImg2_145_EXMPLR, 
      OutputImg2_144_EXMPLR, OutputImg2_143_EXMPLR, OutputImg2_142_EXMPLR, 
      OutputImg2_141_EXMPLR, OutputImg2_140_EXMPLR, OutputImg2_139_EXMPLR, 
      OutputImg2_138_EXMPLR, OutputImg2_137_EXMPLR, OutputImg2_136_EXMPLR, 
      OutputImg2_135_EXMPLR, OutputImg2_134_EXMPLR, OutputImg2_133_EXMPLR, 
      OutputImg2_132_EXMPLR, OutputImg2_131_EXMPLR, OutputImg2_130_EXMPLR, 
      OutputImg2_129_EXMPLR, OutputImg2_128_EXMPLR, OutputImg2_127_EXMPLR, 
      OutputImg2_126_EXMPLR, OutputImg2_125_EXMPLR, OutputImg2_124_EXMPLR, 
      OutputImg2_123_EXMPLR, OutputImg2_122_EXMPLR, OutputImg2_121_EXMPLR, 
      OutputImg2_120_EXMPLR, OutputImg2_119_EXMPLR, OutputImg2_118_EXMPLR, 
      OutputImg2_117_EXMPLR, OutputImg2_116_EXMPLR, OutputImg2_115_EXMPLR, 
      OutputImg2_114_EXMPLR, OutputImg2_113_EXMPLR, OutputImg2_112_EXMPLR, 
      OutputImg2_111_EXMPLR, OutputImg2_110_EXMPLR, OutputImg2_109_EXMPLR, 
      OutputImg2_108_EXMPLR, OutputImg2_107_EXMPLR, OutputImg2_106_EXMPLR, 
      OutputImg2_105_EXMPLR, OutputImg2_104_EXMPLR, OutputImg2_103_EXMPLR, 
      OutputImg2_102_EXMPLR, OutputImg2_101_EXMPLR, OutputImg2_100_EXMPLR, 
      OutputImg2_99_EXMPLR, OutputImg2_98_EXMPLR, OutputImg2_97_EXMPLR, 
      OutputImg2_96_EXMPLR, OutputImg2_95_EXMPLR, OutputImg2_94_EXMPLR, 
      OutputImg2_93_EXMPLR, OutputImg2_92_EXMPLR, OutputImg2_91_EXMPLR, 
      OutputImg2_90_EXMPLR, OutputImg2_89_EXMPLR, OutputImg2_88_EXMPLR, 
      OutputImg2_87_EXMPLR, OutputImg2_86_EXMPLR, OutputImg2_85_EXMPLR, 
      OutputImg2_84_EXMPLR, OutputImg2_83_EXMPLR, OutputImg2_82_EXMPLR, 
      OutputImg2_81_EXMPLR, OutputImg2_80_EXMPLR, OutputImg2_79_EXMPLR, 
      OutputImg2_78_EXMPLR, OutputImg2_77_EXMPLR, OutputImg2_76_EXMPLR, 
      OutputImg2_75_EXMPLR, OutputImg2_74_EXMPLR, OutputImg2_73_EXMPLR, 
      OutputImg2_72_EXMPLR, OutputImg2_71_EXMPLR, OutputImg2_70_EXMPLR, 
      OutputImg2_69_EXMPLR, OutputImg2_68_EXMPLR, OutputImg2_67_EXMPLR, 
      OutputImg2_66_EXMPLR, OutputImg2_65_EXMPLR, OutputImg2_64_EXMPLR, 
      OutputImg2_63_EXMPLR, OutputImg2_62_EXMPLR, OutputImg2_61_EXMPLR, 
      OutputImg2_60_EXMPLR, OutputImg2_59_EXMPLR, OutputImg2_58_EXMPLR, 
      OutputImg2_57_EXMPLR, OutputImg2_56_EXMPLR, OutputImg2_55_EXMPLR, 
      OutputImg2_54_EXMPLR, OutputImg2_53_EXMPLR, OutputImg2_52_EXMPLR, 
      OutputImg2_51_EXMPLR, OutputImg2_50_EXMPLR, OutputImg2_49_EXMPLR, 
      OutputImg2_48_EXMPLR, OutputImg2_47_EXMPLR, OutputImg2_46_EXMPLR, 
      OutputImg2_45_EXMPLR, OutputImg2_44_EXMPLR, OutputImg2_43_EXMPLR, 
      OutputImg2_42_EXMPLR, OutputImg2_41_EXMPLR, OutputImg2_40_EXMPLR, 
      OutputImg2_39_EXMPLR, OutputImg2_38_EXMPLR, OutputImg2_37_EXMPLR, 
      OutputImg2_36_EXMPLR, OutputImg2_35_EXMPLR, OutputImg2_34_EXMPLR, 
      OutputImg2_33_EXMPLR, OutputImg2_32_EXMPLR, OutputImg2_31_EXMPLR, 
      OutputImg2_30_EXMPLR, OutputImg2_29_EXMPLR, OutputImg2_28_EXMPLR, 
      OutputImg2_27_EXMPLR, OutputImg2_26_EXMPLR, OutputImg2_25_EXMPLR, 
      OutputImg2_24_EXMPLR, OutputImg2_23_EXMPLR, OutputImg2_22_EXMPLR, 
      OutputImg2_21_EXMPLR, OutputImg2_20_EXMPLR, OutputImg2_19_EXMPLR, 
      OutputImg2_18_EXMPLR, OutputImg2_17_EXMPLR, OutputImg2_16_EXMPLR, 
      OutputImg2_15_EXMPLR, OutputImg2_14_EXMPLR, OutputImg2_13_EXMPLR, 
      OutputImg2_12_EXMPLR, OutputImg2_11_EXMPLR, OutputImg2_10_EXMPLR, 
      OutputImg2_9_EXMPLR, OutputImg2_8_EXMPLR, OutputImg2_7_EXMPLR, 
      OutputImg2_6_EXMPLR, OutputImg2_5_EXMPLR, OutputImg2_4_EXMPLR, 
      OutputImg2_3_EXMPLR, OutputImg2_2_EXMPLR, OutputImg2_1_EXMPLR, 
      OutputImg2_0_EXMPLR, OutputImg3_447_EXMPLR, OutputImg3_446_EXMPLR, 
      OutputImg3_445_EXMPLR, OutputImg3_444_EXMPLR, OutputImg3_443_EXMPLR, 
      OutputImg3_442_EXMPLR, OutputImg3_441_EXMPLR, OutputImg3_440_EXMPLR, 
      OutputImg3_439_EXMPLR, OutputImg3_438_EXMPLR, OutputImg3_437_EXMPLR, 
      OutputImg3_436_EXMPLR, OutputImg3_435_EXMPLR, OutputImg3_434_EXMPLR, 
      OutputImg3_433_EXMPLR, OutputImg3_432_EXMPLR, OutputImg3_431_EXMPLR, 
      OutputImg3_430_EXMPLR, OutputImg3_429_EXMPLR, OutputImg3_428_EXMPLR, 
      OutputImg3_427_EXMPLR, OutputImg3_426_EXMPLR, OutputImg3_425_EXMPLR, 
      OutputImg3_424_EXMPLR, OutputImg3_423_EXMPLR, OutputImg3_422_EXMPLR, 
      OutputImg3_421_EXMPLR, OutputImg3_420_EXMPLR, OutputImg3_419_EXMPLR, 
      OutputImg3_418_EXMPLR, OutputImg3_417_EXMPLR, OutputImg3_416_EXMPLR, 
      OutputImg3_415_EXMPLR, OutputImg3_414_EXMPLR, OutputImg3_413_EXMPLR, 
      OutputImg3_412_EXMPLR, OutputImg3_411_EXMPLR, OutputImg3_410_EXMPLR, 
      OutputImg3_409_EXMPLR, OutputImg3_408_EXMPLR, OutputImg3_407_EXMPLR, 
      OutputImg3_406_EXMPLR, OutputImg3_405_EXMPLR, OutputImg3_404_EXMPLR, 
      OutputImg3_403_EXMPLR, OutputImg3_402_EXMPLR, OutputImg3_401_EXMPLR, 
      OutputImg3_400_EXMPLR, OutputImg3_399_EXMPLR, OutputImg3_398_EXMPLR, 
      OutputImg3_397_EXMPLR, OutputImg3_396_EXMPLR, OutputImg3_395_EXMPLR, 
      OutputImg3_394_EXMPLR, OutputImg3_393_EXMPLR, OutputImg3_392_EXMPLR, 
      OutputImg3_391_EXMPLR, OutputImg3_390_EXMPLR, OutputImg3_389_EXMPLR, 
      OutputImg3_388_EXMPLR, OutputImg3_387_EXMPLR, OutputImg3_386_EXMPLR, 
      OutputImg3_385_EXMPLR, OutputImg3_384_EXMPLR, OutputImg3_383_EXMPLR, 
      OutputImg3_382_EXMPLR, OutputImg3_381_EXMPLR, OutputImg3_380_EXMPLR, 
      OutputImg3_379_EXMPLR, OutputImg3_378_EXMPLR, OutputImg3_377_EXMPLR, 
      OutputImg3_376_EXMPLR, OutputImg3_375_EXMPLR, OutputImg3_374_EXMPLR, 
      OutputImg3_373_EXMPLR, OutputImg3_372_EXMPLR, OutputImg3_371_EXMPLR, 
      OutputImg3_370_EXMPLR, OutputImg3_369_EXMPLR, OutputImg3_368_EXMPLR, 
      OutputImg3_367_EXMPLR, OutputImg3_366_EXMPLR, OutputImg3_365_EXMPLR, 
      OutputImg3_364_EXMPLR, OutputImg3_363_EXMPLR, OutputImg3_362_EXMPLR, 
      OutputImg3_361_EXMPLR, OutputImg3_360_EXMPLR, OutputImg3_359_EXMPLR, 
      OutputImg3_358_EXMPLR, OutputImg3_357_EXMPLR, OutputImg3_356_EXMPLR, 
      OutputImg3_355_EXMPLR, OutputImg3_354_EXMPLR, OutputImg3_353_EXMPLR, 
      OutputImg3_352_EXMPLR, OutputImg3_351_EXMPLR, OutputImg3_350_EXMPLR, 
      OutputImg3_349_EXMPLR, OutputImg3_348_EXMPLR, OutputImg3_347_EXMPLR, 
      OutputImg3_346_EXMPLR, OutputImg3_345_EXMPLR, OutputImg3_344_EXMPLR, 
      OutputImg3_343_EXMPLR, OutputImg3_342_EXMPLR, OutputImg3_341_EXMPLR, 
      OutputImg3_340_EXMPLR, OutputImg3_339_EXMPLR, OutputImg3_338_EXMPLR, 
      OutputImg3_337_EXMPLR, OutputImg3_336_EXMPLR, OutputImg3_335_EXMPLR, 
      OutputImg3_334_EXMPLR, OutputImg3_333_EXMPLR, OutputImg3_332_EXMPLR, 
      OutputImg3_331_EXMPLR, OutputImg3_330_EXMPLR, OutputImg3_329_EXMPLR, 
      OutputImg3_328_EXMPLR, OutputImg3_327_EXMPLR, OutputImg3_326_EXMPLR, 
      OutputImg3_325_EXMPLR, OutputImg3_324_EXMPLR, OutputImg3_323_EXMPLR, 
      OutputImg3_322_EXMPLR, OutputImg3_321_EXMPLR, OutputImg3_320_EXMPLR, 
      OutputImg3_319_EXMPLR, OutputImg3_318_EXMPLR, OutputImg3_317_EXMPLR, 
      OutputImg3_316_EXMPLR, OutputImg3_315_EXMPLR, OutputImg3_314_EXMPLR, 
      OutputImg3_313_EXMPLR, OutputImg3_312_EXMPLR, OutputImg3_311_EXMPLR, 
      OutputImg3_310_EXMPLR, OutputImg3_309_EXMPLR, OutputImg3_308_EXMPLR, 
      OutputImg3_307_EXMPLR, OutputImg3_306_EXMPLR, OutputImg3_305_EXMPLR, 
      OutputImg3_304_EXMPLR, OutputImg3_303_EXMPLR, OutputImg3_302_EXMPLR, 
      OutputImg3_301_EXMPLR, OutputImg3_300_EXMPLR, OutputImg3_299_EXMPLR, 
      OutputImg3_298_EXMPLR, OutputImg3_297_EXMPLR, OutputImg3_296_EXMPLR, 
      OutputImg3_295_EXMPLR, OutputImg3_294_EXMPLR, OutputImg3_293_EXMPLR, 
      OutputImg3_292_EXMPLR, OutputImg3_291_EXMPLR, OutputImg3_290_EXMPLR, 
      OutputImg3_289_EXMPLR, OutputImg3_288_EXMPLR, OutputImg3_287_EXMPLR, 
      OutputImg3_286_EXMPLR, OutputImg3_285_EXMPLR, OutputImg3_284_EXMPLR, 
      OutputImg3_283_EXMPLR, OutputImg3_282_EXMPLR, OutputImg3_281_EXMPLR, 
      OutputImg3_280_EXMPLR, OutputImg3_279_EXMPLR, OutputImg3_278_EXMPLR, 
      OutputImg3_277_EXMPLR, OutputImg3_276_EXMPLR, OutputImg3_275_EXMPLR, 
      OutputImg3_274_EXMPLR, OutputImg3_273_EXMPLR, OutputImg3_272_EXMPLR, 
      OutputImg3_271_EXMPLR, OutputImg3_270_EXMPLR, OutputImg3_269_EXMPLR, 
      OutputImg3_268_EXMPLR, OutputImg3_267_EXMPLR, OutputImg3_266_EXMPLR, 
      OutputImg3_265_EXMPLR, OutputImg3_264_EXMPLR, OutputImg3_263_EXMPLR, 
      OutputImg3_262_EXMPLR, OutputImg3_261_EXMPLR, OutputImg3_260_EXMPLR, 
      OutputImg3_259_EXMPLR, OutputImg3_258_EXMPLR, OutputImg3_257_EXMPLR, 
      OutputImg3_256_EXMPLR, OutputImg3_255_EXMPLR, OutputImg3_254_EXMPLR, 
      OutputImg3_253_EXMPLR, OutputImg3_252_EXMPLR, OutputImg3_251_EXMPLR, 
      OutputImg3_250_EXMPLR, OutputImg3_249_EXMPLR, OutputImg3_248_EXMPLR, 
      OutputImg3_247_EXMPLR, OutputImg3_246_EXMPLR, OutputImg3_245_EXMPLR, 
      OutputImg3_244_EXMPLR, OutputImg3_243_EXMPLR, OutputImg3_242_EXMPLR, 
      OutputImg3_241_EXMPLR, OutputImg3_240_EXMPLR, OutputImg3_239_EXMPLR, 
      OutputImg3_238_EXMPLR, OutputImg3_237_EXMPLR, OutputImg3_236_EXMPLR, 
      OutputImg3_235_EXMPLR, OutputImg3_234_EXMPLR, OutputImg3_233_EXMPLR, 
      OutputImg3_232_EXMPLR, OutputImg3_231_EXMPLR, OutputImg3_230_EXMPLR, 
      OutputImg3_229_EXMPLR, OutputImg3_228_EXMPLR, OutputImg3_227_EXMPLR, 
      OutputImg3_226_EXMPLR, OutputImg3_225_EXMPLR, OutputImg3_224_EXMPLR, 
      OutputImg3_223_EXMPLR, OutputImg3_222_EXMPLR, OutputImg3_221_EXMPLR, 
      OutputImg3_220_EXMPLR, OutputImg3_219_EXMPLR, OutputImg3_218_EXMPLR, 
      OutputImg3_217_EXMPLR, OutputImg3_216_EXMPLR, OutputImg3_215_EXMPLR, 
      OutputImg3_214_EXMPLR, OutputImg3_213_EXMPLR, OutputImg3_212_EXMPLR, 
      OutputImg3_211_EXMPLR, OutputImg3_210_EXMPLR, OutputImg3_209_EXMPLR, 
      OutputImg3_208_EXMPLR, OutputImg3_207_EXMPLR, OutputImg3_206_EXMPLR, 
      OutputImg3_205_EXMPLR, OutputImg3_204_EXMPLR, OutputImg3_203_EXMPLR, 
      OutputImg3_202_EXMPLR, OutputImg3_201_EXMPLR, OutputImg3_200_EXMPLR, 
      OutputImg3_199_EXMPLR, OutputImg3_198_EXMPLR, OutputImg3_197_EXMPLR, 
      OutputImg3_196_EXMPLR, OutputImg3_195_EXMPLR, OutputImg3_194_EXMPLR, 
      OutputImg3_193_EXMPLR, OutputImg3_192_EXMPLR, OutputImg3_191_EXMPLR, 
      OutputImg3_190_EXMPLR, OutputImg3_189_EXMPLR, OutputImg3_188_EXMPLR, 
      OutputImg3_187_EXMPLR, OutputImg3_186_EXMPLR, OutputImg3_185_EXMPLR, 
      OutputImg3_184_EXMPLR, OutputImg3_183_EXMPLR, OutputImg3_182_EXMPLR, 
      OutputImg3_181_EXMPLR, OutputImg3_180_EXMPLR, OutputImg3_179_EXMPLR, 
      OutputImg3_178_EXMPLR, OutputImg3_177_EXMPLR, OutputImg3_176_EXMPLR, 
      OutputImg3_175_EXMPLR, OutputImg3_174_EXMPLR, OutputImg3_173_EXMPLR, 
      OutputImg3_172_EXMPLR, OutputImg3_171_EXMPLR, OutputImg3_170_EXMPLR, 
      OutputImg3_169_EXMPLR, OutputImg3_168_EXMPLR, OutputImg3_167_EXMPLR, 
      OutputImg3_166_EXMPLR, OutputImg3_165_EXMPLR, OutputImg3_164_EXMPLR, 
      OutputImg3_163_EXMPLR, OutputImg3_162_EXMPLR, OutputImg3_161_EXMPLR, 
      OutputImg3_160_EXMPLR, OutputImg3_159_EXMPLR, OutputImg3_158_EXMPLR, 
      OutputImg3_157_EXMPLR, OutputImg3_156_EXMPLR, OutputImg3_155_EXMPLR, 
      OutputImg3_154_EXMPLR, OutputImg3_153_EXMPLR, OutputImg3_152_EXMPLR, 
      OutputImg3_151_EXMPLR, OutputImg3_150_EXMPLR, OutputImg3_149_EXMPLR, 
      OutputImg3_148_EXMPLR, OutputImg3_147_EXMPLR, OutputImg3_146_EXMPLR, 
      OutputImg3_145_EXMPLR, OutputImg3_144_EXMPLR, OutputImg3_143_EXMPLR, 
      OutputImg3_142_EXMPLR, OutputImg3_141_EXMPLR, OutputImg3_140_EXMPLR, 
      OutputImg3_139_EXMPLR, OutputImg3_138_EXMPLR, OutputImg3_137_EXMPLR, 
      OutputImg3_136_EXMPLR, OutputImg3_135_EXMPLR, OutputImg3_134_EXMPLR, 
      OutputImg3_133_EXMPLR, OutputImg3_132_EXMPLR, OutputImg3_131_EXMPLR, 
      OutputImg3_130_EXMPLR, OutputImg3_129_EXMPLR, OutputImg3_128_EXMPLR, 
      OutputImg3_127_EXMPLR, OutputImg3_126_EXMPLR, OutputImg3_125_EXMPLR, 
      OutputImg3_124_EXMPLR, OutputImg3_123_EXMPLR, OutputImg3_122_EXMPLR, 
      OutputImg3_121_EXMPLR, OutputImg3_120_EXMPLR, OutputImg3_119_EXMPLR, 
      OutputImg3_118_EXMPLR, OutputImg3_117_EXMPLR, OutputImg3_116_EXMPLR, 
      OutputImg3_115_EXMPLR, OutputImg3_114_EXMPLR, OutputImg3_113_EXMPLR, 
      OutputImg3_112_EXMPLR, OutputImg3_111_EXMPLR, OutputImg3_110_EXMPLR, 
      OutputImg3_109_EXMPLR, OutputImg3_108_EXMPLR, OutputImg3_107_EXMPLR, 
      OutputImg3_106_EXMPLR, OutputImg3_105_EXMPLR, OutputImg3_104_EXMPLR, 
      OutputImg3_103_EXMPLR, OutputImg3_102_EXMPLR, OutputImg3_101_EXMPLR, 
      OutputImg3_100_EXMPLR, OutputImg3_99_EXMPLR, OutputImg3_98_EXMPLR, 
      OutputImg3_97_EXMPLR, OutputImg3_96_EXMPLR, OutputImg3_95_EXMPLR, 
      OutputImg3_94_EXMPLR, OutputImg3_93_EXMPLR, OutputImg3_92_EXMPLR, 
      OutputImg3_91_EXMPLR, OutputImg3_90_EXMPLR, OutputImg3_89_EXMPLR, 
      OutputImg3_88_EXMPLR, OutputImg3_87_EXMPLR, OutputImg3_86_EXMPLR, 
      OutputImg3_85_EXMPLR, OutputImg3_84_EXMPLR, OutputImg3_83_EXMPLR, 
      OutputImg3_82_EXMPLR, OutputImg3_81_EXMPLR, OutputImg3_80_EXMPLR, 
      OutputImg3_79_EXMPLR, OutputImg3_78_EXMPLR, OutputImg3_77_EXMPLR, 
      OutputImg3_76_EXMPLR, OutputImg3_75_EXMPLR, OutputImg3_74_EXMPLR, 
      OutputImg3_73_EXMPLR, OutputImg3_72_EXMPLR, OutputImg3_71_EXMPLR, 
      OutputImg3_70_EXMPLR, OutputImg3_69_EXMPLR, OutputImg3_68_EXMPLR, 
      OutputImg3_67_EXMPLR, OutputImg3_66_EXMPLR, OutputImg3_65_EXMPLR, 
      OutputImg3_64_EXMPLR, OutputImg3_63_EXMPLR, OutputImg3_62_EXMPLR, 
      OutputImg3_61_EXMPLR, OutputImg3_60_EXMPLR, OutputImg3_59_EXMPLR, 
      OutputImg3_58_EXMPLR, OutputImg3_57_EXMPLR, OutputImg3_56_EXMPLR, 
      OutputImg3_55_EXMPLR, OutputImg3_54_EXMPLR, OutputImg3_53_EXMPLR, 
      OutputImg3_52_EXMPLR, OutputImg3_51_EXMPLR, OutputImg3_50_EXMPLR, 
      OutputImg3_49_EXMPLR, OutputImg3_48_EXMPLR, OutputImg3_47_EXMPLR, 
      OutputImg3_46_EXMPLR, OutputImg3_45_EXMPLR, OutputImg3_44_EXMPLR, 
      OutputImg3_43_EXMPLR, OutputImg3_42_EXMPLR, OutputImg3_41_EXMPLR, 
      OutputImg3_40_EXMPLR, OutputImg3_39_EXMPLR, OutputImg3_38_EXMPLR, 
      OutputImg3_37_EXMPLR, OutputImg3_36_EXMPLR, OutputImg3_35_EXMPLR, 
      OutputImg3_34_EXMPLR, OutputImg3_33_EXMPLR, OutputImg3_32_EXMPLR, 
      OutputImg3_31_EXMPLR, OutputImg3_30_EXMPLR, OutputImg3_29_EXMPLR, 
      OutputImg3_28_EXMPLR, OutputImg3_27_EXMPLR, OutputImg3_26_EXMPLR, 
      OutputImg3_25_EXMPLR, OutputImg3_24_EXMPLR, OutputImg3_23_EXMPLR, 
      OutputImg3_22_EXMPLR, OutputImg3_21_EXMPLR, OutputImg3_20_EXMPLR, 
      OutputImg3_19_EXMPLR, OutputImg3_18_EXMPLR, OutputImg3_17_EXMPLR, 
      OutputImg3_16_EXMPLR, OutputImg3_15_EXMPLR, OutputImg3_14_EXMPLR, 
      OutputImg3_13_EXMPLR, OutputImg3_12_EXMPLR, OutputImg3_11_EXMPLR, 
      OutputImg3_10_EXMPLR, OutputImg3_9_EXMPLR, OutputImg3_8_EXMPLR, 
      OutputImg3_7_EXMPLR, OutputImg3_6_EXMPLR, OutputImg3_5_EXMPLR, 
      OutputImg3_4_EXMPLR, OutputImg3_3_EXMPLR, OutputImg3_2_EXMPLR, 
      OutputImg3_1_EXMPLR, OutputImg3_0_EXMPLR, OutputImg4_447_EXMPLR, 
      OutputImg4_446_EXMPLR, OutputImg4_445_EXMPLR, OutputImg4_444_EXMPLR, 
      OutputImg4_443_EXMPLR, OutputImg4_442_EXMPLR, OutputImg4_441_EXMPLR, 
      OutputImg4_440_EXMPLR, OutputImg4_439_EXMPLR, OutputImg4_438_EXMPLR, 
      OutputImg4_437_EXMPLR, OutputImg4_436_EXMPLR, OutputImg4_435_EXMPLR, 
      OutputImg4_434_EXMPLR, OutputImg4_433_EXMPLR, OutputImg4_432_EXMPLR, 
      OutputImg4_431_EXMPLR, OutputImg4_430_EXMPLR, OutputImg4_429_EXMPLR, 
      OutputImg4_428_EXMPLR, OutputImg4_427_EXMPLR, OutputImg4_426_EXMPLR, 
      OutputImg4_425_EXMPLR, OutputImg4_424_EXMPLR, OutputImg4_423_EXMPLR, 
      OutputImg4_422_EXMPLR, OutputImg4_421_EXMPLR, OutputImg4_420_EXMPLR, 
      OutputImg4_419_EXMPLR, OutputImg4_418_EXMPLR, OutputImg4_417_EXMPLR, 
      OutputImg4_416_EXMPLR, OutputImg4_415_EXMPLR, OutputImg4_414_EXMPLR, 
      OutputImg4_413_EXMPLR, OutputImg4_412_EXMPLR, OutputImg4_411_EXMPLR, 
      OutputImg4_410_EXMPLR, OutputImg4_409_EXMPLR, OutputImg4_408_EXMPLR, 
      OutputImg4_407_EXMPLR, OutputImg4_406_EXMPLR, OutputImg4_405_EXMPLR, 
      OutputImg4_404_EXMPLR, OutputImg4_403_EXMPLR, OutputImg4_402_EXMPLR, 
      OutputImg4_401_EXMPLR, OutputImg4_400_EXMPLR, OutputImg4_399_EXMPLR, 
      OutputImg4_398_EXMPLR, OutputImg4_397_EXMPLR, OutputImg4_396_EXMPLR, 
      OutputImg4_395_EXMPLR, OutputImg4_394_EXMPLR, OutputImg4_393_EXMPLR, 
      OutputImg4_392_EXMPLR, OutputImg4_391_EXMPLR, OutputImg4_390_EXMPLR, 
      OutputImg4_389_EXMPLR, OutputImg4_388_EXMPLR, OutputImg4_387_EXMPLR, 
      OutputImg4_386_EXMPLR, OutputImg4_385_EXMPLR, OutputImg4_384_EXMPLR, 
      OutputImg4_383_EXMPLR, OutputImg4_382_EXMPLR, OutputImg4_381_EXMPLR, 
      OutputImg4_380_EXMPLR, OutputImg4_379_EXMPLR, OutputImg4_378_EXMPLR, 
      OutputImg4_377_EXMPLR, OutputImg4_376_EXMPLR, OutputImg4_375_EXMPLR, 
      OutputImg4_374_EXMPLR, OutputImg4_373_EXMPLR, OutputImg4_372_EXMPLR, 
      OutputImg4_371_EXMPLR, OutputImg4_370_EXMPLR, OutputImg4_369_EXMPLR, 
      OutputImg4_368_EXMPLR, OutputImg4_367_EXMPLR, OutputImg4_366_EXMPLR, 
      OutputImg4_365_EXMPLR, OutputImg4_364_EXMPLR, OutputImg4_363_EXMPLR, 
      OutputImg4_362_EXMPLR, OutputImg4_361_EXMPLR, OutputImg4_360_EXMPLR, 
      OutputImg4_359_EXMPLR, OutputImg4_358_EXMPLR, OutputImg4_357_EXMPLR, 
      OutputImg4_356_EXMPLR, OutputImg4_355_EXMPLR, OutputImg4_354_EXMPLR, 
      OutputImg4_353_EXMPLR, OutputImg4_352_EXMPLR, OutputImg4_351_EXMPLR, 
      OutputImg4_350_EXMPLR, OutputImg4_349_EXMPLR, OutputImg4_348_EXMPLR, 
      OutputImg4_347_EXMPLR, OutputImg4_346_EXMPLR, OutputImg4_345_EXMPLR, 
      OutputImg4_344_EXMPLR, OutputImg4_343_EXMPLR, OutputImg4_342_EXMPLR, 
      OutputImg4_341_EXMPLR, OutputImg4_340_EXMPLR, OutputImg4_339_EXMPLR, 
      OutputImg4_338_EXMPLR, OutputImg4_337_EXMPLR, OutputImg4_336_EXMPLR, 
      OutputImg4_335_EXMPLR, OutputImg4_334_EXMPLR, OutputImg4_333_EXMPLR, 
      OutputImg4_332_EXMPLR, OutputImg4_331_EXMPLR, OutputImg4_330_EXMPLR, 
      OutputImg4_329_EXMPLR, OutputImg4_328_EXMPLR, OutputImg4_327_EXMPLR, 
      OutputImg4_326_EXMPLR, OutputImg4_325_EXMPLR, OutputImg4_324_EXMPLR, 
      OutputImg4_323_EXMPLR, OutputImg4_322_EXMPLR, OutputImg4_321_EXMPLR, 
      OutputImg4_320_EXMPLR, OutputImg4_319_EXMPLR, OutputImg4_318_EXMPLR, 
      OutputImg4_317_EXMPLR, OutputImg4_316_EXMPLR, OutputImg4_315_EXMPLR, 
      OutputImg4_314_EXMPLR, OutputImg4_313_EXMPLR, OutputImg4_312_EXMPLR, 
      OutputImg4_311_EXMPLR, OutputImg4_310_EXMPLR, OutputImg4_309_EXMPLR, 
      OutputImg4_308_EXMPLR, OutputImg4_307_EXMPLR, OutputImg4_306_EXMPLR, 
      OutputImg4_305_EXMPLR, OutputImg4_304_EXMPLR, OutputImg4_303_EXMPLR, 
      OutputImg4_302_EXMPLR, OutputImg4_301_EXMPLR, OutputImg4_300_EXMPLR, 
      OutputImg4_299_EXMPLR, OutputImg4_298_EXMPLR, OutputImg4_297_EXMPLR, 
      OutputImg4_296_EXMPLR, OutputImg4_295_EXMPLR, OutputImg4_294_EXMPLR, 
      OutputImg4_293_EXMPLR, OutputImg4_292_EXMPLR, OutputImg4_291_EXMPLR, 
      OutputImg4_290_EXMPLR, OutputImg4_289_EXMPLR, OutputImg4_288_EXMPLR, 
      OutputImg4_287_EXMPLR, OutputImg4_286_EXMPLR, OutputImg4_285_EXMPLR, 
      OutputImg4_284_EXMPLR, OutputImg4_283_EXMPLR, OutputImg4_282_EXMPLR, 
      OutputImg4_281_EXMPLR, OutputImg4_280_EXMPLR, OutputImg4_279_EXMPLR, 
      OutputImg4_278_EXMPLR, OutputImg4_277_EXMPLR, OutputImg4_276_EXMPLR, 
      OutputImg4_275_EXMPLR, OutputImg4_274_EXMPLR, OutputImg4_273_EXMPLR, 
      OutputImg4_272_EXMPLR, OutputImg4_271_EXMPLR, OutputImg4_270_EXMPLR, 
      OutputImg4_269_EXMPLR, OutputImg4_268_EXMPLR, OutputImg4_267_EXMPLR, 
      OutputImg4_266_EXMPLR, OutputImg4_265_EXMPLR, OutputImg4_264_EXMPLR, 
      OutputImg4_263_EXMPLR, OutputImg4_262_EXMPLR, OutputImg4_261_EXMPLR, 
      OutputImg4_260_EXMPLR, OutputImg4_259_EXMPLR, OutputImg4_258_EXMPLR, 
      OutputImg4_257_EXMPLR, OutputImg4_256_EXMPLR, OutputImg4_255_EXMPLR, 
      OutputImg4_254_EXMPLR, OutputImg4_253_EXMPLR, OutputImg4_252_EXMPLR, 
      OutputImg4_251_EXMPLR, OutputImg4_250_EXMPLR, OutputImg4_249_EXMPLR, 
      OutputImg4_248_EXMPLR, OutputImg4_247_EXMPLR, OutputImg4_246_EXMPLR, 
      OutputImg4_245_EXMPLR, OutputImg4_244_EXMPLR, OutputImg4_243_EXMPLR, 
      OutputImg4_242_EXMPLR, OutputImg4_241_EXMPLR, OutputImg4_240_EXMPLR, 
      OutputImg4_239_EXMPLR, OutputImg4_238_EXMPLR, OutputImg4_237_EXMPLR, 
      OutputImg4_236_EXMPLR, OutputImg4_235_EXMPLR, OutputImg4_234_EXMPLR, 
      OutputImg4_233_EXMPLR, OutputImg4_232_EXMPLR, OutputImg4_231_EXMPLR, 
      OutputImg4_230_EXMPLR, OutputImg4_229_EXMPLR, OutputImg4_228_EXMPLR, 
      OutputImg4_227_EXMPLR, OutputImg4_226_EXMPLR, OutputImg4_225_EXMPLR, 
      OutputImg4_224_EXMPLR, OutputImg4_223_EXMPLR, OutputImg4_222_EXMPLR, 
      OutputImg4_221_EXMPLR, OutputImg4_220_EXMPLR, OutputImg4_219_EXMPLR, 
      OutputImg4_218_EXMPLR, OutputImg4_217_EXMPLR, OutputImg4_216_EXMPLR, 
      OutputImg4_215_EXMPLR, OutputImg4_214_EXMPLR, OutputImg4_213_EXMPLR, 
      OutputImg4_212_EXMPLR, OutputImg4_211_EXMPLR, OutputImg4_210_EXMPLR, 
      OutputImg4_209_EXMPLR, OutputImg4_208_EXMPLR, OutputImg4_207_EXMPLR, 
      OutputImg4_206_EXMPLR, OutputImg4_205_EXMPLR, OutputImg4_204_EXMPLR, 
      OutputImg4_203_EXMPLR, OutputImg4_202_EXMPLR, OutputImg4_201_EXMPLR, 
      OutputImg4_200_EXMPLR, OutputImg4_199_EXMPLR, OutputImg4_198_EXMPLR, 
      OutputImg4_197_EXMPLR, OutputImg4_196_EXMPLR, OutputImg4_195_EXMPLR, 
      OutputImg4_194_EXMPLR, OutputImg4_193_EXMPLR, OutputImg4_192_EXMPLR, 
      OutputImg4_191_EXMPLR, OutputImg4_190_EXMPLR, OutputImg4_189_EXMPLR, 
      OutputImg4_188_EXMPLR, OutputImg4_187_EXMPLR, OutputImg4_186_EXMPLR, 
      OutputImg4_185_EXMPLR, OutputImg4_184_EXMPLR, OutputImg4_183_EXMPLR, 
      OutputImg4_182_EXMPLR, OutputImg4_181_EXMPLR, OutputImg4_180_EXMPLR, 
      OutputImg4_179_EXMPLR, OutputImg4_178_EXMPLR, OutputImg4_177_EXMPLR, 
      OutputImg4_176_EXMPLR, OutputImg4_175_EXMPLR, OutputImg4_174_EXMPLR, 
      OutputImg4_173_EXMPLR, OutputImg4_172_EXMPLR, OutputImg4_171_EXMPLR, 
      OutputImg4_170_EXMPLR, OutputImg4_169_EXMPLR, OutputImg4_168_EXMPLR, 
      OutputImg4_167_EXMPLR, OutputImg4_166_EXMPLR, OutputImg4_165_EXMPLR, 
      OutputImg4_164_EXMPLR, OutputImg4_163_EXMPLR, OutputImg4_162_EXMPLR, 
      OutputImg4_161_EXMPLR, OutputImg4_160_EXMPLR, OutputImg4_159_EXMPLR, 
      OutputImg4_158_EXMPLR, OutputImg4_157_EXMPLR, OutputImg4_156_EXMPLR, 
      OutputImg4_155_EXMPLR, OutputImg4_154_EXMPLR, OutputImg4_153_EXMPLR, 
      OutputImg4_152_EXMPLR, OutputImg4_151_EXMPLR, OutputImg4_150_EXMPLR, 
      OutputImg4_149_EXMPLR, OutputImg4_148_EXMPLR, OutputImg4_147_EXMPLR, 
      OutputImg4_146_EXMPLR, OutputImg4_145_EXMPLR, OutputImg4_144_EXMPLR, 
      OutputImg4_143_EXMPLR, OutputImg4_142_EXMPLR, OutputImg4_141_EXMPLR, 
      OutputImg4_140_EXMPLR, OutputImg4_139_EXMPLR, OutputImg4_138_EXMPLR, 
      OutputImg4_137_EXMPLR, OutputImg4_136_EXMPLR, OutputImg4_135_EXMPLR, 
      OutputImg4_134_EXMPLR, OutputImg4_133_EXMPLR, OutputImg4_132_EXMPLR, 
      OutputImg4_131_EXMPLR, OutputImg4_130_EXMPLR, OutputImg4_129_EXMPLR, 
      OutputImg4_128_EXMPLR, OutputImg4_127_EXMPLR, OutputImg4_126_EXMPLR, 
      OutputImg4_125_EXMPLR, OutputImg4_124_EXMPLR, OutputImg4_123_EXMPLR, 
      OutputImg4_122_EXMPLR, OutputImg4_121_EXMPLR, OutputImg4_120_EXMPLR, 
      OutputImg4_119_EXMPLR, OutputImg4_118_EXMPLR, OutputImg4_117_EXMPLR, 
      OutputImg4_116_EXMPLR, OutputImg4_115_EXMPLR, OutputImg4_114_EXMPLR, 
      OutputImg4_113_EXMPLR, OutputImg4_112_EXMPLR, OutputImg4_111_EXMPLR, 
      OutputImg4_110_EXMPLR, OutputImg4_109_EXMPLR, OutputImg4_108_EXMPLR, 
      OutputImg4_107_EXMPLR, OutputImg4_106_EXMPLR, OutputImg4_105_EXMPLR, 
      OutputImg4_104_EXMPLR, OutputImg4_103_EXMPLR, OutputImg4_102_EXMPLR, 
      OutputImg4_101_EXMPLR, OutputImg4_100_EXMPLR, OutputImg4_99_EXMPLR, 
      OutputImg4_98_EXMPLR, OutputImg4_97_EXMPLR, OutputImg4_96_EXMPLR, 
      OutputImg4_95_EXMPLR, OutputImg4_94_EXMPLR, OutputImg4_93_EXMPLR, 
      OutputImg4_92_EXMPLR, OutputImg4_91_EXMPLR, OutputImg4_90_EXMPLR, 
      OutputImg4_89_EXMPLR, OutputImg4_88_EXMPLR, OutputImg4_87_EXMPLR, 
      OutputImg4_86_EXMPLR, OutputImg4_85_EXMPLR, OutputImg4_84_EXMPLR, 
      OutputImg4_83_EXMPLR, OutputImg4_82_EXMPLR, OutputImg4_81_EXMPLR, 
      OutputImg4_80_EXMPLR, OutputImg4_79_EXMPLR, OutputImg4_78_EXMPLR, 
      OutputImg4_77_EXMPLR, OutputImg4_76_EXMPLR, OutputImg4_75_EXMPLR, 
      OutputImg4_74_EXMPLR, OutputImg4_73_EXMPLR, OutputImg4_72_EXMPLR, 
      OutputImg4_71_EXMPLR, OutputImg4_70_EXMPLR, OutputImg4_69_EXMPLR, 
      OutputImg4_68_EXMPLR, OutputImg4_67_EXMPLR, OutputImg4_66_EXMPLR, 
      OutputImg4_65_EXMPLR, OutputImg4_64_EXMPLR, OutputImg4_63_EXMPLR, 
      OutputImg4_62_EXMPLR, OutputImg4_61_EXMPLR, OutputImg4_60_EXMPLR, 
      OutputImg4_59_EXMPLR, OutputImg4_58_EXMPLR, OutputImg4_57_EXMPLR, 
      OutputImg4_56_EXMPLR, OutputImg4_55_EXMPLR, OutputImg4_54_EXMPLR, 
      OutputImg4_53_EXMPLR, OutputImg4_52_EXMPLR, OutputImg4_51_EXMPLR, 
      OutputImg4_50_EXMPLR, OutputImg4_49_EXMPLR, OutputImg4_48_EXMPLR, 
      OutputImg4_47_EXMPLR, OutputImg4_46_EXMPLR, OutputImg4_45_EXMPLR, 
      OutputImg4_44_EXMPLR, OutputImg4_43_EXMPLR, OutputImg4_42_EXMPLR, 
      OutputImg4_41_EXMPLR, OutputImg4_40_EXMPLR, OutputImg4_39_EXMPLR, 
      OutputImg4_38_EXMPLR, OutputImg4_37_EXMPLR, OutputImg4_36_EXMPLR, 
      OutputImg4_35_EXMPLR, OutputImg4_34_EXMPLR, OutputImg4_33_EXMPLR, 
      OutputImg4_32_EXMPLR, OutputImg4_31_EXMPLR, OutputImg4_30_EXMPLR, 
      OutputImg4_29_EXMPLR, OutputImg4_28_EXMPLR, OutputImg4_27_EXMPLR, 
      OutputImg4_26_EXMPLR, OutputImg4_25_EXMPLR, OutputImg4_24_EXMPLR, 
      OutputImg4_23_EXMPLR, OutputImg4_22_EXMPLR, OutputImg4_21_EXMPLR, 
      OutputImg4_20_EXMPLR, OutputImg4_19_EXMPLR, OutputImg4_18_EXMPLR, 
      OutputImg4_17_EXMPLR, OutputImg4_16_EXMPLR, OutputImg4_15_EXMPLR, 
      OutputImg4_14_EXMPLR, OutputImg4_13_EXMPLR, OutputImg4_12_EXMPLR, 
      OutputImg4_11_EXMPLR, OutputImg4_10_EXMPLR, OutputImg4_9_EXMPLR, 
      OutputImg4_8_EXMPLR, OutputImg4_7_EXMPLR, OutputImg4_6_EXMPLR, 
      OutputImg4_5_EXMPLR, OutputImg4_4_EXMPLR, OutputImg4_3_EXMPLR, 
      OutputImg4_2_EXMPLR, OutputImg4_1_EXMPLR, OutputImg4_0_EXMPLR, 
      OutputImg5_447_EXMPLR, OutputImg5_446_EXMPLR, OutputImg5_445_EXMPLR, 
      OutputImg5_444_EXMPLR, OutputImg5_443_EXMPLR, OutputImg5_442_EXMPLR, 
      OutputImg5_441_EXMPLR, OutputImg5_440_EXMPLR, OutputImg5_439_EXMPLR, 
      OutputImg5_438_EXMPLR, OutputImg5_437_EXMPLR, OutputImg5_436_EXMPLR, 
      OutputImg5_435_EXMPLR, OutputImg5_434_EXMPLR, OutputImg5_433_EXMPLR, 
      OutputImg5_432_EXMPLR, OutputImg5_431_EXMPLR, OutputImg5_430_EXMPLR, 
      OutputImg5_429_EXMPLR, OutputImg5_428_EXMPLR, OutputImg5_427_EXMPLR, 
      OutputImg5_426_EXMPLR, OutputImg5_425_EXMPLR, OutputImg5_424_EXMPLR, 
      OutputImg5_423_EXMPLR, OutputImg5_422_EXMPLR, OutputImg5_421_EXMPLR, 
      OutputImg5_420_EXMPLR, OutputImg5_419_EXMPLR, OutputImg5_418_EXMPLR, 
      OutputImg5_417_EXMPLR, OutputImg5_416_EXMPLR, OutputImg5_415_EXMPLR, 
      OutputImg5_414_EXMPLR, OutputImg5_413_EXMPLR, OutputImg5_412_EXMPLR, 
      OutputImg5_411_EXMPLR, OutputImg5_410_EXMPLR, OutputImg5_409_EXMPLR, 
      OutputImg5_408_EXMPLR, OutputImg5_407_EXMPLR, OutputImg5_406_EXMPLR, 
      OutputImg5_405_EXMPLR, OutputImg5_404_EXMPLR, OutputImg5_403_EXMPLR, 
      OutputImg5_402_EXMPLR, OutputImg5_401_EXMPLR, OutputImg5_400_EXMPLR, 
      OutputImg5_399_EXMPLR, OutputImg5_398_EXMPLR, OutputImg5_397_EXMPLR, 
      OutputImg5_396_EXMPLR, OutputImg5_395_EXMPLR, OutputImg5_394_EXMPLR, 
      OutputImg5_393_EXMPLR, OutputImg5_392_EXMPLR, OutputImg5_391_EXMPLR, 
      OutputImg5_390_EXMPLR, OutputImg5_389_EXMPLR, OutputImg5_388_EXMPLR, 
      OutputImg5_387_EXMPLR, OutputImg5_386_EXMPLR, OutputImg5_385_EXMPLR, 
      OutputImg5_384_EXMPLR, OutputImg5_383_EXMPLR, OutputImg5_382_EXMPLR, 
      OutputImg5_381_EXMPLR, OutputImg5_380_EXMPLR, OutputImg5_379_EXMPLR, 
      OutputImg5_378_EXMPLR, OutputImg5_377_EXMPLR, OutputImg5_376_EXMPLR, 
      OutputImg5_375_EXMPLR, OutputImg5_374_EXMPLR, OutputImg5_373_EXMPLR, 
      OutputImg5_372_EXMPLR, OutputImg5_371_EXMPLR, OutputImg5_370_EXMPLR, 
      OutputImg5_369_EXMPLR, OutputImg5_368_EXMPLR, OutputImg5_367_EXMPLR, 
      OutputImg5_366_EXMPLR, OutputImg5_365_EXMPLR, OutputImg5_364_EXMPLR, 
      OutputImg5_363_EXMPLR, OutputImg5_362_EXMPLR, OutputImg5_361_EXMPLR, 
      OutputImg5_360_EXMPLR, OutputImg5_359_EXMPLR, OutputImg5_358_EXMPLR, 
      OutputImg5_357_EXMPLR, OutputImg5_356_EXMPLR, OutputImg5_355_EXMPLR, 
      OutputImg5_354_EXMPLR, OutputImg5_353_EXMPLR, OutputImg5_352_EXMPLR, 
      OutputImg5_351_EXMPLR, OutputImg5_350_EXMPLR, OutputImg5_349_EXMPLR, 
      OutputImg5_348_EXMPLR, OutputImg5_347_EXMPLR, OutputImg5_346_EXMPLR, 
      OutputImg5_345_EXMPLR, OutputImg5_344_EXMPLR, OutputImg5_343_EXMPLR, 
      OutputImg5_342_EXMPLR, OutputImg5_341_EXMPLR, OutputImg5_340_EXMPLR, 
      OutputImg5_339_EXMPLR, OutputImg5_338_EXMPLR, OutputImg5_337_EXMPLR, 
      OutputImg5_336_EXMPLR, OutputImg5_335_EXMPLR, OutputImg5_334_EXMPLR, 
      OutputImg5_333_EXMPLR, OutputImg5_332_EXMPLR, OutputImg5_331_EXMPLR, 
      OutputImg5_330_EXMPLR, OutputImg5_329_EXMPLR, OutputImg5_328_EXMPLR, 
      OutputImg5_327_EXMPLR, OutputImg5_326_EXMPLR, OutputImg5_325_EXMPLR, 
      OutputImg5_324_EXMPLR, OutputImg5_323_EXMPLR, OutputImg5_322_EXMPLR, 
      OutputImg5_321_EXMPLR, OutputImg5_320_EXMPLR, OutputImg5_319_EXMPLR, 
      OutputImg5_318_EXMPLR, OutputImg5_317_EXMPLR, OutputImg5_316_EXMPLR, 
      OutputImg5_315_EXMPLR, OutputImg5_314_EXMPLR, OutputImg5_313_EXMPLR, 
      OutputImg5_312_EXMPLR, OutputImg5_311_EXMPLR, OutputImg5_310_EXMPLR, 
      OutputImg5_309_EXMPLR, OutputImg5_308_EXMPLR, OutputImg5_307_EXMPLR, 
      OutputImg5_306_EXMPLR, OutputImg5_305_EXMPLR, OutputImg5_304_EXMPLR, 
      OutputImg5_303_EXMPLR, OutputImg5_302_EXMPLR, OutputImg5_301_EXMPLR, 
      OutputImg5_300_EXMPLR, OutputImg5_299_EXMPLR, OutputImg5_298_EXMPLR, 
      OutputImg5_297_EXMPLR, OutputImg5_296_EXMPLR, OutputImg5_295_EXMPLR, 
      OutputImg5_294_EXMPLR, OutputImg5_293_EXMPLR, OutputImg5_292_EXMPLR, 
      OutputImg5_291_EXMPLR, OutputImg5_290_EXMPLR, OutputImg5_289_EXMPLR, 
      OutputImg5_288_EXMPLR, OutputImg5_287_EXMPLR, OutputImg5_286_EXMPLR, 
      OutputImg5_285_EXMPLR, OutputImg5_284_EXMPLR, OutputImg5_283_EXMPLR, 
      OutputImg5_282_EXMPLR, OutputImg5_281_EXMPLR, OutputImg5_280_EXMPLR, 
      OutputImg5_279_EXMPLR, OutputImg5_278_EXMPLR, OutputImg5_277_EXMPLR, 
      OutputImg5_276_EXMPLR, OutputImg5_275_EXMPLR, OutputImg5_274_EXMPLR, 
      OutputImg5_273_EXMPLR, OutputImg5_272_EXMPLR, OutputImg5_271_EXMPLR, 
      OutputImg5_270_EXMPLR, OutputImg5_269_EXMPLR, OutputImg5_268_EXMPLR, 
      OutputImg5_267_EXMPLR, OutputImg5_266_EXMPLR, OutputImg5_265_EXMPLR, 
      OutputImg5_264_EXMPLR, OutputImg5_263_EXMPLR, OutputImg5_262_EXMPLR, 
      OutputImg5_261_EXMPLR, OutputImg5_260_EXMPLR, OutputImg5_259_EXMPLR, 
      OutputImg5_258_EXMPLR, OutputImg5_257_EXMPLR, OutputImg5_256_EXMPLR, 
      OutputImg5_255_EXMPLR, OutputImg5_254_EXMPLR, OutputImg5_253_EXMPLR, 
      OutputImg5_252_EXMPLR, OutputImg5_251_EXMPLR, OutputImg5_250_EXMPLR, 
      OutputImg5_249_EXMPLR, OutputImg5_248_EXMPLR, OutputImg5_247_EXMPLR, 
      OutputImg5_246_EXMPLR, OutputImg5_245_EXMPLR, OutputImg5_244_EXMPLR, 
      OutputImg5_243_EXMPLR, OutputImg5_242_EXMPLR, OutputImg5_241_EXMPLR, 
      OutputImg5_240_EXMPLR, OutputImg5_239_EXMPLR, OutputImg5_238_EXMPLR, 
      OutputImg5_237_EXMPLR, OutputImg5_236_EXMPLR, OutputImg5_235_EXMPLR, 
      OutputImg5_234_EXMPLR, OutputImg5_233_EXMPLR, OutputImg5_232_EXMPLR, 
      OutputImg5_231_EXMPLR, OutputImg5_230_EXMPLR, OutputImg5_229_EXMPLR, 
      OutputImg5_228_EXMPLR, OutputImg5_227_EXMPLR, OutputImg5_226_EXMPLR, 
      OutputImg5_225_EXMPLR, OutputImg5_224_EXMPLR, OutputImg5_223_EXMPLR, 
      OutputImg5_222_EXMPLR, OutputImg5_221_EXMPLR, OutputImg5_220_EXMPLR, 
      OutputImg5_219_EXMPLR, OutputImg5_218_EXMPLR, OutputImg5_217_EXMPLR, 
      OutputImg5_216_EXMPLR, OutputImg5_215_EXMPLR, OutputImg5_214_EXMPLR, 
      OutputImg5_213_EXMPLR, OutputImg5_212_EXMPLR, OutputImg5_211_EXMPLR, 
      OutputImg5_210_EXMPLR, OutputImg5_209_EXMPLR, OutputImg5_208_EXMPLR, 
      OutputImg5_207_EXMPLR, OutputImg5_206_EXMPLR, OutputImg5_205_EXMPLR, 
      OutputImg5_204_EXMPLR, OutputImg5_203_EXMPLR, OutputImg5_202_EXMPLR, 
      OutputImg5_201_EXMPLR, OutputImg5_200_EXMPLR, OutputImg5_199_EXMPLR, 
      OutputImg5_198_EXMPLR, OutputImg5_197_EXMPLR, OutputImg5_196_EXMPLR, 
      OutputImg5_195_EXMPLR, OutputImg5_194_EXMPLR, OutputImg5_193_EXMPLR, 
      OutputImg5_192_EXMPLR, OutputImg5_191_EXMPLR, OutputImg5_190_EXMPLR, 
      OutputImg5_189_EXMPLR, OutputImg5_188_EXMPLR, OutputImg5_187_EXMPLR, 
      OutputImg5_186_EXMPLR, OutputImg5_185_EXMPLR, OutputImg5_184_EXMPLR, 
      OutputImg5_183_EXMPLR, OutputImg5_182_EXMPLR, OutputImg5_181_EXMPLR, 
      OutputImg5_180_EXMPLR, OutputImg5_179_EXMPLR, OutputImg5_178_EXMPLR, 
      OutputImg5_177_EXMPLR, OutputImg5_176_EXMPLR, OutputImg5_175_EXMPLR, 
      OutputImg5_174_EXMPLR, OutputImg5_173_EXMPLR, OutputImg5_172_EXMPLR, 
      OutputImg5_171_EXMPLR, OutputImg5_170_EXMPLR, OutputImg5_169_EXMPLR, 
      OutputImg5_168_EXMPLR, OutputImg5_167_EXMPLR, OutputImg5_166_EXMPLR, 
      OutputImg5_165_EXMPLR, OutputImg5_164_EXMPLR, OutputImg5_163_EXMPLR, 
      OutputImg5_162_EXMPLR, OutputImg5_161_EXMPLR, OutputImg5_160_EXMPLR, 
      OutputImg5_159_EXMPLR, OutputImg5_158_EXMPLR, OutputImg5_157_EXMPLR, 
      OutputImg5_156_EXMPLR, OutputImg5_155_EXMPLR, OutputImg5_154_EXMPLR, 
      OutputImg5_153_EXMPLR, OutputImg5_152_EXMPLR, OutputImg5_151_EXMPLR, 
      OutputImg5_150_EXMPLR, OutputImg5_149_EXMPLR, OutputImg5_148_EXMPLR, 
      OutputImg5_147_EXMPLR, OutputImg5_146_EXMPLR, OutputImg5_145_EXMPLR, 
      OutputImg5_144_EXMPLR, OutputImg5_143_EXMPLR, OutputImg5_142_EXMPLR, 
      OutputImg5_141_EXMPLR, OutputImg5_140_EXMPLR, OutputImg5_139_EXMPLR, 
      OutputImg5_138_EXMPLR, OutputImg5_137_EXMPLR, OutputImg5_136_EXMPLR, 
      OutputImg5_135_EXMPLR, OutputImg5_134_EXMPLR, OutputImg5_133_EXMPLR, 
      OutputImg5_132_EXMPLR, OutputImg5_131_EXMPLR, OutputImg5_130_EXMPLR, 
      OutputImg5_129_EXMPLR, OutputImg5_128_EXMPLR, OutputImg5_127_EXMPLR, 
      OutputImg5_126_EXMPLR, OutputImg5_125_EXMPLR, OutputImg5_124_EXMPLR, 
      OutputImg5_123_EXMPLR, OutputImg5_122_EXMPLR, OutputImg5_121_EXMPLR, 
      OutputImg5_120_EXMPLR, OutputImg5_119_EXMPLR, OutputImg5_118_EXMPLR, 
      OutputImg5_117_EXMPLR, OutputImg5_116_EXMPLR, OutputImg5_115_EXMPLR, 
      OutputImg5_114_EXMPLR, OutputImg5_113_EXMPLR, OutputImg5_112_EXMPLR, 
      OutputImg5_111_EXMPLR, OutputImg5_110_EXMPLR, OutputImg5_109_EXMPLR, 
      OutputImg5_108_EXMPLR, OutputImg5_107_EXMPLR, OutputImg5_106_EXMPLR, 
      OutputImg5_105_EXMPLR, OutputImg5_104_EXMPLR, OutputImg5_103_EXMPLR, 
      OutputImg5_102_EXMPLR, OutputImg5_101_EXMPLR, OutputImg5_100_EXMPLR, 
      OutputImg5_99_EXMPLR, OutputImg5_98_EXMPLR, OutputImg5_97_EXMPLR, 
      OutputImg5_96_EXMPLR, OutputImg5_95_EXMPLR, OutputImg5_94_EXMPLR, 
      OutputImg5_93_EXMPLR, OutputImg5_92_EXMPLR, OutputImg5_91_EXMPLR, 
      OutputImg5_90_EXMPLR, OutputImg5_89_EXMPLR, OutputImg5_88_EXMPLR, 
      OutputImg5_87_EXMPLR, OutputImg5_86_EXMPLR, OutputImg5_85_EXMPLR, 
      OutputImg5_84_EXMPLR, OutputImg5_83_EXMPLR, OutputImg5_82_EXMPLR, 
      OutputImg5_81_EXMPLR, OutputImg5_80_EXMPLR, OutputImg5_79_EXMPLR, 
      OutputImg5_78_EXMPLR, OutputImg5_77_EXMPLR, OutputImg5_76_EXMPLR, 
      OutputImg5_75_EXMPLR, OutputImg5_74_EXMPLR, OutputImg5_73_EXMPLR, 
      OutputImg5_72_EXMPLR, OutputImg5_71_EXMPLR, OutputImg5_70_EXMPLR, 
      OutputImg5_69_EXMPLR, OutputImg5_68_EXMPLR, OutputImg5_67_EXMPLR, 
      OutputImg5_66_EXMPLR, OutputImg5_65_EXMPLR, OutputImg5_64_EXMPLR, 
      OutputImg5_63_EXMPLR, OutputImg5_62_EXMPLR, OutputImg5_61_EXMPLR, 
      OutputImg5_60_EXMPLR, OutputImg5_59_EXMPLR, OutputImg5_58_EXMPLR, 
      OutputImg5_57_EXMPLR, OutputImg5_56_EXMPLR, OutputImg5_55_EXMPLR, 
      OutputImg5_54_EXMPLR, OutputImg5_53_EXMPLR, OutputImg5_52_EXMPLR, 
      OutputImg5_51_EXMPLR, OutputImg5_50_EXMPLR, OutputImg5_49_EXMPLR, 
      OutputImg5_48_EXMPLR, OutputImg5_47_EXMPLR, OutputImg5_46_EXMPLR, 
      OutputImg5_45_EXMPLR, OutputImg5_44_EXMPLR, OutputImg5_43_EXMPLR, 
      OutputImg5_42_EXMPLR, OutputImg5_41_EXMPLR, OutputImg5_40_EXMPLR, 
      OutputImg5_39_EXMPLR, OutputImg5_38_EXMPLR, OutputImg5_37_EXMPLR, 
      OutputImg5_36_EXMPLR, OutputImg5_35_EXMPLR, OutputImg5_34_EXMPLR, 
      OutputImg5_33_EXMPLR, OutputImg5_32_EXMPLR, OutputImg5_31_EXMPLR, 
      OutputImg5_30_EXMPLR, OutputImg5_29_EXMPLR, OutputImg5_28_EXMPLR, 
      OutputImg5_27_EXMPLR, OutputImg5_26_EXMPLR, OutputImg5_25_EXMPLR, 
      OutputImg5_24_EXMPLR, OutputImg5_23_EXMPLR, OutputImg5_22_EXMPLR, 
      OutputImg5_21_EXMPLR, OutputImg5_20_EXMPLR, OutputImg5_19_EXMPLR, 
      OutputImg5_18_EXMPLR, OutputImg5_17_EXMPLR, OutputImg5_16_EXMPLR, 
      OutputImg5_15_EXMPLR, OutputImg5_14_EXMPLR, OutputImg5_13_EXMPLR, 
      OutputImg5_12_EXMPLR, OutputImg5_11_EXMPLR, OutputImg5_10_EXMPLR, 
      OutputImg5_9_EXMPLR, OutputImg5_8_EXMPLR, OutputImg5_7_EXMPLR, 
      OutputImg5_6_EXMPLR, OutputImg5_5_EXMPLR, OutputImg5_4_EXMPLR, 
      OutputImg5_3_EXMPLR, OutputImg5_2_EXMPLR, OutputImg5_1_EXMPLR, 
      OutputImg5_0_EXMPLR, ImgCounterOuput_2_EXMPLR, 
      ImgCounterOuput_1_EXMPLR, ImgCounterOuput_0_EXMPLR, ImgIndic_0_EXMPLR, 
      ImgEn_5_EXMPLR, ImgEn_4_EXMPLR, ImgEn_3_EXMPLR, ImgEn_2_EXMPLR, 
      ImgEn_1_EXMPLR, ImgEn_0_EXMPLR, newAdd16_12, newAdd16_11, newAdd16_10, 
      newAdd16_9, newAdd16_8, newAdd16_7, newAdd16_6, newAdd16_5, newAdd16_4, 
      newAdd16_3, newAdd16_2, newAdd16_1, newAdd16_0, DFFCLK, DecOutput_5, 
      DecOutput_4, DecOutput_3, DecOutput_2, DecOutput_1, DecOutput_0, 
      ImgReg0IN_447, ImgReg0IN_446, ImgReg0IN_445, ImgReg0IN_444, 
      ImgReg0IN_443, ImgReg0IN_442, ImgReg0IN_441, ImgReg0IN_440, 
      ImgReg0IN_439, ImgReg0IN_438, ImgReg0IN_437, ImgReg0IN_436, 
      ImgReg0IN_435, ImgReg0IN_434, ImgReg0IN_433, ImgReg0IN_432, 
      ImgReg0IN_431, ImgReg0IN_430, ImgReg0IN_429, ImgReg0IN_428, 
      ImgReg0IN_427, ImgReg0IN_426, ImgReg0IN_425, ImgReg0IN_424, 
      ImgReg0IN_423, ImgReg0IN_422, ImgReg0IN_421, ImgReg0IN_420, 
      ImgReg0IN_419, ImgReg0IN_418, ImgReg0IN_417, ImgReg0IN_416, 
      ImgReg0IN_415, ImgReg0IN_414, ImgReg0IN_413, ImgReg0IN_412, 
      ImgReg0IN_411, ImgReg0IN_410, ImgReg0IN_409, ImgReg0IN_408, 
      ImgReg0IN_407, ImgReg0IN_406, ImgReg0IN_405, ImgReg0IN_404, 
      ImgReg0IN_403, ImgReg0IN_402, ImgReg0IN_401, ImgReg0IN_400, 
      ImgReg0IN_399, ImgReg0IN_398, ImgReg0IN_397, ImgReg0IN_396, 
      ImgReg0IN_395, ImgReg0IN_394, ImgReg0IN_393, ImgReg0IN_392, 
      ImgReg0IN_391, ImgReg0IN_390, ImgReg0IN_389, ImgReg0IN_388, 
      ImgReg0IN_387, ImgReg0IN_386, ImgReg0IN_385, ImgReg0IN_384, 
      ImgReg0IN_383, ImgReg0IN_382, ImgReg0IN_381, ImgReg0IN_380, 
      ImgReg0IN_379, ImgReg0IN_378, ImgReg0IN_377, ImgReg0IN_376, 
      ImgReg0IN_375, ImgReg0IN_374, ImgReg0IN_373, ImgReg0IN_372, 
      ImgReg0IN_371, ImgReg0IN_370, ImgReg0IN_369, ImgReg0IN_368, 
      ImgReg0IN_367, ImgReg0IN_366, ImgReg0IN_365, ImgReg0IN_364, 
      ImgReg0IN_363, ImgReg0IN_362, ImgReg0IN_361, ImgReg0IN_360, 
      ImgReg0IN_359, ImgReg0IN_358, ImgReg0IN_357, ImgReg0IN_356, 
      ImgReg0IN_355, ImgReg0IN_354, ImgReg0IN_353, ImgReg0IN_352, 
      ImgReg0IN_351, ImgReg0IN_350, ImgReg0IN_349, ImgReg0IN_348, 
      ImgReg0IN_347, ImgReg0IN_346, ImgReg0IN_345, ImgReg0IN_344, 
      ImgReg0IN_343, ImgReg0IN_342, ImgReg0IN_341, ImgReg0IN_340, 
      ImgReg0IN_339, ImgReg0IN_338, ImgReg0IN_337, ImgReg0IN_336, 
      ImgReg0IN_335, ImgReg0IN_334, ImgReg0IN_333, ImgReg0IN_332, 
      ImgReg0IN_331, ImgReg0IN_330, ImgReg0IN_329, ImgReg0IN_328, 
      ImgReg0IN_327, ImgReg0IN_326, ImgReg0IN_325, ImgReg0IN_324, 
      ImgReg0IN_323, ImgReg0IN_322, ImgReg0IN_321, ImgReg0IN_320, 
      ImgReg0IN_319, ImgReg0IN_318, ImgReg0IN_317, ImgReg0IN_316, 
      ImgReg0IN_315, ImgReg0IN_314, ImgReg0IN_313, ImgReg0IN_312, 
      ImgReg0IN_311, ImgReg0IN_310, ImgReg0IN_309, ImgReg0IN_308, 
      ImgReg0IN_307, ImgReg0IN_306, ImgReg0IN_305, ImgReg0IN_304, 
      ImgReg0IN_303, ImgReg0IN_302, ImgReg0IN_301, ImgReg0IN_300, 
      ImgReg0IN_299, ImgReg0IN_298, ImgReg0IN_297, ImgReg0IN_296, 
      ImgReg0IN_295, ImgReg0IN_294, ImgReg0IN_293, ImgReg0IN_292, 
      ImgReg0IN_291, ImgReg0IN_290, ImgReg0IN_289, ImgReg0IN_288, 
      ImgReg0IN_287, ImgReg0IN_286, ImgReg0IN_285, ImgReg0IN_284, 
      ImgReg0IN_283, ImgReg0IN_282, ImgReg0IN_281, ImgReg0IN_280, 
      ImgReg0IN_279, ImgReg0IN_278, ImgReg0IN_277, ImgReg0IN_276, 
      ImgReg0IN_275, ImgReg0IN_274, ImgReg0IN_273, ImgReg0IN_272, 
      ImgReg0IN_271, ImgReg0IN_270, ImgReg0IN_269, ImgReg0IN_268, 
      ImgReg0IN_267, ImgReg0IN_266, ImgReg0IN_265, ImgReg0IN_264, 
      ImgReg0IN_263, ImgReg0IN_262, ImgReg0IN_261, ImgReg0IN_260, 
      ImgReg0IN_259, ImgReg0IN_258, ImgReg0IN_257, ImgReg0IN_256, 
      ImgReg0IN_255, ImgReg0IN_254, ImgReg0IN_253, ImgReg0IN_252, 
      ImgReg0IN_251, ImgReg0IN_250, ImgReg0IN_249, ImgReg0IN_248, 
      ImgReg0IN_247, ImgReg0IN_246, ImgReg0IN_245, ImgReg0IN_244, 
      ImgReg0IN_243, ImgReg0IN_242, ImgReg0IN_241, ImgReg0IN_240, 
      ImgReg0IN_239, ImgReg0IN_238, ImgReg0IN_237, ImgReg0IN_236, 
      ImgReg0IN_235, ImgReg0IN_234, ImgReg0IN_233, ImgReg0IN_232, 
      ImgReg0IN_231, ImgReg0IN_230, ImgReg0IN_229, ImgReg0IN_228, 
      ImgReg0IN_227, ImgReg0IN_226, ImgReg0IN_225, ImgReg0IN_224, 
      ImgReg0IN_223, ImgReg0IN_222, ImgReg0IN_221, ImgReg0IN_220, 
      ImgReg0IN_219, ImgReg0IN_218, ImgReg0IN_217, ImgReg0IN_216, 
      ImgReg0IN_215, ImgReg0IN_214, ImgReg0IN_213, ImgReg0IN_212, 
      ImgReg0IN_211, ImgReg0IN_210, ImgReg0IN_209, ImgReg0IN_208, 
      ImgReg0IN_207, ImgReg0IN_206, ImgReg0IN_205, ImgReg0IN_204, 
      ImgReg0IN_203, ImgReg0IN_202, ImgReg0IN_201, ImgReg0IN_200, 
      ImgReg0IN_199, ImgReg0IN_198, ImgReg0IN_197, ImgReg0IN_196, 
      ImgReg0IN_195, ImgReg0IN_194, ImgReg0IN_193, ImgReg0IN_192, 
      ImgReg0IN_191, ImgReg0IN_190, ImgReg0IN_189, ImgReg0IN_188, 
      ImgReg0IN_187, ImgReg0IN_186, ImgReg0IN_185, ImgReg0IN_184, 
      ImgReg0IN_183, ImgReg0IN_182, ImgReg0IN_181, ImgReg0IN_180, 
      ImgReg0IN_179, ImgReg0IN_178, ImgReg0IN_177, ImgReg0IN_176, 
      ImgReg0IN_175, ImgReg0IN_174, ImgReg0IN_173, ImgReg0IN_172, 
      ImgReg0IN_171, ImgReg0IN_170, ImgReg0IN_169, ImgReg0IN_168, 
      ImgReg0IN_167, ImgReg0IN_166, ImgReg0IN_165, ImgReg0IN_164, 
      ImgReg0IN_163, ImgReg0IN_162, ImgReg0IN_161, ImgReg0IN_160, 
      ImgReg0IN_159, ImgReg0IN_158, ImgReg0IN_157, ImgReg0IN_156, 
      ImgReg0IN_155, ImgReg0IN_154, ImgReg0IN_153, ImgReg0IN_152, 
      ImgReg0IN_151, ImgReg0IN_150, ImgReg0IN_149, ImgReg0IN_148, 
      ImgReg0IN_147, ImgReg0IN_146, ImgReg0IN_145, ImgReg0IN_144, 
      ImgReg0IN_143, ImgReg0IN_142, ImgReg0IN_141, ImgReg0IN_140, 
      ImgReg0IN_139, ImgReg0IN_138, ImgReg0IN_137, ImgReg0IN_136, 
      ImgReg0IN_135, ImgReg0IN_134, ImgReg0IN_133, ImgReg0IN_132, 
      ImgReg0IN_131, ImgReg0IN_130, ImgReg0IN_129, ImgReg0IN_128, 
      ImgReg0IN_127, ImgReg0IN_126, ImgReg0IN_125, ImgReg0IN_124, 
      ImgReg0IN_123, ImgReg0IN_122, ImgReg0IN_121, ImgReg0IN_120, 
      ImgReg0IN_119, ImgReg0IN_118, ImgReg0IN_117, ImgReg0IN_116, 
      ImgReg0IN_115, ImgReg0IN_114, ImgReg0IN_113, ImgReg0IN_112, 
      ImgReg0IN_111, ImgReg0IN_110, ImgReg0IN_109, ImgReg0IN_108, 
      ImgReg0IN_107, ImgReg0IN_106, ImgReg0IN_105, ImgReg0IN_104, 
      ImgReg0IN_103, ImgReg0IN_102, ImgReg0IN_101, ImgReg0IN_100, 
      ImgReg0IN_99, ImgReg0IN_98, ImgReg0IN_97, ImgReg0IN_96, ImgReg0IN_95, 
      ImgReg0IN_94, ImgReg0IN_93, ImgReg0IN_92, ImgReg0IN_91, ImgReg0IN_90, 
      ImgReg0IN_89, ImgReg0IN_88, ImgReg0IN_87, ImgReg0IN_86, ImgReg0IN_85, 
      ImgReg0IN_84, ImgReg0IN_83, ImgReg0IN_82, ImgReg0IN_81, ImgReg0IN_80, 
      ImgReg0IN_79, ImgReg0IN_78, ImgReg0IN_77, ImgReg0IN_76, ImgReg0IN_75, 
      ImgReg0IN_74, ImgReg0IN_73, ImgReg0IN_72, ImgReg0IN_71, ImgReg0IN_70, 
      ImgReg0IN_69, ImgReg0IN_68, ImgReg0IN_67, ImgReg0IN_66, ImgReg0IN_65, 
      ImgReg0IN_64, ImgReg0IN_63, ImgReg0IN_62, ImgReg0IN_61, ImgReg0IN_60, 
      ImgReg0IN_59, ImgReg0IN_58, ImgReg0IN_57, ImgReg0IN_56, ImgReg0IN_55, 
      ImgReg0IN_54, ImgReg0IN_53, ImgReg0IN_52, ImgReg0IN_51, ImgReg0IN_50, 
      ImgReg0IN_49, ImgReg0IN_48, ImgReg0IN_47, ImgReg0IN_46, ImgReg0IN_45, 
      ImgReg0IN_44, ImgReg0IN_43, ImgReg0IN_42, ImgReg0IN_41, ImgReg0IN_40, 
      ImgReg0IN_39, ImgReg0IN_38, ImgReg0IN_37, ImgReg0IN_36, ImgReg0IN_35, 
      ImgReg0IN_34, ImgReg0IN_33, ImgReg0IN_32, ImgReg0IN_31, ImgReg0IN_30, 
      ImgReg0IN_29, ImgReg0IN_28, ImgReg0IN_27, ImgReg0IN_26, ImgReg0IN_25, 
      ImgReg0IN_24, ImgReg0IN_23, ImgReg0IN_22, ImgReg0IN_21, ImgReg0IN_20, 
      ImgReg0IN_19, ImgReg0IN_18, ImgReg0IN_17, ImgReg0IN_16, ImgReg0IN_15, 
      ImgReg0IN_14, ImgReg0IN_13, ImgReg0IN_12, ImgReg0IN_11, ImgReg0IN_10, 
      ImgReg0IN_9, ImgReg0IN_8, ImgReg0IN_7, ImgReg0IN_6, ImgReg0IN_5, 
      ImgReg0IN_4, ImgReg0IN_3, ImgReg0IN_2, ImgReg0IN_1, ImgReg0IN_0, 
      ImgReg1IN_447, ImgReg1IN_446, ImgReg1IN_445, ImgReg1IN_444, 
      ImgReg1IN_443, ImgReg1IN_442, ImgReg1IN_441, ImgReg1IN_440, 
      ImgReg1IN_439, ImgReg1IN_438, ImgReg1IN_437, ImgReg1IN_436, 
      ImgReg1IN_435, ImgReg1IN_434, ImgReg1IN_433, ImgReg1IN_432, 
      ImgReg1IN_431, ImgReg1IN_430, ImgReg1IN_429, ImgReg1IN_428, 
      ImgReg1IN_427, ImgReg1IN_426, ImgReg1IN_425, ImgReg1IN_424, 
      ImgReg1IN_423, ImgReg1IN_422, ImgReg1IN_421, ImgReg1IN_420, 
      ImgReg1IN_419, ImgReg1IN_418, ImgReg1IN_417, ImgReg1IN_416, 
      ImgReg1IN_415, ImgReg1IN_414, ImgReg1IN_413, ImgReg1IN_412, 
      ImgReg1IN_411, ImgReg1IN_410, ImgReg1IN_409, ImgReg1IN_408, 
      ImgReg1IN_407, ImgReg1IN_406, ImgReg1IN_405, ImgReg1IN_404, 
      ImgReg1IN_403, ImgReg1IN_402, ImgReg1IN_401, ImgReg1IN_400, 
      ImgReg1IN_399, ImgReg1IN_398, ImgReg1IN_397, ImgReg1IN_396, 
      ImgReg1IN_395, ImgReg1IN_394, ImgReg1IN_393, ImgReg1IN_392, 
      ImgReg1IN_391, ImgReg1IN_390, ImgReg1IN_389, ImgReg1IN_388, 
      ImgReg1IN_387, ImgReg1IN_386, ImgReg1IN_385, ImgReg1IN_384, 
      ImgReg1IN_383, ImgReg1IN_382, ImgReg1IN_381, ImgReg1IN_380, 
      ImgReg1IN_379, ImgReg1IN_378, ImgReg1IN_377, ImgReg1IN_376, 
      ImgReg1IN_375, ImgReg1IN_374, ImgReg1IN_373, ImgReg1IN_372, 
      ImgReg1IN_371, ImgReg1IN_370, ImgReg1IN_369, ImgReg1IN_368, 
      ImgReg1IN_367, ImgReg1IN_366, ImgReg1IN_365, ImgReg1IN_364, 
      ImgReg1IN_363, ImgReg1IN_362, ImgReg1IN_361, ImgReg1IN_360, 
      ImgReg1IN_359, ImgReg1IN_358, ImgReg1IN_357, ImgReg1IN_356, 
      ImgReg1IN_355, ImgReg1IN_354, ImgReg1IN_353, ImgReg1IN_352, 
      ImgReg1IN_351, ImgReg1IN_350, ImgReg1IN_349, ImgReg1IN_348, 
      ImgReg1IN_347, ImgReg1IN_346, ImgReg1IN_345, ImgReg1IN_344, 
      ImgReg1IN_343, ImgReg1IN_342, ImgReg1IN_341, ImgReg1IN_340, 
      ImgReg1IN_339, ImgReg1IN_338, ImgReg1IN_337, ImgReg1IN_336, 
      ImgReg1IN_335, ImgReg1IN_334, ImgReg1IN_333, ImgReg1IN_332, 
      ImgReg1IN_331, ImgReg1IN_330, ImgReg1IN_329, ImgReg1IN_328, 
      ImgReg1IN_327, ImgReg1IN_326, ImgReg1IN_325, ImgReg1IN_324, 
      ImgReg1IN_323, ImgReg1IN_322, ImgReg1IN_321, ImgReg1IN_320, 
      ImgReg1IN_319, ImgReg1IN_318, ImgReg1IN_317, ImgReg1IN_316, 
      ImgReg1IN_315, ImgReg1IN_314, ImgReg1IN_313, ImgReg1IN_312, 
      ImgReg1IN_311, ImgReg1IN_310, ImgReg1IN_309, ImgReg1IN_308, 
      ImgReg1IN_307, ImgReg1IN_306, ImgReg1IN_305, ImgReg1IN_304, 
      ImgReg1IN_303, ImgReg1IN_302, ImgReg1IN_301, ImgReg1IN_300, 
      ImgReg1IN_299, ImgReg1IN_298, ImgReg1IN_297, ImgReg1IN_296, 
      ImgReg1IN_295, ImgReg1IN_294, ImgReg1IN_293, ImgReg1IN_292, 
      ImgReg1IN_291, ImgReg1IN_290, ImgReg1IN_289, ImgReg1IN_288, 
      ImgReg1IN_287, ImgReg1IN_286, ImgReg1IN_285, ImgReg1IN_284, 
      ImgReg1IN_283, ImgReg1IN_282, ImgReg1IN_281, ImgReg1IN_280, 
      ImgReg1IN_279, ImgReg1IN_278, ImgReg1IN_277, ImgReg1IN_276, 
      ImgReg1IN_275, ImgReg1IN_274, ImgReg1IN_273, ImgReg1IN_272, 
      ImgReg1IN_271, ImgReg1IN_270, ImgReg1IN_269, ImgReg1IN_268, 
      ImgReg1IN_267, ImgReg1IN_266, ImgReg1IN_265, ImgReg1IN_264, 
      ImgReg1IN_263, ImgReg1IN_262, ImgReg1IN_261, ImgReg1IN_260, 
      ImgReg1IN_259, ImgReg1IN_258, ImgReg1IN_257, ImgReg1IN_256, 
      ImgReg1IN_255, ImgReg1IN_254, ImgReg1IN_253, ImgReg1IN_252, 
      ImgReg1IN_251, ImgReg1IN_250, ImgReg1IN_249, ImgReg1IN_248, 
      ImgReg1IN_247, ImgReg1IN_246, ImgReg1IN_245, ImgReg1IN_244, 
      ImgReg1IN_243, ImgReg1IN_242, ImgReg1IN_241, ImgReg1IN_240, 
      ImgReg1IN_239, ImgReg1IN_238, ImgReg1IN_237, ImgReg1IN_236, 
      ImgReg1IN_235, ImgReg1IN_234, ImgReg1IN_233, ImgReg1IN_232, 
      ImgReg1IN_231, ImgReg1IN_230, ImgReg1IN_229, ImgReg1IN_228, 
      ImgReg1IN_227, ImgReg1IN_226, ImgReg1IN_225, ImgReg1IN_224, 
      ImgReg1IN_223, ImgReg1IN_222, ImgReg1IN_221, ImgReg1IN_220, 
      ImgReg1IN_219, ImgReg1IN_218, ImgReg1IN_217, ImgReg1IN_216, 
      ImgReg1IN_215, ImgReg1IN_214, ImgReg1IN_213, ImgReg1IN_212, 
      ImgReg1IN_211, ImgReg1IN_210, ImgReg1IN_209, ImgReg1IN_208, 
      ImgReg1IN_207, ImgReg1IN_206, ImgReg1IN_205, ImgReg1IN_204, 
      ImgReg1IN_203, ImgReg1IN_202, ImgReg1IN_201, ImgReg1IN_200, 
      ImgReg1IN_199, ImgReg1IN_198, ImgReg1IN_197, ImgReg1IN_196, 
      ImgReg1IN_195, ImgReg1IN_194, ImgReg1IN_193, ImgReg1IN_192, 
      ImgReg1IN_191, ImgReg1IN_190, ImgReg1IN_189, ImgReg1IN_188, 
      ImgReg1IN_187, ImgReg1IN_186, ImgReg1IN_185, ImgReg1IN_184, 
      ImgReg1IN_183, ImgReg1IN_182, ImgReg1IN_181, ImgReg1IN_180, 
      ImgReg1IN_179, ImgReg1IN_178, ImgReg1IN_177, ImgReg1IN_176, 
      ImgReg1IN_175, ImgReg1IN_174, ImgReg1IN_173, ImgReg1IN_172, 
      ImgReg1IN_171, ImgReg1IN_170, ImgReg1IN_169, ImgReg1IN_168, 
      ImgReg1IN_167, ImgReg1IN_166, ImgReg1IN_165, ImgReg1IN_164, 
      ImgReg1IN_163, ImgReg1IN_162, ImgReg1IN_161, ImgReg1IN_160, 
      ImgReg1IN_159, ImgReg1IN_158, ImgReg1IN_157, ImgReg1IN_156, 
      ImgReg1IN_155, ImgReg1IN_154, ImgReg1IN_153, ImgReg1IN_152, 
      ImgReg1IN_151, ImgReg1IN_150, ImgReg1IN_149, ImgReg1IN_148, 
      ImgReg1IN_147, ImgReg1IN_146, ImgReg1IN_145, ImgReg1IN_144, 
      ImgReg1IN_143, ImgReg1IN_142, ImgReg1IN_141, ImgReg1IN_140, 
      ImgReg1IN_139, ImgReg1IN_138, ImgReg1IN_137, ImgReg1IN_136, 
      ImgReg1IN_135, ImgReg1IN_134, ImgReg1IN_133, ImgReg1IN_132, 
      ImgReg1IN_131, ImgReg1IN_130, ImgReg1IN_129, ImgReg1IN_128, 
      ImgReg1IN_127, ImgReg1IN_126, ImgReg1IN_125, ImgReg1IN_124, 
      ImgReg1IN_123, ImgReg1IN_122, ImgReg1IN_121, ImgReg1IN_120, 
      ImgReg1IN_119, ImgReg1IN_118, ImgReg1IN_117, ImgReg1IN_116, 
      ImgReg1IN_115, ImgReg1IN_114, ImgReg1IN_113, ImgReg1IN_112, 
      ImgReg1IN_111, ImgReg1IN_110, ImgReg1IN_109, ImgReg1IN_108, 
      ImgReg1IN_107, ImgReg1IN_106, ImgReg1IN_105, ImgReg1IN_104, 
      ImgReg1IN_103, ImgReg1IN_102, ImgReg1IN_101, ImgReg1IN_100, 
      ImgReg1IN_99, ImgReg1IN_98, ImgReg1IN_97, ImgReg1IN_96, ImgReg1IN_95, 
      ImgReg1IN_94, ImgReg1IN_93, ImgReg1IN_92, ImgReg1IN_91, ImgReg1IN_90, 
      ImgReg1IN_89, ImgReg1IN_88, ImgReg1IN_87, ImgReg1IN_86, ImgReg1IN_85, 
      ImgReg1IN_84, ImgReg1IN_83, ImgReg1IN_82, ImgReg1IN_81, ImgReg1IN_80, 
      ImgReg1IN_79, ImgReg1IN_78, ImgReg1IN_77, ImgReg1IN_76, ImgReg1IN_75, 
      ImgReg1IN_74, ImgReg1IN_73, ImgReg1IN_72, ImgReg1IN_71, ImgReg1IN_70, 
      ImgReg1IN_69, ImgReg1IN_68, ImgReg1IN_67, ImgReg1IN_66, ImgReg1IN_65, 
      ImgReg1IN_64, ImgReg1IN_63, ImgReg1IN_62, ImgReg1IN_61, ImgReg1IN_60, 
      ImgReg1IN_59, ImgReg1IN_58, ImgReg1IN_57, ImgReg1IN_56, ImgReg1IN_55, 
      ImgReg1IN_54, ImgReg1IN_53, ImgReg1IN_52, ImgReg1IN_51, ImgReg1IN_50, 
      ImgReg1IN_49, ImgReg1IN_48, ImgReg1IN_47, ImgReg1IN_46, ImgReg1IN_45, 
      ImgReg1IN_44, ImgReg1IN_43, ImgReg1IN_42, ImgReg1IN_41, ImgReg1IN_40, 
      ImgReg1IN_39, ImgReg1IN_38, ImgReg1IN_37, ImgReg1IN_36, ImgReg1IN_35, 
      ImgReg1IN_34, ImgReg1IN_33, ImgReg1IN_32, ImgReg1IN_31, ImgReg1IN_30, 
      ImgReg1IN_29, ImgReg1IN_28, ImgReg1IN_27, ImgReg1IN_26, ImgReg1IN_25, 
      ImgReg1IN_24, ImgReg1IN_23, ImgReg1IN_22, ImgReg1IN_21, ImgReg1IN_20, 
      ImgReg1IN_19, ImgReg1IN_18, ImgReg1IN_17, ImgReg1IN_16, ImgReg1IN_15, 
      ImgReg1IN_14, ImgReg1IN_13, ImgReg1IN_12, ImgReg1IN_11, ImgReg1IN_10, 
      ImgReg1IN_9, ImgReg1IN_8, ImgReg1IN_7, ImgReg1IN_6, ImgReg1IN_5, 
      ImgReg1IN_4, ImgReg1IN_3, ImgReg1IN_2, ImgReg1IN_1, ImgReg1IN_0, 
      ImgReg2IN_447, ImgReg2IN_446, ImgReg2IN_445, ImgReg2IN_444, 
      ImgReg2IN_443, ImgReg2IN_442, ImgReg2IN_441, ImgReg2IN_440, 
      ImgReg2IN_439, ImgReg2IN_438, ImgReg2IN_437, ImgReg2IN_436, 
      ImgReg2IN_435, ImgReg2IN_434, ImgReg2IN_433, ImgReg2IN_432, 
      ImgReg2IN_431, ImgReg2IN_430, ImgReg2IN_429, ImgReg2IN_428, 
      ImgReg2IN_427, ImgReg2IN_426, ImgReg2IN_425, ImgReg2IN_424, 
      ImgReg2IN_423, ImgReg2IN_422, ImgReg2IN_421, ImgReg2IN_420, 
      ImgReg2IN_419, ImgReg2IN_418, ImgReg2IN_417, ImgReg2IN_416, 
      ImgReg2IN_415, ImgReg2IN_414, ImgReg2IN_413, ImgReg2IN_412, 
      ImgReg2IN_411, ImgReg2IN_410, ImgReg2IN_409, ImgReg2IN_408, 
      ImgReg2IN_407, ImgReg2IN_406, ImgReg2IN_405, ImgReg2IN_404, 
      ImgReg2IN_403, ImgReg2IN_402, ImgReg2IN_401, ImgReg2IN_400, 
      ImgReg2IN_399, ImgReg2IN_398, ImgReg2IN_397, ImgReg2IN_396, 
      ImgReg2IN_395, ImgReg2IN_394, ImgReg2IN_393, ImgReg2IN_392, 
      ImgReg2IN_391, ImgReg2IN_390, ImgReg2IN_389, ImgReg2IN_388, 
      ImgReg2IN_387, ImgReg2IN_386, ImgReg2IN_385, ImgReg2IN_384, 
      ImgReg2IN_383, ImgReg2IN_382, ImgReg2IN_381, ImgReg2IN_380, 
      ImgReg2IN_379, ImgReg2IN_378, ImgReg2IN_377, ImgReg2IN_376, 
      ImgReg2IN_375, ImgReg2IN_374, ImgReg2IN_373, ImgReg2IN_372, 
      ImgReg2IN_371, ImgReg2IN_370, ImgReg2IN_369, ImgReg2IN_368, 
      ImgReg2IN_367, ImgReg2IN_366, ImgReg2IN_365, ImgReg2IN_364, 
      ImgReg2IN_363, ImgReg2IN_362, ImgReg2IN_361, ImgReg2IN_360, 
      ImgReg2IN_359, ImgReg2IN_358, ImgReg2IN_357, ImgReg2IN_356, 
      ImgReg2IN_355, ImgReg2IN_354, ImgReg2IN_353, ImgReg2IN_352, 
      ImgReg2IN_351, ImgReg2IN_350, ImgReg2IN_349, ImgReg2IN_348, 
      ImgReg2IN_347, ImgReg2IN_346, ImgReg2IN_345, ImgReg2IN_344, 
      ImgReg2IN_343, ImgReg2IN_342, ImgReg2IN_341, ImgReg2IN_340, 
      ImgReg2IN_339, ImgReg2IN_338, ImgReg2IN_337, ImgReg2IN_336, 
      ImgReg2IN_335, ImgReg2IN_334, ImgReg2IN_333, ImgReg2IN_332, 
      ImgReg2IN_331, ImgReg2IN_330, ImgReg2IN_329, ImgReg2IN_328, 
      ImgReg2IN_327, ImgReg2IN_326, ImgReg2IN_325, ImgReg2IN_324, 
      ImgReg2IN_323, ImgReg2IN_322, ImgReg2IN_321, ImgReg2IN_320, 
      ImgReg2IN_319, ImgReg2IN_318, ImgReg2IN_317, ImgReg2IN_316, 
      ImgReg2IN_315, ImgReg2IN_314, ImgReg2IN_313, ImgReg2IN_312, 
      ImgReg2IN_311, ImgReg2IN_310, ImgReg2IN_309, ImgReg2IN_308, 
      ImgReg2IN_307, ImgReg2IN_306, ImgReg2IN_305, ImgReg2IN_304, 
      ImgReg2IN_303, ImgReg2IN_302, ImgReg2IN_301, ImgReg2IN_300, 
      ImgReg2IN_299, ImgReg2IN_298, ImgReg2IN_297, ImgReg2IN_296, 
      ImgReg2IN_295, ImgReg2IN_294, ImgReg2IN_293, ImgReg2IN_292, 
      ImgReg2IN_291, ImgReg2IN_290, ImgReg2IN_289, ImgReg2IN_288, 
      ImgReg2IN_287, ImgReg2IN_286, ImgReg2IN_285, ImgReg2IN_284, 
      ImgReg2IN_283, ImgReg2IN_282, ImgReg2IN_281, ImgReg2IN_280, 
      ImgReg2IN_279, ImgReg2IN_278, ImgReg2IN_277, ImgReg2IN_276, 
      ImgReg2IN_275, ImgReg2IN_274, ImgReg2IN_273, ImgReg2IN_272, 
      ImgReg2IN_271, ImgReg2IN_270, ImgReg2IN_269, ImgReg2IN_268, 
      ImgReg2IN_267, ImgReg2IN_266, ImgReg2IN_265, ImgReg2IN_264, 
      ImgReg2IN_263, ImgReg2IN_262, ImgReg2IN_261, ImgReg2IN_260, 
      ImgReg2IN_259, ImgReg2IN_258, ImgReg2IN_257, ImgReg2IN_256, 
      ImgReg2IN_255, ImgReg2IN_254, ImgReg2IN_253, ImgReg2IN_252, 
      ImgReg2IN_251, ImgReg2IN_250, ImgReg2IN_249, ImgReg2IN_248, 
      ImgReg2IN_247, ImgReg2IN_246, ImgReg2IN_245, ImgReg2IN_244, 
      ImgReg2IN_243, ImgReg2IN_242, ImgReg2IN_241, ImgReg2IN_240, 
      ImgReg2IN_239, ImgReg2IN_238, ImgReg2IN_237, ImgReg2IN_236, 
      ImgReg2IN_235, ImgReg2IN_234, ImgReg2IN_233, ImgReg2IN_232, 
      ImgReg2IN_231, ImgReg2IN_230, ImgReg2IN_229, ImgReg2IN_228, 
      ImgReg2IN_227, ImgReg2IN_226, ImgReg2IN_225, ImgReg2IN_224, 
      ImgReg2IN_223, ImgReg2IN_222, ImgReg2IN_221, ImgReg2IN_220, 
      ImgReg2IN_219, ImgReg2IN_218, ImgReg2IN_217, ImgReg2IN_216, 
      ImgReg2IN_215, ImgReg2IN_214, ImgReg2IN_213, ImgReg2IN_212, 
      ImgReg2IN_211, ImgReg2IN_210, ImgReg2IN_209, ImgReg2IN_208, 
      ImgReg2IN_207, ImgReg2IN_206, ImgReg2IN_205, ImgReg2IN_204, 
      ImgReg2IN_203, ImgReg2IN_202, ImgReg2IN_201, ImgReg2IN_200, 
      ImgReg2IN_199, ImgReg2IN_198, ImgReg2IN_197, ImgReg2IN_196, 
      ImgReg2IN_195, ImgReg2IN_194, ImgReg2IN_193, ImgReg2IN_192, 
      ImgReg2IN_191, ImgReg2IN_190, ImgReg2IN_189, ImgReg2IN_188, 
      ImgReg2IN_187, ImgReg2IN_186, ImgReg2IN_185, ImgReg2IN_184, 
      ImgReg2IN_183, ImgReg2IN_182, ImgReg2IN_181, ImgReg2IN_180, 
      ImgReg2IN_179, ImgReg2IN_178, ImgReg2IN_177, ImgReg2IN_176, 
      ImgReg2IN_175, ImgReg2IN_174, ImgReg2IN_173, ImgReg2IN_172, 
      ImgReg2IN_171, ImgReg2IN_170, ImgReg2IN_169, ImgReg2IN_168, 
      ImgReg2IN_167, ImgReg2IN_166, ImgReg2IN_165, ImgReg2IN_164, 
      ImgReg2IN_163, ImgReg2IN_162, ImgReg2IN_161, ImgReg2IN_160, 
      ImgReg2IN_159, ImgReg2IN_158, ImgReg2IN_157, ImgReg2IN_156, 
      ImgReg2IN_155, ImgReg2IN_154, ImgReg2IN_153, ImgReg2IN_152, 
      ImgReg2IN_151, ImgReg2IN_150, ImgReg2IN_149, ImgReg2IN_148, 
      ImgReg2IN_147, ImgReg2IN_146, ImgReg2IN_145, ImgReg2IN_144, 
      ImgReg2IN_143, ImgReg2IN_142, ImgReg2IN_141, ImgReg2IN_140, 
      ImgReg2IN_139, ImgReg2IN_138, ImgReg2IN_137, ImgReg2IN_136, 
      ImgReg2IN_135, ImgReg2IN_134, ImgReg2IN_133, ImgReg2IN_132, 
      ImgReg2IN_131, ImgReg2IN_130, ImgReg2IN_129, ImgReg2IN_128, 
      ImgReg2IN_127, ImgReg2IN_126, ImgReg2IN_125, ImgReg2IN_124, 
      ImgReg2IN_123, ImgReg2IN_122, ImgReg2IN_121, ImgReg2IN_120, 
      ImgReg2IN_119, ImgReg2IN_118, ImgReg2IN_117, ImgReg2IN_116, 
      ImgReg2IN_115, ImgReg2IN_114, ImgReg2IN_113, ImgReg2IN_112, 
      ImgReg2IN_111, ImgReg2IN_110, ImgReg2IN_109, ImgReg2IN_108, 
      ImgReg2IN_107, ImgReg2IN_106, ImgReg2IN_105, ImgReg2IN_104, 
      ImgReg2IN_103, ImgReg2IN_102, ImgReg2IN_101, ImgReg2IN_100, 
      ImgReg2IN_99, ImgReg2IN_98, ImgReg2IN_97, ImgReg2IN_96, ImgReg2IN_95, 
      ImgReg2IN_94, ImgReg2IN_93, ImgReg2IN_92, ImgReg2IN_91, ImgReg2IN_90, 
      ImgReg2IN_89, ImgReg2IN_88, ImgReg2IN_87, ImgReg2IN_86, ImgReg2IN_85, 
      ImgReg2IN_84, ImgReg2IN_83, ImgReg2IN_82, ImgReg2IN_81, ImgReg2IN_80, 
      ImgReg2IN_79, ImgReg2IN_78, ImgReg2IN_77, ImgReg2IN_76, ImgReg2IN_75, 
      ImgReg2IN_74, ImgReg2IN_73, ImgReg2IN_72, ImgReg2IN_71, ImgReg2IN_70, 
      ImgReg2IN_69, ImgReg2IN_68, ImgReg2IN_67, ImgReg2IN_66, ImgReg2IN_65, 
      ImgReg2IN_64, ImgReg2IN_63, ImgReg2IN_62, ImgReg2IN_61, ImgReg2IN_60, 
      ImgReg2IN_59, ImgReg2IN_58, ImgReg2IN_57, ImgReg2IN_56, ImgReg2IN_55, 
      ImgReg2IN_54, ImgReg2IN_53, ImgReg2IN_52, ImgReg2IN_51, ImgReg2IN_50, 
      ImgReg2IN_49, ImgReg2IN_48, ImgReg2IN_47, ImgReg2IN_46, ImgReg2IN_45, 
      ImgReg2IN_44, ImgReg2IN_43, ImgReg2IN_42, ImgReg2IN_41, ImgReg2IN_40, 
      ImgReg2IN_39, ImgReg2IN_38, ImgReg2IN_37, ImgReg2IN_36, ImgReg2IN_35, 
      ImgReg2IN_34, ImgReg2IN_33, ImgReg2IN_32, ImgReg2IN_31, ImgReg2IN_30, 
      ImgReg2IN_29, ImgReg2IN_28, ImgReg2IN_27, ImgReg2IN_26, ImgReg2IN_25, 
      ImgReg2IN_24, ImgReg2IN_23, ImgReg2IN_22, ImgReg2IN_21, ImgReg2IN_20, 
      ImgReg2IN_19, ImgReg2IN_18, ImgReg2IN_17, ImgReg2IN_16, ImgReg2IN_15, 
      ImgReg2IN_14, ImgReg2IN_13, ImgReg2IN_12, ImgReg2IN_11, ImgReg2IN_10, 
      ImgReg2IN_9, ImgReg2IN_8, ImgReg2IN_7, ImgReg2IN_6, ImgReg2IN_5, 
      ImgReg2IN_4, ImgReg2IN_3, ImgReg2IN_2, ImgReg2IN_1, ImgReg2IN_0, 
      ImgReg3IN_447, ImgReg3IN_446, ImgReg3IN_445, ImgReg3IN_444, 
      ImgReg3IN_443, ImgReg3IN_442, ImgReg3IN_441, ImgReg3IN_440, 
      ImgReg3IN_439, ImgReg3IN_438, ImgReg3IN_437, ImgReg3IN_436, 
      ImgReg3IN_435, ImgReg3IN_434, ImgReg3IN_433, ImgReg3IN_432, 
      ImgReg3IN_431, ImgReg3IN_430, ImgReg3IN_429, ImgReg3IN_428, 
      ImgReg3IN_427, ImgReg3IN_426, ImgReg3IN_425, ImgReg3IN_424, 
      ImgReg3IN_423, ImgReg3IN_422, ImgReg3IN_421, ImgReg3IN_420, 
      ImgReg3IN_419, ImgReg3IN_418, ImgReg3IN_417, ImgReg3IN_416, 
      ImgReg3IN_415, ImgReg3IN_414, ImgReg3IN_413, ImgReg3IN_412, 
      ImgReg3IN_411, ImgReg3IN_410, ImgReg3IN_409, ImgReg3IN_408, 
      ImgReg3IN_407, ImgReg3IN_406, ImgReg3IN_405, ImgReg3IN_404, 
      ImgReg3IN_403, ImgReg3IN_402, ImgReg3IN_401, ImgReg3IN_400, 
      ImgReg3IN_399, ImgReg3IN_398, ImgReg3IN_397, ImgReg3IN_396, 
      ImgReg3IN_395, ImgReg3IN_394, ImgReg3IN_393, ImgReg3IN_392, 
      ImgReg3IN_391, ImgReg3IN_390, ImgReg3IN_389, ImgReg3IN_388, 
      ImgReg3IN_387, ImgReg3IN_386, ImgReg3IN_385, ImgReg3IN_384, 
      ImgReg3IN_383, ImgReg3IN_382, ImgReg3IN_381, ImgReg3IN_380, 
      ImgReg3IN_379, ImgReg3IN_378, ImgReg3IN_377, ImgReg3IN_376, 
      ImgReg3IN_375, ImgReg3IN_374, ImgReg3IN_373, ImgReg3IN_372, 
      ImgReg3IN_371, ImgReg3IN_370, ImgReg3IN_369, ImgReg3IN_368, 
      ImgReg3IN_367, ImgReg3IN_366, ImgReg3IN_365, ImgReg3IN_364, 
      ImgReg3IN_363, ImgReg3IN_362, ImgReg3IN_361, ImgReg3IN_360, 
      ImgReg3IN_359, ImgReg3IN_358, ImgReg3IN_357, ImgReg3IN_356, 
      ImgReg3IN_355, ImgReg3IN_354, ImgReg3IN_353, ImgReg3IN_352, 
      ImgReg3IN_351, ImgReg3IN_350, ImgReg3IN_349, ImgReg3IN_348, 
      ImgReg3IN_347, ImgReg3IN_346, ImgReg3IN_345, ImgReg3IN_344, 
      ImgReg3IN_343, ImgReg3IN_342, ImgReg3IN_341, ImgReg3IN_340, 
      ImgReg3IN_339, ImgReg3IN_338, ImgReg3IN_337, ImgReg3IN_336, 
      ImgReg3IN_335, ImgReg3IN_334, ImgReg3IN_333, ImgReg3IN_332, 
      ImgReg3IN_331, ImgReg3IN_330, ImgReg3IN_329, ImgReg3IN_328, 
      ImgReg3IN_327, ImgReg3IN_326, ImgReg3IN_325, ImgReg3IN_324, 
      ImgReg3IN_323, ImgReg3IN_322, ImgReg3IN_321, ImgReg3IN_320, 
      ImgReg3IN_319, ImgReg3IN_318, ImgReg3IN_317, ImgReg3IN_316, 
      ImgReg3IN_315, ImgReg3IN_314, ImgReg3IN_313, ImgReg3IN_312, 
      ImgReg3IN_311, ImgReg3IN_310, ImgReg3IN_309, ImgReg3IN_308, 
      ImgReg3IN_307, ImgReg3IN_306, ImgReg3IN_305, ImgReg3IN_304, 
      ImgReg3IN_303, ImgReg3IN_302, ImgReg3IN_301, ImgReg3IN_300, 
      ImgReg3IN_299, ImgReg3IN_298, ImgReg3IN_297, ImgReg3IN_296, 
      ImgReg3IN_295, ImgReg3IN_294, ImgReg3IN_293, ImgReg3IN_292, 
      ImgReg3IN_291, ImgReg3IN_290, ImgReg3IN_289, ImgReg3IN_288, 
      ImgReg3IN_287, ImgReg3IN_286, ImgReg3IN_285, ImgReg3IN_284, 
      ImgReg3IN_283, ImgReg3IN_282, ImgReg3IN_281, ImgReg3IN_280, 
      ImgReg3IN_279, ImgReg3IN_278, ImgReg3IN_277, ImgReg3IN_276, 
      ImgReg3IN_275, ImgReg3IN_274, ImgReg3IN_273, ImgReg3IN_272, 
      ImgReg3IN_271, ImgReg3IN_270, ImgReg3IN_269, ImgReg3IN_268, 
      ImgReg3IN_267, ImgReg3IN_266, ImgReg3IN_265, ImgReg3IN_264, 
      ImgReg3IN_263, ImgReg3IN_262, ImgReg3IN_261, ImgReg3IN_260, 
      ImgReg3IN_259, ImgReg3IN_258, ImgReg3IN_257, ImgReg3IN_256, 
      ImgReg3IN_255, ImgReg3IN_254, ImgReg3IN_253, ImgReg3IN_252, 
      ImgReg3IN_251, ImgReg3IN_250, ImgReg3IN_249, ImgReg3IN_248, 
      ImgReg3IN_247, ImgReg3IN_246, ImgReg3IN_245, ImgReg3IN_244, 
      ImgReg3IN_243, ImgReg3IN_242, ImgReg3IN_241, ImgReg3IN_240, 
      ImgReg3IN_239, ImgReg3IN_238, ImgReg3IN_237, ImgReg3IN_236, 
      ImgReg3IN_235, ImgReg3IN_234, ImgReg3IN_233, ImgReg3IN_232, 
      ImgReg3IN_231, ImgReg3IN_230, ImgReg3IN_229, ImgReg3IN_228, 
      ImgReg3IN_227, ImgReg3IN_226, ImgReg3IN_225, ImgReg3IN_224, 
      ImgReg3IN_223, ImgReg3IN_222, ImgReg3IN_221, ImgReg3IN_220, 
      ImgReg3IN_219, ImgReg3IN_218, ImgReg3IN_217, ImgReg3IN_216, 
      ImgReg3IN_215, ImgReg3IN_214, ImgReg3IN_213, ImgReg3IN_212, 
      ImgReg3IN_211, ImgReg3IN_210, ImgReg3IN_209, ImgReg3IN_208, 
      ImgReg3IN_207, ImgReg3IN_206, ImgReg3IN_205, ImgReg3IN_204, 
      ImgReg3IN_203, ImgReg3IN_202, ImgReg3IN_201, ImgReg3IN_200, 
      ImgReg3IN_199, ImgReg3IN_198, ImgReg3IN_197, ImgReg3IN_196, 
      ImgReg3IN_195, ImgReg3IN_194, ImgReg3IN_193, ImgReg3IN_192, 
      ImgReg3IN_191, ImgReg3IN_190, ImgReg3IN_189, ImgReg3IN_188, 
      ImgReg3IN_187, ImgReg3IN_186, ImgReg3IN_185, ImgReg3IN_184, 
      ImgReg3IN_183, ImgReg3IN_182, ImgReg3IN_181, ImgReg3IN_180, 
      ImgReg3IN_179, ImgReg3IN_178, ImgReg3IN_177, ImgReg3IN_176, 
      ImgReg3IN_175, ImgReg3IN_174, ImgReg3IN_173, ImgReg3IN_172, 
      ImgReg3IN_171, ImgReg3IN_170, ImgReg3IN_169, ImgReg3IN_168, 
      ImgReg3IN_167, ImgReg3IN_166, ImgReg3IN_165, ImgReg3IN_164, 
      ImgReg3IN_163, ImgReg3IN_162, ImgReg3IN_161, ImgReg3IN_160, 
      ImgReg3IN_159, ImgReg3IN_158, ImgReg3IN_157, ImgReg3IN_156, 
      ImgReg3IN_155, ImgReg3IN_154, ImgReg3IN_153, ImgReg3IN_152, 
      ImgReg3IN_151, ImgReg3IN_150, ImgReg3IN_149, ImgReg3IN_148, 
      ImgReg3IN_147, ImgReg3IN_146, ImgReg3IN_145, ImgReg3IN_144, 
      ImgReg3IN_143, ImgReg3IN_142, ImgReg3IN_141, ImgReg3IN_140, 
      ImgReg3IN_139, ImgReg3IN_138, ImgReg3IN_137, ImgReg3IN_136, 
      ImgReg3IN_135, ImgReg3IN_134, ImgReg3IN_133, ImgReg3IN_132, 
      ImgReg3IN_131, ImgReg3IN_130, ImgReg3IN_129, ImgReg3IN_128, 
      ImgReg3IN_127, ImgReg3IN_126, ImgReg3IN_125, ImgReg3IN_124, 
      ImgReg3IN_123, ImgReg3IN_122, ImgReg3IN_121, ImgReg3IN_120, 
      ImgReg3IN_119, ImgReg3IN_118, ImgReg3IN_117, ImgReg3IN_116, 
      ImgReg3IN_115, ImgReg3IN_114, ImgReg3IN_113, ImgReg3IN_112, 
      ImgReg3IN_111, ImgReg3IN_110, ImgReg3IN_109, ImgReg3IN_108, 
      ImgReg3IN_107, ImgReg3IN_106, ImgReg3IN_105, ImgReg3IN_104, 
      ImgReg3IN_103, ImgReg3IN_102, ImgReg3IN_101, ImgReg3IN_100, 
      ImgReg3IN_99, ImgReg3IN_98, ImgReg3IN_97, ImgReg3IN_96, ImgReg3IN_95, 
      ImgReg3IN_94, ImgReg3IN_93, ImgReg3IN_92, ImgReg3IN_91, ImgReg3IN_90, 
      ImgReg3IN_89, ImgReg3IN_88, ImgReg3IN_87, ImgReg3IN_86, ImgReg3IN_85, 
      ImgReg3IN_84, ImgReg3IN_83, ImgReg3IN_82, ImgReg3IN_81, ImgReg3IN_80, 
      ImgReg3IN_79, ImgReg3IN_78, ImgReg3IN_77, ImgReg3IN_76, ImgReg3IN_75, 
      ImgReg3IN_74, ImgReg3IN_73, ImgReg3IN_72, ImgReg3IN_71, ImgReg3IN_70, 
      ImgReg3IN_69, ImgReg3IN_68, ImgReg3IN_67, ImgReg3IN_66, ImgReg3IN_65, 
      ImgReg3IN_64, ImgReg3IN_63, ImgReg3IN_62, ImgReg3IN_61, ImgReg3IN_60, 
      ImgReg3IN_59, ImgReg3IN_58, ImgReg3IN_57, ImgReg3IN_56, ImgReg3IN_55, 
      ImgReg3IN_54, ImgReg3IN_53, ImgReg3IN_52, ImgReg3IN_51, ImgReg3IN_50, 
      ImgReg3IN_49, ImgReg3IN_48, ImgReg3IN_47, ImgReg3IN_46, ImgReg3IN_45, 
      ImgReg3IN_44, ImgReg3IN_43, ImgReg3IN_42, ImgReg3IN_41, ImgReg3IN_40, 
      ImgReg3IN_39, ImgReg3IN_38, ImgReg3IN_37, ImgReg3IN_36, ImgReg3IN_35, 
      ImgReg3IN_34, ImgReg3IN_33, ImgReg3IN_32, ImgReg3IN_31, ImgReg3IN_30, 
      ImgReg3IN_29, ImgReg3IN_28, ImgReg3IN_27, ImgReg3IN_26, ImgReg3IN_25, 
      ImgReg3IN_24, ImgReg3IN_23, ImgReg3IN_22, ImgReg3IN_21, ImgReg3IN_20, 
      ImgReg3IN_19, ImgReg3IN_18, ImgReg3IN_17, ImgReg3IN_16, ImgReg3IN_15, 
      ImgReg3IN_14, ImgReg3IN_13, ImgReg3IN_12, ImgReg3IN_11, ImgReg3IN_10, 
      ImgReg3IN_9, ImgReg3IN_8, ImgReg3IN_7, ImgReg3IN_6, ImgReg3IN_5, 
      ImgReg3IN_4, ImgReg3IN_3, ImgReg3IN_2, ImgReg3IN_1, ImgReg3IN_0, 
      ImgReg4IN_447, ImgReg4IN_446, ImgReg4IN_445, ImgReg4IN_444, 
      ImgReg4IN_443, ImgReg4IN_442, ImgReg4IN_441, ImgReg4IN_440, 
      ImgReg4IN_439, ImgReg4IN_438, ImgReg4IN_437, ImgReg4IN_436, 
      ImgReg4IN_435, ImgReg4IN_434, ImgReg4IN_433, ImgReg4IN_432, 
      ImgReg4IN_431, ImgReg4IN_430, ImgReg4IN_429, ImgReg4IN_428, 
      ImgReg4IN_427, ImgReg4IN_426, ImgReg4IN_425, ImgReg4IN_424, 
      ImgReg4IN_423, ImgReg4IN_422, ImgReg4IN_421, ImgReg4IN_420, 
      ImgReg4IN_419, ImgReg4IN_418, ImgReg4IN_417, ImgReg4IN_416, 
      ImgReg4IN_415, ImgReg4IN_414, ImgReg4IN_413, ImgReg4IN_412, 
      ImgReg4IN_411, ImgReg4IN_410, ImgReg4IN_409, ImgReg4IN_408, 
      ImgReg4IN_407, ImgReg4IN_406, ImgReg4IN_405, ImgReg4IN_404, 
      ImgReg4IN_403, ImgReg4IN_402, ImgReg4IN_401, ImgReg4IN_400, 
      ImgReg4IN_399, ImgReg4IN_398, ImgReg4IN_397, ImgReg4IN_396, 
      ImgReg4IN_395, ImgReg4IN_394, ImgReg4IN_393, ImgReg4IN_392, 
      ImgReg4IN_391, ImgReg4IN_390, ImgReg4IN_389, ImgReg4IN_388, 
      ImgReg4IN_387, ImgReg4IN_386, ImgReg4IN_385, ImgReg4IN_384, 
      ImgReg4IN_383, ImgReg4IN_382, ImgReg4IN_381, ImgReg4IN_380, 
      ImgReg4IN_379, ImgReg4IN_378, ImgReg4IN_377, ImgReg4IN_376, 
      ImgReg4IN_375, ImgReg4IN_374, ImgReg4IN_373, ImgReg4IN_372, 
      ImgReg4IN_371, ImgReg4IN_370, ImgReg4IN_369, ImgReg4IN_368, 
      ImgReg4IN_367, ImgReg4IN_366, ImgReg4IN_365, ImgReg4IN_364, 
      ImgReg4IN_363, ImgReg4IN_362, ImgReg4IN_361, ImgReg4IN_360, 
      ImgReg4IN_359, ImgReg4IN_358, ImgReg4IN_357, ImgReg4IN_356, 
      ImgReg4IN_355, ImgReg4IN_354, ImgReg4IN_353, ImgReg4IN_352, 
      ImgReg4IN_351, ImgReg4IN_350, ImgReg4IN_349, ImgReg4IN_348, 
      ImgReg4IN_347, ImgReg4IN_346, ImgReg4IN_345, ImgReg4IN_344, 
      ImgReg4IN_343, ImgReg4IN_342, ImgReg4IN_341, ImgReg4IN_340, 
      ImgReg4IN_339, ImgReg4IN_338, ImgReg4IN_337, ImgReg4IN_336, 
      ImgReg4IN_335, ImgReg4IN_334, ImgReg4IN_333, ImgReg4IN_332, 
      ImgReg4IN_331, ImgReg4IN_330, ImgReg4IN_329, ImgReg4IN_328, 
      ImgReg4IN_327, ImgReg4IN_326, ImgReg4IN_325, ImgReg4IN_324, 
      ImgReg4IN_323, ImgReg4IN_322, ImgReg4IN_321, ImgReg4IN_320, 
      ImgReg4IN_319, ImgReg4IN_318, ImgReg4IN_317, ImgReg4IN_316, 
      ImgReg4IN_315, ImgReg4IN_314, ImgReg4IN_313, ImgReg4IN_312, 
      ImgReg4IN_311, ImgReg4IN_310, ImgReg4IN_309, ImgReg4IN_308, 
      ImgReg4IN_307, ImgReg4IN_306, ImgReg4IN_305, ImgReg4IN_304, 
      ImgReg4IN_303, ImgReg4IN_302, ImgReg4IN_301, ImgReg4IN_300, 
      ImgReg4IN_299, ImgReg4IN_298, ImgReg4IN_297, ImgReg4IN_296, 
      ImgReg4IN_295, ImgReg4IN_294, ImgReg4IN_293, ImgReg4IN_292, 
      ImgReg4IN_291, ImgReg4IN_290, ImgReg4IN_289, ImgReg4IN_288, 
      ImgReg4IN_287, ImgReg4IN_286, ImgReg4IN_285, ImgReg4IN_284, 
      ImgReg4IN_283, ImgReg4IN_282, ImgReg4IN_281, ImgReg4IN_280, 
      ImgReg4IN_279, ImgReg4IN_278, ImgReg4IN_277, ImgReg4IN_276, 
      ImgReg4IN_275, ImgReg4IN_274, ImgReg4IN_273, ImgReg4IN_272, 
      ImgReg4IN_271, ImgReg4IN_270, ImgReg4IN_269, ImgReg4IN_268, 
      ImgReg4IN_267, ImgReg4IN_266, ImgReg4IN_265, ImgReg4IN_264, 
      ImgReg4IN_263, ImgReg4IN_262, ImgReg4IN_261, ImgReg4IN_260, 
      ImgReg4IN_259, ImgReg4IN_258, ImgReg4IN_257, ImgReg4IN_256, 
      ImgReg4IN_255, ImgReg4IN_254, ImgReg4IN_253, ImgReg4IN_252, 
      ImgReg4IN_251, ImgReg4IN_250, ImgReg4IN_249, ImgReg4IN_248, 
      ImgReg4IN_247, ImgReg4IN_246, ImgReg4IN_245, ImgReg4IN_244, 
      ImgReg4IN_243, ImgReg4IN_242, ImgReg4IN_241, ImgReg4IN_240, 
      ImgReg4IN_239, ImgReg4IN_238, ImgReg4IN_237, ImgReg4IN_236, 
      ImgReg4IN_235, ImgReg4IN_234, ImgReg4IN_233, ImgReg4IN_232, 
      ImgReg4IN_231, ImgReg4IN_230, ImgReg4IN_229, ImgReg4IN_228, 
      ImgReg4IN_227, ImgReg4IN_226, ImgReg4IN_225, ImgReg4IN_224, 
      ImgReg4IN_223, ImgReg4IN_222, ImgReg4IN_221, ImgReg4IN_220, 
      ImgReg4IN_219, ImgReg4IN_218, ImgReg4IN_217, ImgReg4IN_216, 
      ImgReg4IN_215, ImgReg4IN_214, ImgReg4IN_213, ImgReg4IN_212, 
      ImgReg4IN_211, ImgReg4IN_210, ImgReg4IN_209, ImgReg4IN_208, 
      ImgReg4IN_207, ImgReg4IN_206, ImgReg4IN_205, ImgReg4IN_204, 
      ImgReg4IN_203, ImgReg4IN_202, ImgReg4IN_201, ImgReg4IN_200, 
      ImgReg4IN_199, ImgReg4IN_198, ImgReg4IN_197, ImgReg4IN_196, 
      ImgReg4IN_195, ImgReg4IN_194, ImgReg4IN_193, ImgReg4IN_192, 
      ImgReg4IN_191, ImgReg4IN_190, ImgReg4IN_189, ImgReg4IN_188, 
      ImgReg4IN_187, ImgReg4IN_186, ImgReg4IN_185, ImgReg4IN_184, 
      ImgReg4IN_183, ImgReg4IN_182, ImgReg4IN_181, ImgReg4IN_180, 
      ImgReg4IN_179, ImgReg4IN_178, ImgReg4IN_177, ImgReg4IN_176, 
      ImgReg4IN_175, ImgReg4IN_174, ImgReg4IN_173, ImgReg4IN_172, 
      ImgReg4IN_171, ImgReg4IN_170, ImgReg4IN_169, ImgReg4IN_168, 
      ImgReg4IN_167, ImgReg4IN_166, ImgReg4IN_165, ImgReg4IN_164, 
      ImgReg4IN_163, ImgReg4IN_162, ImgReg4IN_161, ImgReg4IN_160, 
      ImgReg4IN_159, ImgReg4IN_158, ImgReg4IN_157, ImgReg4IN_156, 
      ImgReg4IN_155, ImgReg4IN_154, ImgReg4IN_153, ImgReg4IN_152, 
      ImgReg4IN_151, ImgReg4IN_150, ImgReg4IN_149, ImgReg4IN_148, 
      ImgReg4IN_147, ImgReg4IN_146, ImgReg4IN_145, ImgReg4IN_144, 
      ImgReg4IN_143, ImgReg4IN_142, ImgReg4IN_141, ImgReg4IN_140, 
      ImgReg4IN_139, ImgReg4IN_138, ImgReg4IN_137, ImgReg4IN_136, 
      ImgReg4IN_135, ImgReg4IN_134, ImgReg4IN_133, ImgReg4IN_132, 
      ImgReg4IN_131, ImgReg4IN_130, ImgReg4IN_129, ImgReg4IN_128, 
      ImgReg4IN_127, ImgReg4IN_126, ImgReg4IN_125, ImgReg4IN_124, 
      ImgReg4IN_123, ImgReg4IN_122, ImgReg4IN_121, ImgReg4IN_120, 
      ImgReg4IN_119, ImgReg4IN_118, ImgReg4IN_117, ImgReg4IN_116, 
      ImgReg4IN_115, ImgReg4IN_114, ImgReg4IN_113, ImgReg4IN_112, 
      ImgReg4IN_111, ImgReg4IN_110, ImgReg4IN_109, ImgReg4IN_108, 
      ImgReg4IN_107, ImgReg4IN_106, ImgReg4IN_105, ImgReg4IN_104, 
      ImgReg4IN_103, ImgReg4IN_102, ImgReg4IN_101, ImgReg4IN_100, 
      ImgReg4IN_99, ImgReg4IN_98, ImgReg4IN_97, ImgReg4IN_96, ImgReg4IN_95, 
      ImgReg4IN_94, ImgReg4IN_93, ImgReg4IN_92, ImgReg4IN_91, ImgReg4IN_90, 
      ImgReg4IN_89, ImgReg4IN_88, ImgReg4IN_87, ImgReg4IN_86, ImgReg4IN_85, 
      ImgReg4IN_84, ImgReg4IN_83, ImgReg4IN_82, ImgReg4IN_81, ImgReg4IN_80, 
      ImgReg4IN_79, ImgReg4IN_78, ImgReg4IN_77, ImgReg4IN_76, ImgReg4IN_75, 
      ImgReg4IN_74, ImgReg4IN_73, ImgReg4IN_72, ImgReg4IN_71, ImgReg4IN_70, 
      ImgReg4IN_69, ImgReg4IN_68, ImgReg4IN_67, ImgReg4IN_66, ImgReg4IN_65, 
      ImgReg4IN_64, ImgReg4IN_63, ImgReg4IN_62, ImgReg4IN_61, ImgReg4IN_60, 
      ImgReg4IN_59, ImgReg4IN_58, ImgReg4IN_57, ImgReg4IN_56, ImgReg4IN_55, 
      ImgReg4IN_54, ImgReg4IN_53, ImgReg4IN_52, ImgReg4IN_51, ImgReg4IN_50, 
      ImgReg4IN_49, ImgReg4IN_48, ImgReg4IN_47, ImgReg4IN_46, ImgReg4IN_45, 
      ImgReg4IN_44, ImgReg4IN_43, ImgReg4IN_42, ImgReg4IN_41, ImgReg4IN_40, 
      ImgReg4IN_39, ImgReg4IN_38, ImgReg4IN_37, ImgReg4IN_36, ImgReg4IN_35, 
      ImgReg4IN_34, ImgReg4IN_33, ImgReg4IN_32, ImgReg4IN_31, ImgReg4IN_30, 
      ImgReg4IN_29, ImgReg4IN_28, ImgReg4IN_27, ImgReg4IN_26, ImgReg4IN_25, 
      ImgReg4IN_24, ImgReg4IN_23, ImgReg4IN_22, ImgReg4IN_21, ImgReg4IN_20, 
      ImgReg4IN_19, ImgReg4IN_18, ImgReg4IN_17, ImgReg4IN_16, ImgReg4IN_15, 
      ImgReg4IN_14, ImgReg4IN_13, ImgReg4IN_12, ImgReg4IN_11, ImgReg4IN_10, 
      ImgReg4IN_9, ImgReg4IN_8, ImgReg4IN_7, ImgReg4IN_6, ImgReg4IN_5, 
      ImgReg4IN_4, ImgReg4IN_3, ImgReg4IN_2, ImgReg4IN_1, ImgReg4IN_0, 
      ImgReg5IN_447, ImgReg5IN_446, ImgReg5IN_445, ImgReg5IN_444, 
      ImgReg5IN_443, ImgReg5IN_442, ImgReg5IN_441, ImgReg5IN_440, 
      ImgReg5IN_439, ImgReg5IN_438, ImgReg5IN_437, ImgReg5IN_436, 
      ImgReg5IN_435, ImgReg5IN_434, ImgReg5IN_433, ImgReg5IN_432, 
      ImgReg5IN_431, ImgReg5IN_430, ImgReg5IN_429, ImgReg5IN_428, 
      ImgReg5IN_427, ImgReg5IN_426, ImgReg5IN_425, ImgReg5IN_424, 
      ImgReg5IN_423, ImgReg5IN_422, ImgReg5IN_421, ImgReg5IN_420, 
      ImgReg5IN_419, ImgReg5IN_418, ImgReg5IN_417, ImgReg5IN_416, 
      ImgReg5IN_415, ImgReg5IN_414, ImgReg5IN_413, ImgReg5IN_412, 
      ImgReg5IN_411, ImgReg5IN_410, ImgReg5IN_409, ImgReg5IN_408, 
      ImgReg5IN_407, ImgReg5IN_406, ImgReg5IN_405, ImgReg5IN_404, 
      ImgReg5IN_403, ImgReg5IN_402, ImgReg5IN_401, ImgReg5IN_400, 
      ImgReg5IN_399, ImgReg5IN_398, ImgReg5IN_397, ImgReg5IN_396, 
      ImgReg5IN_395, ImgReg5IN_394, ImgReg5IN_393, ImgReg5IN_392, 
      ImgReg5IN_391, ImgReg5IN_390, ImgReg5IN_389, ImgReg5IN_388, 
      ImgReg5IN_387, ImgReg5IN_386, ImgReg5IN_385, ImgReg5IN_384, 
      ImgReg5IN_383, ImgReg5IN_382, ImgReg5IN_381, ImgReg5IN_380, 
      ImgReg5IN_379, ImgReg5IN_378, ImgReg5IN_377, ImgReg5IN_376, 
      ImgReg5IN_375, ImgReg5IN_374, ImgReg5IN_373, ImgReg5IN_372, 
      ImgReg5IN_371, ImgReg5IN_370, ImgReg5IN_369, ImgReg5IN_368, 
      ImgReg5IN_367, ImgReg5IN_366, ImgReg5IN_365, ImgReg5IN_364, 
      ImgReg5IN_363, ImgReg5IN_362, ImgReg5IN_361, ImgReg5IN_360, 
      ImgReg5IN_359, ImgReg5IN_358, ImgReg5IN_357, ImgReg5IN_356, 
      ImgReg5IN_355, ImgReg5IN_354, ImgReg5IN_353, ImgReg5IN_352, 
      ImgReg5IN_351, ImgReg5IN_350, ImgReg5IN_349, ImgReg5IN_348, 
      ImgReg5IN_347, ImgReg5IN_346, ImgReg5IN_345, ImgReg5IN_344, 
      ImgReg5IN_343, ImgReg5IN_342, ImgReg5IN_341, ImgReg5IN_340, 
      ImgReg5IN_339, ImgReg5IN_338, ImgReg5IN_337, ImgReg5IN_336, 
      ImgReg5IN_335, ImgReg5IN_334, ImgReg5IN_333, ImgReg5IN_332, 
      ImgReg5IN_331, ImgReg5IN_330, ImgReg5IN_329, ImgReg5IN_328, 
      ImgReg5IN_327, ImgReg5IN_326, ImgReg5IN_325, ImgReg5IN_324, 
      ImgReg5IN_323, ImgReg5IN_322, ImgReg5IN_321, ImgReg5IN_320, 
      ImgReg5IN_319, ImgReg5IN_318, ImgReg5IN_317, ImgReg5IN_316, 
      ImgReg5IN_315, ImgReg5IN_314, ImgReg5IN_313, ImgReg5IN_312, 
      ImgReg5IN_311, ImgReg5IN_310, ImgReg5IN_309, ImgReg5IN_308, 
      ImgReg5IN_307, ImgReg5IN_306, ImgReg5IN_305, ImgReg5IN_304, 
      ImgReg5IN_303, ImgReg5IN_302, ImgReg5IN_301, ImgReg5IN_300, 
      ImgReg5IN_299, ImgReg5IN_298, ImgReg5IN_297, ImgReg5IN_296, 
      ImgReg5IN_295, ImgReg5IN_294, ImgReg5IN_293, ImgReg5IN_292, 
      ImgReg5IN_291, ImgReg5IN_290, ImgReg5IN_289, ImgReg5IN_288, 
      ImgReg5IN_287, ImgReg5IN_286, ImgReg5IN_285, ImgReg5IN_284, 
      ImgReg5IN_283, ImgReg5IN_282, ImgReg5IN_281, ImgReg5IN_280, 
      ImgReg5IN_279, ImgReg5IN_278, ImgReg5IN_277, ImgReg5IN_276, 
      ImgReg5IN_275, ImgReg5IN_274, ImgReg5IN_273, ImgReg5IN_272, 
      ImgReg5IN_271, ImgReg5IN_270, ImgReg5IN_269, ImgReg5IN_268, 
      ImgReg5IN_267, ImgReg5IN_266, ImgReg5IN_265, ImgReg5IN_264, 
      ImgReg5IN_263, ImgReg5IN_262, ImgReg5IN_261, ImgReg5IN_260, 
      ImgReg5IN_259, ImgReg5IN_258, ImgReg5IN_257, ImgReg5IN_256, 
      ImgReg5IN_255, ImgReg5IN_254, ImgReg5IN_253, ImgReg5IN_252, 
      ImgReg5IN_251, ImgReg5IN_250, ImgReg5IN_249, ImgReg5IN_248, 
      ImgReg5IN_247, ImgReg5IN_246, ImgReg5IN_245, ImgReg5IN_244, 
      ImgReg5IN_243, ImgReg5IN_242, ImgReg5IN_241, ImgReg5IN_240, 
      ImgReg5IN_239, ImgReg5IN_238, ImgReg5IN_237, ImgReg5IN_236, 
      ImgReg5IN_235, ImgReg5IN_234, ImgReg5IN_233, ImgReg5IN_232, 
      ImgReg5IN_231, ImgReg5IN_230, ImgReg5IN_229, ImgReg5IN_228, 
      ImgReg5IN_227, ImgReg5IN_226, ImgReg5IN_225, ImgReg5IN_224, 
      ImgReg5IN_223, ImgReg5IN_222, ImgReg5IN_221, ImgReg5IN_220, 
      ImgReg5IN_219, ImgReg5IN_218, ImgReg5IN_217, ImgReg5IN_216, 
      ImgReg5IN_215, ImgReg5IN_214, ImgReg5IN_213, ImgReg5IN_212, 
      ImgReg5IN_211, ImgReg5IN_210, ImgReg5IN_209, ImgReg5IN_208, 
      ImgReg5IN_207, ImgReg5IN_206, ImgReg5IN_205, ImgReg5IN_204, 
      ImgReg5IN_203, ImgReg5IN_202, ImgReg5IN_201, ImgReg5IN_200, 
      ImgReg5IN_199, ImgReg5IN_198, ImgReg5IN_197, ImgReg5IN_196, 
      ImgReg5IN_195, ImgReg5IN_194, ImgReg5IN_193, ImgReg5IN_192, 
      ImgReg5IN_191, ImgReg5IN_190, ImgReg5IN_189, ImgReg5IN_188, 
      ImgReg5IN_187, ImgReg5IN_186, ImgReg5IN_185, ImgReg5IN_184, 
      ImgReg5IN_183, ImgReg5IN_182, ImgReg5IN_181, ImgReg5IN_180, 
      ImgReg5IN_179, ImgReg5IN_178, ImgReg5IN_177, ImgReg5IN_176, 
      ImgReg5IN_175, ImgReg5IN_174, ImgReg5IN_173, ImgReg5IN_172, 
      ImgReg5IN_171, ImgReg5IN_170, ImgReg5IN_169, ImgReg5IN_168, 
      ImgReg5IN_167, ImgReg5IN_166, ImgReg5IN_165, ImgReg5IN_164, 
      ImgReg5IN_163, ImgReg5IN_162, ImgReg5IN_161, ImgReg5IN_160, 
      ImgReg5IN_159, ImgReg5IN_158, ImgReg5IN_157, ImgReg5IN_156, 
      ImgReg5IN_155, ImgReg5IN_154, ImgReg5IN_153, ImgReg5IN_152, 
      ImgReg5IN_151, ImgReg5IN_150, ImgReg5IN_149, ImgReg5IN_148, 
      ImgReg5IN_147, ImgReg5IN_146, ImgReg5IN_145, ImgReg5IN_144, 
      ImgReg5IN_143, ImgReg5IN_142, ImgReg5IN_141, ImgReg5IN_140, 
      ImgReg5IN_139, ImgReg5IN_138, ImgReg5IN_137, ImgReg5IN_136, 
      ImgReg5IN_135, ImgReg5IN_134, ImgReg5IN_133, ImgReg5IN_132, 
      ImgReg5IN_131, ImgReg5IN_130, ImgReg5IN_129, ImgReg5IN_128, 
      ImgReg5IN_127, ImgReg5IN_126, ImgReg5IN_125, ImgReg5IN_124, 
      ImgReg5IN_123, ImgReg5IN_122, ImgReg5IN_121, ImgReg5IN_120, 
      ImgReg5IN_119, ImgReg5IN_118, ImgReg5IN_117, ImgReg5IN_116, 
      ImgReg5IN_115, ImgReg5IN_114, ImgReg5IN_113, ImgReg5IN_112, 
      ImgReg5IN_111, ImgReg5IN_110, ImgReg5IN_109, ImgReg5IN_108, 
      ImgReg5IN_107, ImgReg5IN_106, ImgReg5IN_105, ImgReg5IN_104, 
      ImgReg5IN_103, ImgReg5IN_102, ImgReg5IN_101, ImgReg5IN_100, 
      ImgReg5IN_99, ImgReg5IN_98, ImgReg5IN_97, ImgReg5IN_96, ImgReg5IN_95, 
      ImgReg5IN_94, ImgReg5IN_93, ImgReg5IN_92, ImgReg5IN_91, ImgReg5IN_90, 
      ImgReg5IN_89, ImgReg5IN_88, ImgReg5IN_87, ImgReg5IN_86, ImgReg5IN_85, 
      ImgReg5IN_84, ImgReg5IN_83, ImgReg5IN_82, ImgReg5IN_81, ImgReg5IN_80, 
      ImgReg5IN_79, ImgReg5IN_78, ImgReg5IN_77, ImgReg5IN_76, ImgReg5IN_75, 
      ImgReg5IN_74, ImgReg5IN_73, ImgReg5IN_72, ImgReg5IN_71, ImgReg5IN_70, 
      ImgReg5IN_69, ImgReg5IN_68, ImgReg5IN_67, ImgReg5IN_66, ImgReg5IN_65, 
      ImgReg5IN_64, ImgReg5IN_63, ImgReg5IN_62, ImgReg5IN_61, ImgReg5IN_60, 
      ImgReg5IN_59, ImgReg5IN_58, ImgReg5IN_57, ImgReg5IN_56, ImgReg5IN_55, 
      ImgReg5IN_54, ImgReg5IN_53, ImgReg5IN_52, ImgReg5IN_51, ImgReg5IN_50, 
      ImgReg5IN_49, ImgReg5IN_48, ImgReg5IN_47, ImgReg5IN_46, ImgReg5IN_45, 
      ImgReg5IN_44, ImgReg5IN_43, ImgReg5IN_42, ImgReg5IN_41, ImgReg5IN_40, 
      ImgReg5IN_39, ImgReg5IN_38, ImgReg5IN_37, ImgReg5IN_36, ImgReg5IN_35, 
      ImgReg5IN_34, ImgReg5IN_33, ImgReg5IN_32, ImgReg5IN_31, ImgReg5IN_30, 
      ImgReg5IN_29, ImgReg5IN_28, ImgReg5IN_27, ImgReg5IN_26, ImgReg5IN_25, 
      ImgReg5IN_24, ImgReg5IN_23, ImgReg5IN_22, ImgReg5IN_21, ImgReg5IN_20, 
      ImgReg5IN_19, ImgReg5IN_18, ImgReg5IN_17, ImgReg5IN_16, ImgReg5IN_15, 
      ImgReg5IN_14, ImgReg5IN_13, ImgReg5IN_12, ImgReg5IN_11, ImgReg5IN_10, 
      ImgReg5IN_9, ImgReg5IN_8, ImgReg5IN_7, ImgReg5IN_6, ImgReg5IN_5, 
      ImgReg5IN_4, ImgReg5IN_3, ImgReg5IN_2, ImgReg5IN_1, ImgReg5IN_0, 
      TriAddEn, IndRst, cReset, cEnable, TriImgRegEn, TriImgLeftEn, PWR, 
      firstOperand_15, nx2, nx20, nx34, NOT_ImgIndic_0, nx23568, nx23573, 
      nx23580, nx23583, nx23592, nx23594, nx23596, nx23598, nx23600, nx23604, 
      nx23606, nx23608, nx23610, nx23612, nx23616, nx23618, nx23620, nx23622, 
      nx23624, nx23628, nx23630, nx23632, nx23634, nx23636, nx23640, nx23642, 
      nx23644, nx23646, nx23648, nx23652, nx23654, nx23656, nx23658, nx23660, 
      nx23664, nx23666, nx23668, nx23670, nx23672, nx23674, nx23676, nx23678, 
      nx23680, nx23682, nx23684, nx23686, nx23688, nx23690, nx23692, nx23694, 
      nx23696, nx23698, nx23700, nx23702, nx23704, nx23706, nx23708, nx23710, 
      nx23712, nx23716, nx23718, nx23720, nx23722, nx23724, nx23726, nx23728, 
      nx23730, nx23732, nx23734, nx23736, nx23738, nx23740, nx23742, nx23744, 
      nx23746, nx23748, nx23750, nx23752, nx23754, nx23756, nx23758, nx23760, 
      nx23762, nx23764, nx23766, nx23768, nx23770, nx23772, nx23774, nx23776, 
      nx23778, nx23780, nx23786, nx23788, nx23790, nx23792, nx23794, nx23796, 
      nx23798, nx23800, nx23802, nx23804, nx23806, nx23808, nx23810, nx23812, 
      nx23814, nx23816, nx23818, nx23820, nx23822, nx23824, nx23828, nx23830, 
      nx23832, nx23834, nx23836, nx23838, nx23840, nx23842, nx23844, nx23846, 
      nx23848, nx23850, nx23852, nx23854, nx23856, nx23858, nx23860, nx23862, 
      nx23864, nx23866, nx23868, nx23870, nx23872, nx23874, nx23876, nx23878, 
      nx23880, nx23882, nx23884, nx23886, nx23888, nx23890, nx23892, nx23894, 
      nx23896, nx23898, nx23900, nx23902, nx23904, nx23906, nx23908, nx23910, 
      nx23912, nx23914, nx23916, nx23918, nx23920, nx23922, nx23924, nx23926, 
      nx23928, nx23930, nx23932, nx23934, nx23936, nx23938, nx23940, nx23942, 
      nx23944, nx23946, nx23948, nx23950, nx23952, nx23954, nx23956, nx23958, 
      nx23960, nx23962, nx23964, nx23966, nx23968, nx23970, nx23972, nx23974, 
      nx23976, nx23978, nx23980, nx23982, nx23984, nx23986, nx23988, nx23990, 
      nx23992, nx23994, nx23996, nx23998, nx24000, nx24002, nx24004, nx24006, 
      nx24008, nx24010, nx24012, nx24014, nx24016, nx24018, nx24020, nx24022, 
      nx24024, nx24026, nx24028, nx24030, nx24032, nx24038, nx24040: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (3 downto 0 );

begin
   OutputImg0(447) <= OutputImg0_447_EXMPLR ;
   OutputImg0(446) <= OutputImg0_446_EXMPLR ;
   OutputImg0(445) <= OutputImg0_445_EXMPLR ;
   OutputImg0(444) <= OutputImg0_444_EXMPLR ;
   OutputImg0(443) <= OutputImg0_443_EXMPLR ;
   OutputImg0(442) <= OutputImg0_442_EXMPLR ;
   OutputImg0(441) <= OutputImg0_441_EXMPLR ;
   OutputImg0(440) <= OutputImg0_440_EXMPLR ;
   OutputImg0(439) <= OutputImg0_439_EXMPLR ;
   OutputImg0(438) <= OutputImg0_438_EXMPLR ;
   OutputImg0(437) <= OutputImg0_437_EXMPLR ;
   OutputImg0(436) <= OutputImg0_436_EXMPLR ;
   OutputImg0(435) <= OutputImg0_435_EXMPLR ;
   OutputImg0(434) <= OutputImg0_434_EXMPLR ;
   OutputImg0(433) <= OutputImg0_433_EXMPLR ;
   OutputImg0(432) <= OutputImg0_432_EXMPLR ;
   OutputImg0(431) <= OutputImg0_431_EXMPLR ;
   OutputImg0(430) <= OutputImg0_430_EXMPLR ;
   OutputImg0(429) <= OutputImg0_429_EXMPLR ;
   OutputImg0(428) <= OutputImg0_428_EXMPLR ;
   OutputImg0(427) <= OutputImg0_427_EXMPLR ;
   OutputImg0(426) <= OutputImg0_426_EXMPLR ;
   OutputImg0(425) <= OutputImg0_425_EXMPLR ;
   OutputImg0(424) <= OutputImg0_424_EXMPLR ;
   OutputImg0(423) <= OutputImg0_423_EXMPLR ;
   OutputImg0(422) <= OutputImg0_422_EXMPLR ;
   OutputImg0(421) <= OutputImg0_421_EXMPLR ;
   OutputImg0(420) <= OutputImg0_420_EXMPLR ;
   OutputImg0(419) <= OutputImg0_419_EXMPLR ;
   OutputImg0(418) <= OutputImg0_418_EXMPLR ;
   OutputImg0(417) <= OutputImg0_417_EXMPLR ;
   OutputImg0(416) <= OutputImg0_416_EXMPLR ;
   OutputImg0(415) <= OutputImg0_415_EXMPLR ;
   OutputImg0(414) <= OutputImg0_414_EXMPLR ;
   OutputImg0(413) <= OutputImg0_413_EXMPLR ;
   OutputImg0(412) <= OutputImg0_412_EXMPLR ;
   OutputImg0(411) <= OutputImg0_411_EXMPLR ;
   OutputImg0(410) <= OutputImg0_410_EXMPLR ;
   OutputImg0(409) <= OutputImg0_409_EXMPLR ;
   OutputImg0(408) <= OutputImg0_408_EXMPLR ;
   OutputImg0(407) <= OutputImg0_407_EXMPLR ;
   OutputImg0(406) <= OutputImg0_406_EXMPLR ;
   OutputImg0(405) <= OutputImg0_405_EXMPLR ;
   OutputImg0(404) <= OutputImg0_404_EXMPLR ;
   OutputImg0(403) <= OutputImg0_403_EXMPLR ;
   OutputImg0(402) <= OutputImg0_402_EXMPLR ;
   OutputImg0(401) <= OutputImg0_401_EXMPLR ;
   OutputImg0(400) <= OutputImg0_400_EXMPLR ;
   OutputImg0(399) <= OutputImg0_399_EXMPLR ;
   OutputImg0(398) <= OutputImg0_398_EXMPLR ;
   OutputImg0(397) <= OutputImg0_397_EXMPLR ;
   OutputImg0(396) <= OutputImg0_396_EXMPLR ;
   OutputImg0(395) <= OutputImg0_395_EXMPLR ;
   OutputImg0(394) <= OutputImg0_394_EXMPLR ;
   OutputImg0(393) <= OutputImg0_393_EXMPLR ;
   OutputImg0(392) <= OutputImg0_392_EXMPLR ;
   OutputImg0(391) <= OutputImg0_391_EXMPLR ;
   OutputImg0(390) <= OutputImg0_390_EXMPLR ;
   OutputImg0(389) <= OutputImg0_389_EXMPLR ;
   OutputImg0(388) <= OutputImg0_388_EXMPLR ;
   OutputImg0(387) <= OutputImg0_387_EXMPLR ;
   OutputImg0(386) <= OutputImg0_386_EXMPLR ;
   OutputImg0(385) <= OutputImg0_385_EXMPLR ;
   OutputImg0(384) <= OutputImg0_384_EXMPLR ;
   OutputImg0(383) <= OutputImg0_383_EXMPLR ;
   OutputImg0(382) <= OutputImg0_382_EXMPLR ;
   OutputImg0(381) <= OutputImg0_381_EXMPLR ;
   OutputImg0(380) <= OutputImg0_380_EXMPLR ;
   OutputImg0(379) <= OutputImg0_379_EXMPLR ;
   OutputImg0(378) <= OutputImg0_378_EXMPLR ;
   OutputImg0(377) <= OutputImg0_377_EXMPLR ;
   OutputImg0(376) <= OutputImg0_376_EXMPLR ;
   OutputImg0(375) <= OutputImg0_375_EXMPLR ;
   OutputImg0(374) <= OutputImg0_374_EXMPLR ;
   OutputImg0(373) <= OutputImg0_373_EXMPLR ;
   OutputImg0(372) <= OutputImg0_372_EXMPLR ;
   OutputImg0(371) <= OutputImg0_371_EXMPLR ;
   OutputImg0(370) <= OutputImg0_370_EXMPLR ;
   OutputImg0(369) <= OutputImg0_369_EXMPLR ;
   OutputImg0(368) <= OutputImg0_368_EXMPLR ;
   OutputImg0(367) <= OutputImg0_367_EXMPLR ;
   OutputImg0(366) <= OutputImg0_366_EXMPLR ;
   OutputImg0(365) <= OutputImg0_365_EXMPLR ;
   OutputImg0(364) <= OutputImg0_364_EXMPLR ;
   OutputImg0(363) <= OutputImg0_363_EXMPLR ;
   OutputImg0(362) <= OutputImg0_362_EXMPLR ;
   OutputImg0(361) <= OutputImg0_361_EXMPLR ;
   OutputImg0(360) <= OutputImg0_360_EXMPLR ;
   OutputImg0(359) <= OutputImg0_359_EXMPLR ;
   OutputImg0(358) <= OutputImg0_358_EXMPLR ;
   OutputImg0(357) <= OutputImg0_357_EXMPLR ;
   OutputImg0(356) <= OutputImg0_356_EXMPLR ;
   OutputImg0(355) <= OutputImg0_355_EXMPLR ;
   OutputImg0(354) <= OutputImg0_354_EXMPLR ;
   OutputImg0(353) <= OutputImg0_353_EXMPLR ;
   OutputImg0(352) <= OutputImg0_352_EXMPLR ;
   OutputImg0(351) <= OutputImg0_351_EXMPLR ;
   OutputImg0(350) <= OutputImg0_350_EXMPLR ;
   OutputImg0(349) <= OutputImg0_349_EXMPLR ;
   OutputImg0(348) <= OutputImg0_348_EXMPLR ;
   OutputImg0(347) <= OutputImg0_347_EXMPLR ;
   OutputImg0(346) <= OutputImg0_346_EXMPLR ;
   OutputImg0(345) <= OutputImg0_345_EXMPLR ;
   OutputImg0(344) <= OutputImg0_344_EXMPLR ;
   OutputImg0(343) <= OutputImg0_343_EXMPLR ;
   OutputImg0(342) <= OutputImg0_342_EXMPLR ;
   OutputImg0(341) <= OutputImg0_341_EXMPLR ;
   OutputImg0(340) <= OutputImg0_340_EXMPLR ;
   OutputImg0(339) <= OutputImg0_339_EXMPLR ;
   OutputImg0(338) <= OutputImg0_338_EXMPLR ;
   OutputImg0(337) <= OutputImg0_337_EXMPLR ;
   OutputImg0(336) <= OutputImg0_336_EXMPLR ;
   OutputImg0(335) <= OutputImg0_335_EXMPLR ;
   OutputImg0(334) <= OutputImg0_334_EXMPLR ;
   OutputImg0(333) <= OutputImg0_333_EXMPLR ;
   OutputImg0(332) <= OutputImg0_332_EXMPLR ;
   OutputImg0(331) <= OutputImg0_331_EXMPLR ;
   OutputImg0(330) <= OutputImg0_330_EXMPLR ;
   OutputImg0(329) <= OutputImg0_329_EXMPLR ;
   OutputImg0(328) <= OutputImg0_328_EXMPLR ;
   OutputImg0(327) <= OutputImg0_327_EXMPLR ;
   OutputImg0(326) <= OutputImg0_326_EXMPLR ;
   OutputImg0(325) <= OutputImg0_325_EXMPLR ;
   OutputImg0(324) <= OutputImg0_324_EXMPLR ;
   OutputImg0(323) <= OutputImg0_323_EXMPLR ;
   OutputImg0(322) <= OutputImg0_322_EXMPLR ;
   OutputImg0(321) <= OutputImg0_321_EXMPLR ;
   OutputImg0(320) <= OutputImg0_320_EXMPLR ;
   OutputImg0(319) <= OutputImg0_319_EXMPLR ;
   OutputImg0(318) <= OutputImg0_318_EXMPLR ;
   OutputImg0(317) <= OutputImg0_317_EXMPLR ;
   OutputImg0(316) <= OutputImg0_316_EXMPLR ;
   OutputImg0(315) <= OutputImg0_315_EXMPLR ;
   OutputImg0(314) <= OutputImg0_314_EXMPLR ;
   OutputImg0(313) <= OutputImg0_313_EXMPLR ;
   OutputImg0(312) <= OutputImg0_312_EXMPLR ;
   OutputImg0(311) <= OutputImg0_311_EXMPLR ;
   OutputImg0(310) <= OutputImg0_310_EXMPLR ;
   OutputImg0(309) <= OutputImg0_309_EXMPLR ;
   OutputImg0(308) <= OutputImg0_308_EXMPLR ;
   OutputImg0(307) <= OutputImg0_307_EXMPLR ;
   OutputImg0(306) <= OutputImg0_306_EXMPLR ;
   OutputImg0(305) <= OutputImg0_305_EXMPLR ;
   OutputImg0(304) <= OutputImg0_304_EXMPLR ;
   OutputImg0(303) <= OutputImg0_303_EXMPLR ;
   OutputImg0(302) <= OutputImg0_302_EXMPLR ;
   OutputImg0(301) <= OutputImg0_301_EXMPLR ;
   OutputImg0(300) <= OutputImg0_300_EXMPLR ;
   OutputImg0(299) <= OutputImg0_299_EXMPLR ;
   OutputImg0(298) <= OutputImg0_298_EXMPLR ;
   OutputImg0(297) <= OutputImg0_297_EXMPLR ;
   OutputImg0(296) <= OutputImg0_296_EXMPLR ;
   OutputImg0(295) <= OutputImg0_295_EXMPLR ;
   OutputImg0(294) <= OutputImg0_294_EXMPLR ;
   OutputImg0(293) <= OutputImg0_293_EXMPLR ;
   OutputImg0(292) <= OutputImg0_292_EXMPLR ;
   OutputImg0(291) <= OutputImg0_291_EXMPLR ;
   OutputImg0(290) <= OutputImg0_290_EXMPLR ;
   OutputImg0(289) <= OutputImg0_289_EXMPLR ;
   OutputImg0(288) <= OutputImg0_288_EXMPLR ;
   OutputImg0(287) <= OutputImg0_287_EXMPLR ;
   OutputImg0(286) <= OutputImg0_286_EXMPLR ;
   OutputImg0(285) <= OutputImg0_285_EXMPLR ;
   OutputImg0(284) <= OutputImg0_284_EXMPLR ;
   OutputImg0(283) <= OutputImg0_283_EXMPLR ;
   OutputImg0(282) <= OutputImg0_282_EXMPLR ;
   OutputImg0(281) <= OutputImg0_281_EXMPLR ;
   OutputImg0(280) <= OutputImg0_280_EXMPLR ;
   OutputImg0(279) <= OutputImg0_279_EXMPLR ;
   OutputImg0(278) <= OutputImg0_278_EXMPLR ;
   OutputImg0(277) <= OutputImg0_277_EXMPLR ;
   OutputImg0(276) <= OutputImg0_276_EXMPLR ;
   OutputImg0(275) <= OutputImg0_275_EXMPLR ;
   OutputImg0(274) <= OutputImg0_274_EXMPLR ;
   OutputImg0(273) <= OutputImg0_273_EXMPLR ;
   OutputImg0(272) <= OutputImg0_272_EXMPLR ;
   OutputImg0(271) <= OutputImg0_271_EXMPLR ;
   OutputImg0(270) <= OutputImg0_270_EXMPLR ;
   OutputImg0(269) <= OutputImg0_269_EXMPLR ;
   OutputImg0(268) <= OutputImg0_268_EXMPLR ;
   OutputImg0(267) <= OutputImg0_267_EXMPLR ;
   OutputImg0(266) <= OutputImg0_266_EXMPLR ;
   OutputImg0(265) <= OutputImg0_265_EXMPLR ;
   OutputImg0(264) <= OutputImg0_264_EXMPLR ;
   OutputImg0(263) <= OutputImg0_263_EXMPLR ;
   OutputImg0(262) <= OutputImg0_262_EXMPLR ;
   OutputImg0(261) <= OutputImg0_261_EXMPLR ;
   OutputImg0(260) <= OutputImg0_260_EXMPLR ;
   OutputImg0(259) <= OutputImg0_259_EXMPLR ;
   OutputImg0(258) <= OutputImg0_258_EXMPLR ;
   OutputImg0(257) <= OutputImg0_257_EXMPLR ;
   OutputImg0(256) <= OutputImg0_256_EXMPLR ;
   OutputImg0(255) <= OutputImg0_255_EXMPLR ;
   OutputImg0(254) <= OutputImg0_254_EXMPLR ;
   OutputImg0(253) <= OutputImg0_253_EXMPLR ;
   OutputImg0(252) <= OutputImg0_252_EXMPLR ;
   OutputImg0(251) <= OutputImg0_251_EXMPLR ;
   OutputImg0(250) <= OutputImg0_250_EXMPLR ;
   OutputImg0(249) <= OutputImg0_249_EXMPLR ;
   OutputImg0(248) <= OutputImg0_248_EXMPLR ;
   OutputImg0(247) <= OutputImg0_247_EXMPLR ;
   OutputImg0(246) <= OutputImg0_246_EXMPLR ;
   OutputImg0(245) <= OutputImg0_245_EXMPLR ;
   OutputImg0(244) <= OutputImg0_244_EXMPLR ;
   OutputImg0(243) <= OutputImg0_243_EXMPLR ;
   OutputImg0(242) <= OutputImg0_242_EXMPLR ;
   OutputImg0(241) <= OutputImg0_241_EXMPLR ;
   OutputImg0(240) <= OutputImg0_240_EXMPLR ;
   OutputImg0(239) <= OutputImg0_239_EXMPLR ;
   OutputImg0(238) <= OutputImg0_238_EXMPLR ;
   OutputImg0(237) <= OutputImg0_237_EXMPLR ;
   OutputImg0(236) <= OutputImg0_236_EXMPLR ;
   OutputImg0(235) <= OutputImg0_235_EXMPLR ;
   OutputImg0(234) <= OutputImg0_234_EXMPLR ;
   OutputImg0(233) <= OutputImg0_233_EXMPLR ;
   OutputImg0(232) <= OutputImg0_232_EXMPLR ;
   OutputImg0(231) <= OutputImg0_231_EXMPLR ;
   OutputImg0(230) <= OutputImg0_230_EXMPLR ;
   OutputImg0(229) <= OutputImg0_229_EXMPLR ;
   OutputImg0(228) <= OutputImg0_228_EXMPLR ;
   OutputImg0(227) <= OutputImg0_227_EXMPLR ;
   OutputImg0(226) <= OutputImg0_226_EXMPLR ;
   OutputImg0(225) <= OutputImg0_225_EXMPLR ;
   OutputImg0(224) <= OutputImg0_224_EXMPLR ;
   OutputImg0(223) <= OutputImg0_223_EXMPLR ;
   OutputImg0(222) <= OutputImg0_222_EXMPLR ;
   OutputImg0(221) <= OutputImg0_221_EXMPLR ;
   OutputImg0(220) <= OutputImg0_220_EXMPLR ;
   OutputImg0(219) <= OutputImg0_219_EXMPLR ;
   OutputImg0(218) <= OutputImg0_218_EXMPLR ;
   OutputImg0(217) <= OutputImg0_217_EXMPLR ;
   OutputImg0(216) <= OutputImg0_216_EXMPLR ;
   OutputImg0(215) <= OutputImg0_215_EXMPLR ;
   OutputImg0(214) <= OutputImg0_214_EXMPLR ;
   OutputImg0(213) <= OutputImg0_213_EXMPLR ;
   OutputImg0(212) <= OutputImg0_212_EXMPLR ;
   OutputImg0(211) <= OutputImg0_211_EXMPLR ;
   OutputImg0(210) <= OutputImg0_210_EXMPLR ;
   OutputImg0(209) <= OutputImg0_209_EXMPLR ;
   OutputImg0(208) <= OutputImg0_208_EXMPLR ;
   OutputImg0(207) <= OutputImg0_207_EXMPLR ;
   OutputImg0(206) <= OutputImg0_206_EXMPLR ;
   OutputImg0(205) <= OutputImg0_205_EXMPLR ;
   OutputImg0(204) <= OutputImg0_204_EXMPLR ;
   OutputImg0(203) <= OutputImg0_203_EXMPLR ;
   OutputImg0(202) <= OutputImg0_202_EXMPLR ;
   OutputImg0(201) <= OutputImg0_201_EXMPLR ;
   OutputImg0(200) <= OutputImg0_200_EXMPLR ;
   OutputImg0(199) <= OutputImg0_199_EXMPLR ;
   OutputImg0(198) <= OutputImg0_198_EXMPLR ;
   OutputImg0(197) <= OutputImg0_197_EXMPLR ;
   OutputImg0(196) <= OutputImg0_196_EXMPLR ;
   OutputImg0(195) <= OutputImg0_195_EXMPLR ;
   OutputImg0(194) <= OutputImg0_194_EXMPLR ;
   OutputImg0(193) <= OutputImg0_193_EXMPLR ;
   OutputImg0(192) <= OutputImg0_192_EXMPLR ;
   OutputImg0(191) <= OutputImg0_191_EXMPLR ;
   OutputImg0(190) <= OutputImg0_190_EXMPLR ;
   OutputImg0(189) <= OutputImg0_189_EXMPLR ;
   OutputImg0(188) <= OutputImg0_188_EXMPLR ;
   OutputImg0(187) <= OutputImg0_187_EXMPLR ;
   OutputImg0(186) <= OutputImg0_186_EXMPLR ;
   OutputImg0(185) <= OutputImg0_185_EXMPLR ;
   OutputImg0(184) <= OutputImg0_184_EXMPLR ;
   OutputImg0(183) <= OutputImg0_183_EXMPLR ;
   OutputImg0(182) <= OutputImg0_182_EXMPLR ;
   OutputImg0(181) <= OutputImg0_181_EXMPLR ;
   OutputImg0(180) <= OutputImg0_180_EXMPLR ;
   OutputImg0(179) <= OutputImg0_179_EXMPLR ;
   OutputImg0(178) <= OutputImg0_178_EXMPLR ;
   OutputImg0(177) <= OutputImg0_177_EXMPLR ;
   OutputImg0(176) <= OutputImg0_176_EXMPLR ;
   OutputImg0(175) <= OutputImg0_175_EXMPLR ;
   OutputImg0(174) <= OutputImg0_174_EXMPLR ;
   OutputImg0(173) <= OutputImg0_173_EXMPLR ;
   OutputImg0(172) <= OutputImg0_172_EXMPLR ;
   OutputImg0(171) <= OutputImg0_171_EXMPLR ;
   OutputImg0(170) <= OutputImg0_170_EXMPLR ;
   OutputImg0(169) <= OutputImg0_169_EXMPLR ;
   OutputImg0(168) <= OutputImg0_168_EXMPLR ;
   OutputImg0(167) <= OutputImg0_167_EXMPLR ;
   OutputImg0(166) <= OutputImg0_166_EXMPLR ;
   OutputImg0(165) <= OutputImg0_165_EXMPLR ;
   OutputImg0(164) <= OutputImg0_164_EXMPLR ;
   OutputImg0(163) <= OutputImg0_163_EXMPLR ;
   OutputImg0(162) <= OutputImg0_162_EXMPLR ;
   OutputImg0(161) <= OutputImg0_161_EXMPLR ;
   OutputImg0(160) <= OutputImg0_160_EXMPLR ;
   OutputImg0(159) <= OutputImg0_159_EXMPLR ;
   OutputImg0(158) <= OutputImg0_158_EXMPLR ;
   OutputImg0(157) <= OutputImg0_157_EXMPLR ;
   OutputImg0(156) <= OutputImg0_156_EXMPLR ;
   OutputImg0(155) <= OutputImg0_155_EXMPLR ;
   OutputImg0(154) <= OutputImg0_154_EXMPLR ;
   OutputImg0(153) <= OutputImg0_153_EXMPLR ;
   OutputImg0(152) <= OutputImg0_152_EXMPLR ;
   OutputImg0(151) <= OutputImg0_151_EXMPLR ;
   OutputImg0(150) <= OutputImg0_150_EXMPLR ;
   OutputImg0(149) <= OutputImg0_149_EXMPLR ;
   OutputImg0(148) <= OutputImg0_148_EXMPLR ;
   OutputImg0(147) <= OutputImg0_147_EXMPLR ;
   OutputImg0(146) <= OutputImg0_146_EXMPLR ;
   OutputImg0(145) <= OutputImg0_145_EXMPLR ;
   OutputImg0(144) <= OutputImg0_144_EXMPLR ;
   OutputImg0(143) <= OutputImg0_143_EXMPLR ;
   OutputImg0(142) <= OutputImg0_142_EXMPLR ;
   OutputImg0(141) <= OutputImg0_141_EXMPLR ;
   OutputImg0(140) <= OutputImg0_140_EXMPLR ;
   OutputImg0(139) <= OutputImg0_139_EXMPLR ;
   OutputImg0(138) <= OutputImg0_138_EXMPLR ;
   OutputImg0(137) <= OutputImg0_137_EXMPLR ;
   OutputImg0(136) <= OutputImg0_136_EXMPLR ;
   OutputImg0(135) <= OutputImg0_135_EXMPLR ;
   OutputImg0(134) <= OutputImg0_134_EXMPLR ;
   OutputImg0(133) <= OutputImg0_133_EXMPLR ;
   OutputImg0(132) <= OutputImg0_132_EXMPLR ;
   OutputImg0(131) <= OutputImg0_131_EXMPLR ;
   OutputImg0(130) <= OutputImg0_130_EXMPLR ;
   OutputImg0(129) <= OutputImg0_129_EXMPLR ;
   OutputImg0(128) <= OutputImg0_128_EXMPLR ;
   OutputImg0(127) <= OutputImg0_127_EXMPLR ;
   OutputImg0(126) <= OutputImg0_126_EXMPLR ;
   OutputImg0(125) <= OutputImg0_125_EXMPLR ;
   OutputImg0(124) <= OutputImg0_124_EXMPLR ;
   OutputImg0(123) <= OutputImg0_123_EXMPLR ;
   OutputImg0(122) <= OutputImg0_122_EXMPLR ;
   OutputImg0(121) <= OutputImg0_121_EXMPLR ;
   OutputImg0(120) <= OutputImg0_120_EXMPLR ;
   OutputImg0(119) <= OutputImg0_119_EXMPLR ;
   OutputImg0(118) <= OutputImg0_118_EXMPLR ;
   OutputImg0(117) <= OutputImg0_117_EXMPLR ;
   OutputImg0(116) <= OutputImg0_116_EXMPLR ;
   OutputImg0(115) <= OutputImg0_115_EXMPLR ;
   OutputImg0(114) <= OutputImg0_114_EXMPLR ;
   OutputImg0(113) <= OutputImg0_113_EXMPLR ;
   OutputImg0(112) <= OutputImg0_112_EXMPLR ;
   OutputImg0(111) <= OutputImg0_111_EXMPLR ;
   OutputImg0(110) <= OutputImg0_110_EXMPLR ;
   OutputImg0(109) <= OutputImg0_109_EXMPLR ;
   OutputImg0(108) <= OutputImg0_108_EXMPLR ;
   OutputImg0(107) <= OutputImg0_107_EXMPLR ;
   OutputImg0(106) <= OutputImg0_106_EXMPLR ;
   OutputImg0(105) <= OutputImg0_105_EXMPLR ;
   OutputImg0(104) <= OutputImg0_104_EXMPLR ;
   OutputImg0(103) <= OutputImg0_103_EXMPLR ;
   OutputImg0(102) <= OutputImg0_102_EXMPLR ;
   OutputImg0(101) <= OutputImg0_101_EXMPLR ;
   OutputImg0(100) <= OutputImg0_100_EXMPLR ;
   OutputImg0(99) <= OutputImg0_99_EXMPLR ;
   OutputImg0(98) <= OutputImg0_98_EXMPLR ;
   OutputImg0(97) <= OutputImg0_97_EXMPLR ;
   OutputImg0(96) <= OutputImg0_96_EXMPLR ;
   OutputImg0(95) <= OutputImg0_95_EXMPLR ;
   OutputImg0(94) <= OutputImg0_94_EXMPLR ;
   OutputImg0(93) <= OutputImg0_93_EXMPLR ;
   OutputImg0(92) <= OutputImg0_92_EXMPLR ;
   OutputImg0(91) <= OutputImg0_91_EXMPLR ;
   OutputImg0(90) <= OutputImg0_90_EXMPLR ;
   OutputImg0(89) <= OutputImg0_89_EXMPLR ;
   OutputImg0(88) <= OutputImg0_88_EXMPLR ;
   OutputImg0(87) <= OutputImg0_87_EXMPLR ;
   OutputImg0(86) <= OutputImg0_86_EXMPLR ;
   OutputImg0(85) <= OutputImg0_85_EXMPLR ;
   OutputImg0(84) <= OutputImg0_84_EXMPLR ;
   OutputImg0(83) <= OutputImg0_83_EXMPLR ;
   OutputImg0(82) <= OutputImg0_82_EXMPLR ;
   OutputImg0(81) <= OutputImg0_81_EXMPLR ;
   OutputImg0(80) <= OutputImg0_80_EXMPLR ;
   OutputImg0(79) <= OutputImg0_79_EXMPLR ;
   OutputImg0(78) <= OutputImg0_78_EXMPLR ;
   OutputImg0(77) <= OutputImg0_77_EXMPLR ;
   OutputImg0(76) <= OutputImg0_76_EXMPLR ;
   OutputImg0(75) <= OutputImg0_75_EXMPLR ;
   OutputImg0(74) <= OutputImg0_74_EXMPLR ;
   OutputImg0(73) <= OutputImg0_73_EXMPLR ;
   OutputImg0(72) <= OutputImg0_72_EXMPLR ;
   OutputImg0(71) <= OutputImg0_71_EXMPLR ;
   OutputImg0(70) <= OutputImg0_70_EXMPLR ;
   OutputImg0(69) <= OutputImg0_69_EXMPLR ;
   OutputImg0(68) <= OutputImg0_68_EXMPLR ;
   OutputImg0(67) <= OutputImg0_67_EXMPLR ;
   OutputImg0(66) <= OutputImg0_66_EXMPLR ;
   OutputImg0(65) <= OutputImg0_65_EXMPLR ;
   OutputImg0(64) <= OutputImg0_64_EXMPLR ;
   OutputImg0(63) <= OutputImg0_63_EXMPLR ;
   OutputImg0(62) <= OutputImg0_62_EXMPLR ;
   OutputImg0(61) <= OutputImg0_61_EXMPLR ;
   OutputImg0(60) <= OutputImg0_60_EXMPLR ;
   OutputImg0(59) <= OutputImg0_59_EXMPLR ;
   OutputImg0(58) <= OutputImg0_58_EXMPLR ;
   OutputImg0(57) <= OutputImg0_57_EXMPLR ;
   OutputImg0(56) <= OutputImg0_56_EXMPLR ;
   OutputImg0(55) <= OutputImg0_55_EXMPLR ;
   OutputImg0(54) <= OutputImg0_54_EXMPLR ;
   OutputImg0(53) <= OutputImg0_53_EXMPLR ;
   OutputImg0(52) <= OutputImg0_52_EXMPLR ;
   OutputImg0(51) <= OutputImg0_51_EXMPLR ;
   OutputImg0(50) <= OutputImg0_50_EXMPLR ;
   OutputImg0(49) <= OutputImg0_49_EXMPLR ;
   OutputImg0(48) <= OutputImg0_48_EXMPLR ;
   OutputImg0(47) <= OutputImg0_47_EXMPLR ;
   OutputImg0(46) <= OutputImg0_46_EXMPLR ;
   OutputImg0(45) <= OutputImg0_45_EXMPLR ;
   OutputImg0(44) <= OutputImg0_44_EXMPLR ;
   OutputImg0(43) <= OutputImg0_43_EXMPLR ;
   OutputImg0(42) <= OutputImg0_42_EXMPLR ;
   OutputImg0(41) <= OutputImg0_41_EXMPLR ;
   OutputImg0(40) <= OutputImg0_40_EXMPLR ;
   OutputImg0(39) <= OutputImg0_39_EXMPLR ;
   OutputImg0(38) <= OutputImg0_38_EXMPLR ;
   OutputImg0(37) <= OutputImg0_37_EXMPLR ;
   OutputImg0(36) <= OutputImg0_36_EXMPLR ;
   OutputImg0(35) <= OutputImg0_35_EXMPLR ;
   OutputImg0(34) <= OutputImg0_34_EXMPLR ;
   OutputImg0(33) <= OutputImg0_33_EXMPLR ;
   OutputImg0(32) <= OutputImg0_32_EXMPLR ;
   OutputImg0(31) <= OutputImg0_31_EXMPLR ;
   OutputImg0(30) <= OutputImg0_30_EXMPLR ;
   OutputImg0(29) <= OutputImg0_29_EXMPLR ;
   OutputImg0(28) <= OutputImg0_28_EXMPLR ;
   OutputImg0(27) <= OutputImg0_27_EXMPLR ;
   OutputImg0(26) <= OutputImg0_26_EXMPLR ;
   OutputImg0(25) <= OutputImg0_25_EXMPLR ;
   OutputImg0(24) <= OutputImg0_24_EXMPLR ;
   OutputImg0(23) <= OutputImg0_23_EXMPLR ;
   OutputImg0(22) <= OutputImg0_22_EXMPLR ;
   OutputImg0(21) <= OutputImg0_21_EXMPLR ;
   OutputImg0(20) <= OutputImg0_20_EXMPLR ;
   OutputImg0(19) <= OutputImg0_19_EXMPLR ;
   OutputImg0(18) <= OutputImg0_18_EXMPLR ;
   OutputImg0(17) <= OutputImg0_17_EXMPLR ;
   OutputImg0(16) <= OutputImg0_16_EXMPLR ;
   OutputImg0(15) <= OutputImg0_15_EXMPLR ;
   OutputImg0(14) <= OutputImg0_14_EXMPLR ;
   OutputImg0(13) <= OutputImg0_13_EXMPLR ;
   OutputImg0(12) <= OutputImg0_12_EXMPLR ;
   OutputImg0(11) <= OutputImg0_11_EXMPLR ;
   OutputImg0(10) <= OutputImg0_10_EXMPLR ;
   OutputImg0(9) <= OutputImg0_9_EXMPLR ;
   OutputImg0(8) <= OutputImg0_8_EXMPLR ;
   OutputImg0(7) <= OutputImg0_7_EXMPLR ;
   OutputImg0(6) <= OutputImg0_6_EXMPLR ;
   OutputImg0(5) <= OutputImg0_5_EXMPLR ;
   OutputImg0(4) <= OutputImg0_4_EXMPLR ;
   OutputImg0(3) <= OutputImg0_3_EXMPLR ;
   OutputImg0(2) <= OutputImg0_2_EXMPLR ;
   OutputImg0(1) <= OutputImg0_1_EXMPLR ;
   OutputImg0(0) <= OutputImg0_0_EXMPLR ;
   OutputImg1(447) <= OutputImg1_447_EXMPLR ;
   OutputImg1(446) <= OutputImg1_446_EXMPLR ;
   OutputImg1(445) <= OutputImg1_445_EXMPLR ;
   OutputImg1(444) <= OutputImg1_444_EXMPLR ;
   OutputImg1(443) <= OutputImg1_443_EXMPLR ;
   OutputImg1(442) <= OutputImg1_442_EXMPLR ;
   OutputImg1(441) <= OutputImg1_441_EXMPLR ;
   OutputImg1(440) <= OutputImg1_440_EXMPLR ;
   OutputImg1(439) <= OutputImg1_439_EXMPLR ;
   OutputImg1(438) <= OutputImg1_438_EXMPLR ;
   OutputImg1(437) <= OutputImg1_437_EXMPLR ;
   OutputImg1(436) <= OutputImg1_436_EXMPLR ;
   OutputImg1(435) <= OutputImg1_435_EXMPLR ;
   OutputImg1(434) <= OutputImg1_434_EXMPLR ;
   OutputImg1(433) <= OutputImg1_433_EXMPLR ;
   OutputImg1(432) <= OutputImg1_432_EXMPLR ;
   OutputImg1(431) <= OutputImg1_431_EXMPLR ;
   OutputImg1(430) <= OutputImg1_430_EXMPLR ;
   OutputImg1(429) <= OutputImg1_429_EXMPLR ;
   OutputImg1(428) <= OutputImg1_428_EXMPLR ;
   OutputImg1(427) <= OutputImg1_427_EXMPLR ;
   OutputImg1(426) <= OutputImg1_426_EXMPLR ;
   OutputImg1(425) <= OutputImg1_425_EXMPLR ;
   OutputImg1(424) <= OutputImg1_424_EXMPLR ;
   OutputImg1(423) <= OutputImg1_423_EXMPLR ;
   OutputImg1(422) <= OutputImg1_422_EXMPLR ;
   OutputImg1(421) <= OutputImg1_421_EXMPLR ;
   OutputImg1(420) <= OutputImg1_420_EXMPLR ;
   OutputImg1(419) <= OutputImg1_419_EXMPLR ;
   OutputImg1(418) <= OutputImg1_418_EXMPLR ;
   OutputImg1(417) <= OutputImg1_417_EXMPLR ;
   OutputImg1(416) <= OutputImg1_416_EXMPLR ;
   OutputImg1(415) <= OutputImg1_415_EXMPLR ;
   OutputImg1(414) <= OutputImg1_414_EXMPLR ;
   OutputImg1(413) <= OutputImg1_413_EXMPLR ;
   OutputImg1(412) <= OutputImg1_412_EXMPLR ;
   OutputImg1(411) <= OutputImg1_411_EXMPLR ;
   OutputImg1(410) <= OutputImg1_410_EXMPLR ;
   OutputImg1(409) <= OutputImg1_409_EXMPLR ;
   OutputImg1(408) <= OutputImg1_408_EXMPLR ;
   OutputImg1(407) <= OutputImg1_407_EXMPLR ;
   OutputImg1(406) <= OutputImg1_406_EXMPLR ;
   OutputImg1(405) <= OutputImg1_405_EXMPLR ;
   OutputImg1(404) <= OutputImg1_404_EXMPLR ;
   OutputImg1(403) <= OutputImg1_403_EXMPLR ;
   OutputImg1(402) <= OutputImg1_402_EXMPLR ;
   OutputImg1(401) <= OutputImg1_401_EXMPLR ;
   OutputImg1(400) <= OutputImg1_400_EXMPLR ;
   OutputImg1(399) <= OutputImg1_399_EXMPLR ;
   OutputImg1(398) <= OutputImg1_398_EXMPLR ;
   OutputImg1(397) <= OutputImg1_397_EXMPLR ;
   OutputImg1(396) <= OutputImg1_396_EXMPLR ;
   OutputImg1(395) <= OutputImg1_395_EXMPLR ;
   OutputImg1(394) <= OutputImg1_394_EXMPLR ;
   OutputImg1(393) <= OutputImg1_393_EXMPLR ;
   OutputImg1(392) <= OutputImg1_392_EXMPLR ;
   OutputImg1(391) <= OutputImg1_391_EXMPLR ;
   OutputImg1(390) <= OutputImg1_390_EXMPLR ;
   OutputImg1(389) <= OutputImg1_389_EXMPLR ;
   OutputImg1(388) <= OutputImg1_388_EXMPLR ;
   OutputImg1(387) <= OutputImg1_387_EXMPLR ;
   OutputImg1(386) <= OutputImg1_386_EXMPLR ;
   OutputImg1(385) <= OutputImg1_385_EXMPLR ;
   OutputImg1(384) <= OutputImg1_384_EXMPLR ;
   OutputImg1(383) <= OutputImg1_383_EXMPLR ;
   OutputImg1(382) <= OutputImg1_382_EXMPLR ;
   OutputImg1(381) <= OutputImg1_381_EXMPLR ;
   OutputImg1(380) <= OutputImg1_380_EXMPLR ;
   OutputImg1(379) <= OutputImg1_379_EXMPLR ;
   OutputImg1(378) <= OutputImg1_378_EXMPLR ;
   OutputImg1(377) <= OutputImg1_377_EXMPLR ;
   OutputImg1(376) <= OutputImg1_376_EXMPLR ;
   OutputImg1(375) <= OutputImg1_375_EXMPLR ;
   OutputImg1(374) <= OutputImg1_374_EXMPLR ;
   OutputImg1(373) <= OutputImg1_373_EXMPLR ;
   OutputImg1(372) <= OutputImg1_372_EXMPLR ;
   OutputImg1(371) <= OutputImg1_371_EXMPLR ;
   OutputImg1(370) <= OutputImg1_370_EXMPLR ;
   OutputImg1(369) <= OutputImg1_369_EXMPLR ;
   OutputImg1(368) <= OutputImg1_368_EXMPLR ;
   OutputImg1(367) <= OutputImg1_367_EXMPLR ;
   OutputImg1(366) <= OutputImg1_366_EXMPLR ;
   OutputImg1(365) <= OutputImg1_365_EXMPLR ;
   OutputImg1(364) <= OutputImg1_364_EXMPLR ;
   OutputImg1(363) <= OutputImg1_363_EXMPLR ;
   OutputImg1(362) <= OutputImg1_362_EXMPLR ;
   OutputImg1(361) <= OutputImg1_361_EXMPLR ;
   OutputImg1(360) <= OutputImg1_360_EXMPLR ;
   OutputImg1(359) <= OutputImg1_359_EXMPLR ;
   OutputImg1(358) <= OutputImg1_358_EXMPLR ;
   OutputImg1(357) <= OutputImg1_357_EXMPLR ;
   OutputImg1(356) <= OutputImg1_356_EXMPLR ;
   OutputImg1(355) <= OutputImg1_355_EXMPLR ;
   OutputImg1(354) <= OutputImg1_354_EXMPLR ;
   OutputImg1(353) <= OutputImg1_353_EXMPLR ;
   OutputImg1(352) <= OutputImg1_352_EXMPLR ;
   OutputImg1(351) <= OutputImg1_351_EXMPLR ;
   OutputImg1(350) <= OutputImg1_350_EXMPLR ;
   OutputImg1(349) <= OutputImg1_349_EXMPLR ;
   OutputImg1(348) <= OutputImg1_348_EXMPLR ;
   OutputImg1(347) <= OutputImg1_347_EXMPLR ;
   OutputImg1(346) <= OutputImg1_346_EXMPLR ;
   OutputImg1(345) <= OutputImg1_345_EXMPLR ;
   OutputImg1(344) <= OutputImg1_344_EXMPLR ;
   OutputImg1(343) <= OutputImg1_343_EXMPLR ;
   OutputImg1(342) <= OutputImg1_342_EXMPLR ;
   OutputImg1(341) <= OutputImg1_341_EXMPLR ;
   OutputImg1(340) <= OutputImg1_340_EXMPLR ;
   OutputImg1(339) <= OutputImg1_339_EXMPLR ;
   OutputImg1(338) <= OutputImg1_338_EXMPLR ;
   OutputImg1(337) <= OutputImg1_337_EXMPLR ;
   OutputImg1(336) <= OutputImg1_336_EXMPLR ;
   OutputImg1(335) <= OutputImg1_335_EXMPLR ;
   OutputImg1(334) <= OutputImg1_334_EXMPLR ;
   OutputImg1(333) <= OutputImg1_333_EXMPLR ;
   OutputImg1(332) <= OutputImg1_332_EXMPLR ;
   OutputImg1(331) <= OutputImg1_331_EXMPLR ;
   OutputImg1(330) <= OutputImg1_330_EXMPLR ;
   OutputImg1(329) <= OutputImg1_329_EXMPLR ;
   OutputImg1(328) <= OutputImg1_328_EXMPLR ;
   OutputImg1(327) <= OutputImg1_327_EXMPLR ;
   OutputImg1(326) <= OutputImg1_326_EXMPLR ;
   OutputImg1(325) <= OutputImg1_325_EXMPLR ;
   OutputImg1(324) <= OutputImg1_324_EXMPLR ;
   OutputImg1(323) <= OutputImg1_323_EXMPLR ;
   OutputImg1(322) <= OutputImg1_322_EXMPLR ;
   OutputImg1(321) <= OutputImg1_321_EXMPLR ;
   OutputImg1(320) <= OutputImg1_320_EXMPLR ;
   OutputImg1(319) <= OutputImg1_319_EXMPLR ;
   OutputImg1(318) <= OutputImg1_318_EXMPLR ;
   OutputImg1(317) <= OutputImg1_317_EXMPLR ;
   OutputImg1(316) <= OutputImg1_316_EXMPLR ;
   OutputImg1(315) <= OutputImg1_315_EXMPLR ;
   OutputImg1(314) <= OutputImg1_314_EXMPLR ;
   OutputImg1(313) <= OutputImg1_313_EXMPLR ;
   OutputImg1(312) <= OutputImg1_312_EXMPLR ;
   OutputImg1(311) <= OutputImg1_311_EXMPLR ;
   OutputImg1(310) <= OutputImg1_310_EXMPLR ;
   OutputImg1(309) <= OutputImg1_309_EXMPLR ;
   OutputImg1(308) <= OutputImg1_308_EXMPLR ;
   OutputImg1(307) <= OutputImg1_307_EXMPLR ;
   OutputImg1(306) <= OutputImg1_306_EXMPLR ;
   OutputImg1(305) <= OutputImg1_305_EXMPLR ;
   OutputImg1(304) <= OutputImg1_304_EXMPLR ;
   OutputImg1(303) <= OutputImg1_303_EXMPLR ;
   OutputImg1(302) <= OutputImg1_302_EXMPLR ;
   OutputImg1(301) <= OutputImg1_301_EXMPLR ;
   OutputImg1(300) <= OutputImg1_300_EXMPLR ;
   OutputImg1(299) <= OutputImg1_299_EXMPLR ;
   OutputImg1(298) <= OutputImg1_298_EXMPLR ;
   OutputImg1(297) <= OutputImg1_297_EXMPLR ;
   OutputImg1(296) <= OutputImg1_296_EXMPLR ;
   OutputImg1(295) <= OutputImg1_295_EXMPLR ;
   OutputImg1(294) <= OutputImg1_294_EXMPLR ;
   OutputImg1(293) <= OutputImg1_293_EXMPLR ;
   OutputImg1(292) <= OutputImg1_292_EXMPLR ;
   OutputImg1(291) <= OutputImg1_291_EXMPLR ;
   OutputImg1(290) <= OutputImg1_290_EXMPLR ;
   OutputImg1(289) <= OutputImg1_289_EXMPLR ;
   OutputImg1(288) <= OutputImg1_288_EXMPLR ;
   OutputImg1(287) <= OutputImg1_287_EXMPLR ;
   OutputImg1(286) <= OutputImg1_286_EXMPLR ;
   OutputImg1(285) <= OutputImg1_285_EXMPLR ;
   OutputImg1(284) <= OutputImg1_284_EXMPLR ;
   OutputImg1(283) <= OutputImg1_283_EXMPLR ;
   OutputImg1(282) <= OutputImg1_282_EXMPLR ;
   OutputImg1(281) <= OutputImg1_281_EXMPLR ;
   OutputImg1(280) <= OutputImg1_280_EXMPLR ;
   OutputImg1(279) <= OutputImg1_279_EXMPLR ;
   OutputImg1(278) <= OutputImg1_278_EXMPLR ;
   OutputImg1(277) <= OutputImg1_277_EXMPLR ;
   OutputImg1(276) <= OutputImg1_276_EXMPLR ;
   OutputImg1(275) <= OutputImg1_275_EXMPLR ;
   OutputImg1(274) <= OutputImg1_274_EXMPLR ;
   OutputImg1(273) <= OutputImg1_273_EXMPLR ;
   OutputImg1(272) <= OutputImg1_272_EXMPLR ;
   OutputImg1(271) <= OutputImg1_271_EXMPLR ;
   OutputImg1(270) <= OutputImg1_270_EXMPLR ;
   OutputImg1(269) <= OutputImg1_269_EXMPLR ;
   OutputImg1(268) <= OutputImg1_268_EXMPLR ;
   OutputImg1(267) <= OutputImg1_267_EXMPLR ;
   OutputImg1(266) <= OutputImg1_266_EXMPLR ;
   OutputImg1(265) <= OutputImg1_265_EXMPLR ;
   OutputImg1(264) <= OutputImg1_264_EXMPLR ;
   OutputImg1(263) <= OutputImg1_263_EXMPLR ;
   OutputImg1(262) <= OutputImg1_262_EXMPLR ;
   OutputImg1(261) <= OutputImg1_261_EXMPLR ;
   OutputImg1(260) <= OutputImg1_260_EXMPLR ;
   OutputImg1(259) <= OutputImg1_259_EXMPLR ;
   OutputImg1(258) <= OutputImg1_258_EXMPLR ;
   OutputImg1(257) <= OutputImg1_257_EXMPLR ;
   OutputImg1(256) <= OutputImg1_256_EXMPLR ;
   OutputImg1(255) <= OutputImg1_255_EXMPLR ;
   OutputImg1(254) <= OutputImg1_254_EXMPLR ;
   OutputImg1(253) <= OutputImg1_253_EXMPLR ;
   OutputImg1(252) <= OutputImg1_252_EXMPLR ;
   OutputImg1(251) <= OutputImg1_251_EXMPLR ;
   OutputImg1(250) <= OutputImg1_250_EXMPLR ;
   OutputImg1(249) <= OutputImg1_249_EXMPLR ;
   OutputImg1(248) <= OutputImg1_248_EXMPLR ;
   OutputImg1(247) <= OutputImg1_247_EXMPLR ;
   OutputImg1(246) <= OutputImg1_246_EXMPLR ;
   OutputImg1(245) <= OutputImg1_245_EXMPLR ;
   OutputImg1(244) <= OutputImg1_244_EXMPLR ;
   OutputImg1(243) <= OutputImg1_243_EXMPLR ;
   OutputImg1(242) <= OutputImg1_242_EXMPLR ;
   OutputImg1(241) <= OutputImg1_241_EXMPLR ;
   OutputImg1(240) <= OutputImg1_240_EXMPLR ;
   OutputImg1(239) <= OutputImg1_239_EXMPLR ;
   OutputImg1(238) <= OutputImg1_238_EXMPLR ;
   OutputImg1(237) <= OutputImg1_237_EXMPLR ;
   OutputImg1(236) <= OutputImg1_236_EXMPLR ;
   OutputImg1(235) <= OutputImg1_235_EXMPLR ;
   OutputImg1(234) <= OutputImg1_234_EXMPLR ;
   OutputImg1(233) <= OutputImg1_233_EXMPLR ;
   OutputImg1(232) <= OutputImg1_232_EXMPLR ;
   OutputImg1(231) <= OutputImg1_231_EXMPLR ;
   OutputImg1(230) <= OutputImg1_230_EXMPLR ;
   OutputImg1(229) <= OutputImg1_229_EXMPLR ;
   OutputImg1(228) <= OutputImg1_228_EXMPLR ;
   OutputImg1(227) <= OutputImg1_227_EXMPLR ;
   OutputImg1(226) <= OutputImg1_226_EXMPLR ;
   OutputImg1(225) <= OutputImg1_225_EXMPLR ;
   OutputImg1(224) <= OutputImg1_224_EXMPLR ;
   OutputImg1(223) <= OutputImg1_223_EXMPLR ;
   OutputImg1(222) <= OutputImg1_222_EXMPLR ;
   OutputImg1(221) <= OutputImg1_221_EXMPLR ;
   OutputImg1(220) <= OutputImg1_220_EXMPLR ;
   OutputImg1(219) <= OutputImg1_219_EXMPLR ;
   OutputImg1(218) <= OutputImg1_218_EXMPLR ;
   OutputImg1(217) <= OutputImg1_217_EXMPLR ;
   OutputImg1(216) <= OutputImg1_216_EXMPLR ;
   OutputImg1(215) <= OutputImg1_215_EXMPLR ;
   OutputImg1(214) <= OutputImg1_214_EXMPLR ;
   OutputImg1(213) <= OutputImg1_213_EXMPLR ;
   OutputImg1(212) <= OutputImg1_212_EXMPLR ;
   OutputImg1(211) <= OutputImg1_211_EXMPLR ;
   OutputImg1(210) <= OutputImg1_210_EXMPLR ;
   OutputImg1(209) <= OutputImg1_209_EXMPLR ;
   OutputImg1(208) <= OutputImg1_208_EXMPLR ;
   OutputImg1(207) <= OutputImg1_207_EXMPLR ;
   OutputImg1(206) <= OutputImg1_206_EXMPLR ;
   OutputImg1(205) <= OutputImg1_205_EXMPLR ;
   OutputImg1(204) <= OutputImg1_204_EXMPLR ;
   OutputImg1(203) <= OutputImg1_203_EXMPLR ;
   OutputImg1(202) <= OutputImg1_202_EXMPLR ;
   OutputImg1(201) <= OutputImg1_201_EXMPLR ;
   OutputImg1(200) <= OutputImg1_200_EXMPLR ;
   OutputImg1(199) <= OutputImg1_199_EXMPLR ;
   OutputImg1(198) <= OutputImg1_198_EXMPLR ;
   OutputImg1(197) <= OutputImg1_197_EXMPLR ;
   OutputImg1(196) <= OutputImg1_196_EXMPLR ;
   OutputImg1(195) <= OutputImg1_195_EXMPLR ;
   OutputImg1(194) <= OutputImg1_194_EXMPLR ;
   OutputImg1(193) <= OutputImg1_193_EXMPLR ;
   OutputImg1(192) <= OutputImg1_192_EXMPLR ;
   OutputImg1(191) <= OutputImg1_191_EXMPLR ;
   OutputImg1(190) <= OutputImg1_190_EXMPLR ;
   OutputImg1(189) <= OutputImg1_189_EXMPLR ;
   OutputImg1(188) <= OutputImg1_188_EXMPLR ;
   OutputImg1(187) <= OutputImg1_187_EXMPLR ;
   OutputImg1(186) <= OutputImg1_186_EXMPLR ;
   OutputImg1(185) <= OutputImg1_185_EXMPLR ;
   OutputImg1(184) <= OutputImg1_184_EXMPLR ;
   OutputImg1(183) <= OutputImg1_183_EXMPLR ;
   OutputImg1(182) <= OutputImg1_182_EXMPLR ;
   OutputImg1(181) <= OutputImg1_181_EXMPLR ;
   OutputImg1(180) <= OutputImg1_180_EXMPLR ;
   OutputImg1(179) <= OutputImg1_179_EXMPLR ;
   OutputImg1(178) <= OutputImg1_178_EXMPLR ;
   OutputImg1(177) <= OutputImg1_177_EXMPLR ;
   OutputImg1(176) <= OutputImg1_176_EXMPLR ;
   OutputImg1(175) <= OutputImg1_175_EXMPLR ;
   OutputImg1(174) <= OutputImg1_174_EXMPLR ;
   OutputImg1(173) <= OutputImg1_173_EXMPLR ;
   OutputImg1(172) <= OutputImg1_172_EXMPLR ;
   OutputImg1(171) <= OutputImg1_171_EXMPLR ;
   OutputImg1(170) <= OutputImg1_170_EXMPLR ;
   OutputImg1(169) <= OutputImg1_169_EXMPLR ;
   OutputImg1(168) <= OutputImg1_168_EXMPLR ;
   OutputImg1(167) <= OutputImg1_167_EXMPLR ;
   OutputImg1(166) <= OutputImg1_166_EXMPLR ;
   OutputImg1(165) <= OutputImg1_165_EXMPLR ;
   OutputImg1(164) <= OutputImg1_164_EXMPLR ;
   OutputImg1(163) <= OutputImg1_163_EXMPLR ;
   OutputImg1(162) <= OutputImg1_162_EXMPLR ;
   OutputImg1(161) <= OutputImg1_161_EXMPLR ;
   OutputImg1(160) <= OutputImg1_160_EXMPLR ;
   OutputImg1(159) <= OutputImg1_159_EXMPLR ;
   OutputImg1(158) <= OutputImg1_158_EXMPLR ;
   OutputImg1(157) <= OutputImg1_157_EXMPLR ;
   OutputImg1(156) <= OutputImg1_156_EXMPLR ;
   OutputImg1(155) <= OutputImg1_155_EXMPLR ;
   OutputImg1(154) <= OutputImg1_154_EXMPLR ;
   OutputImg1(153) <= OutputImg1_153_EXMPLR ;
   OutputImg1(152) <= OutputImg1_152_EXMPLR ;
   OutputImg1(151) <= OutputImg1_151_EXMPLR ;
   OutputImg1(150) <= OutputImg1_150_EXMPLR ;
   OutputImg1(149) <= OutputImg1_149_EXMPLR ;
   OutputImg1(148) <= OutputImg1_148_EXMPLR ;
   OutputImg1(147) <= OutputImg1_147_EXMPLR ;
   OutputImg1(146) <= OutputImg1_146_EXMPLR ;
   OutputImg1(145) <= OutputImg1_145_EXMPLR ;
   OutputImg1(144) <= OutputImg1_144_EXMPLR ;
   OutputImg1(143) <= OutputImg1_143_EXMPLR ;
   OutputImg1(142) <= OutputImg1_142_EXMPLR ;
   OutputImg1(141) <= OutputImg1_141_EXMPLR ;
   OutputImg1(140) <= OutputImg1_140_EXMPLR ;
   OutputImg1(139) <= OutputImg1_139_EXMPLR ;
   OutputImg1(138) <= OutputImg1_138_EXMPLR ;
   OutputImg1(137) <= OutputImg1_137_EXMPLR ;
   OutputImg1(136) <= OutputImg1_136_EXMPLR ;
   OutputImg1(135) <= OutputImg1_135_EXMPLR ;
   OutputImg1(134) <= OutputImg1_134_EXMPLR ;
   OutputImg1(133) <= OutputImg1_133_EXMPLR ;
   OutputImg1(132) <= OutputImg1_132_EXMPLR ;
   OutputImg1(131) <= OutputImg1_131_EXMPLR ;
   OutputImg1(130) <= OutputImg1_130_EXMPLR ;
   OutputImg1(129) <= OutputImg1_129_EXMPLR ;
   OutputImg1(128) <= OutputImg1_128_EXMPLR ;
   OutputImg1(127) <= OutputImg1_127_EXMPLR ;
   OutputImg1(126) <= OutputImg1_126_EXMPLR ;
   OutputImg1(125) <= OutputImg1_125_EXMPLR ;
   OutputImg1(124) <= OutputImg1_124_EXMPLR ;
   OutputImg1(123) <= OutputImg1_123_EXMPLR ;
   OutputImg1(122) <= OutputImg1_122_EXMPLR ;
   OutputImg1(121) <= OutputImg1_121_EXMPLR ;
   OutputImg1(120) <= OutputImg1_120_EXMPLR ;
   OutputImg1(119) <= OutputImg1_119_EXMPLR ;
   OutputImg1(118) <= OutputImg1_118_EXMPLR ;
   OutputImg1(117) <= OutputImg1_117_EXMPLR ;
   OutputImg1(116) <= OutputImg1_116_EXMPLR ;
   OutputImg1(115) <= OutputImg1_115_EXMPLR ;
   OutputImg1(114) <= OutputImg1_114_EXMPLR ;
   OutputImg1(113) <= OutputImg1_113_EXMPLR ;
   OutputImg1(112) <= OutputImg1_112_EXMPLR ;
   OutputImg1(111) <= OutputImg1_111_EXMPLR ;
   OutputImg1(110) <= OutputImg1_110_EXMPLR ;
   OutputImg1(109) <= OutputImg1_109_EXMPLR ;
   OutputImg1(108) <= OutputImg1_108_EXMPLR ;
   OutputImg1(107) <= OutputImg1_107_EXMPLR ;
   OutputImg1(106) <= OutputImg1_106_EXMPLR ;
   OutputImg1(105) <= OutputImg1_105_EXMPLR ;
   OutputImg1(104) <= OutputImg1_104_EXMPLR ;
   OutputImg1(103) <= OutputImg1_103_EXMPLR ;
   OutputImg1(102) <= OutputImg1_102_EXMPLR ;
   OutputImg1(101) <= OutputImg1_101_EXMPLR ;
   OutputImg1(100) <= OutputImg1_100_EXMPLR ;
   OutputImg1(99) <= OutputImg1_99_EXMPLR ;
   OutputImg1(98) <= OutputImg1_98_EXMPLR ;
   OutputImg1(97) <= OutputImg1_97_EXMPLR ;
   OutputImg1(96) <= OutputImg1_96_EXMPLR ;
   OutputImg1(95) <= OutputImg1_95_EXMPLR ;
   OutputImg1(94) <= OutputImg1_94_EXMPLR ;
   OutputImg1(93) <= OutputImg1_93_EXMPLR ;
   OutputImg1(92) <= OutputImg1_92_EXMPLR ;
   OutputImg1(91) <= OutputImg1_91_EXMPLR ;
   OutputImg1(90) <= OutputImg1_90_EXMPLR ;
   OutputImg1(89) <= OutputImg1_89_EXMPLR ;
   OutputImg1(88) <= OutputImg1_88_EXMPLR ;
   OutputImg1(87) <= OutputImg1_87_EXMPLR ;
   OutputImg1(86) <= OutputImg1_86_EXMPLR ;
   OutputImg1(85) <= OutputImg1_85_EXMPLR ;
   OutputImg1(84) <= OutputImg1_84_EXMPLR ;
   OutputImg1(83) <= OutputImg1_83_EXMPLR ;
   OutputImg1(82) <= OutputImg1_82_EXMPLR ;
   OutputImg1(81) <= OutputImg1_81_EXMPLR ;
   OutputImg1(80) <= OutputImg1_80_EXMPLR ;
   OutputImg1(79) <= OutputImg1_79_EXMPLR ;
   OutputImg1(78) <= OutputImg1_78_EXMPLR ;
   OutputImg1(77) <= OutputImg1_77_EXMPLR ;
   OutputImg1(76) <= OutputImg1_76_EXMPLR ;
   OutputImg1(75) <= OutputImg1_75_EXMPLR ;
   OutputImg1(74) <= OutputImg1_74_EXMPLR ;
   OutputImg1(73) <= OutputImg1_73_EXMPLR ;
   OutputImg1(72) <= OutputImg1_72_EXMPLR ;
   OutputImg1(71) <= OutputImg1_71_EXMPLR ;
   OutputImg1(70) <= OutputImg1_70_EXMPLR ;
   OutputImg1(69) <= OutputImg1_69_EXMPLR ;
   OutputImg1(68) <= OutputImg1_68_EXMPLR ;
   OutputImg1(67) <= OutputImg1_67_EXMPLR ;
   OutputImg1(66) <= OutputImg1_66_EXMPLR ;
   OutputImg1(65) <= OutputImg1_65_EXMPLR ;
   OutputImg1(64) <= OutputImg1_64_EXMPLR ;
   OutputImg1(63) <= OutputImg1_63_EXMPLR ;
   OutputImg1(62) <= OutputImg1_62_EXMPLR ;
   OutputImg1(61) <= OutputImg1_61_EXMPLR ;
   OutputImg1(60) <= OutputImg1_60_EXMPLR ;
   OutputImg1(59) <= OutputImg1_59_EXMPLR ;
   OutputImg1(58) <= OutputImg1_58_EXMPLR ;
   OutputImg1(57) <= OutputImg1_57_EXMPLR ;
   OutputImg1(56) <= OutputImg1_56_EXMPLR ;
   OutputImg1(55) <= OutputImg1_55_EXMPLR ;
   OutputImg1(54) <= OutputImg1_54_EXMPLR ;
   OutputImg1(53) <= OutputImg1_53_EXMPLR ;
   OutputImg1(52) <= OutputImg1_52_EXMPLR ;
   OutputImg1(51) <= OutputImg1_51_EXMPLR ;
   OutputImg1(50) <= OutputImg1_50_EXMPLR ;
   OutputImg1(49) <= OutputImg1_49_EXMPLR ;
   OutputImg1(48) <= OutputImg1_48_EXMPLR ;
   OutputImg1(47) <= OutputImg1_47_EXMPLR ;
   OutputImg1(46) <= OutputImg1_46_EXMPLR ;
   OutputImg1(45) <= OutputImg1_45_EXMPLR ;
   OutputImg1(44) <= OutputImg1_44_EXMPLR ;
   OutputImg1(43) <= OutputImg1_43_EXMPLR ;
   OutputImg1(42) <= OutputImg1_42_EXMPLR ;
   OutputImg1(41) <= OutputImg1_41_EXMPLR ;
   OutputImg1(40) <= OutputImg1_40_EXMPLR ;
   OutputImg1(39) <= OutputImg1_39_EXMPLR ;
   OutputImg1(38) <= OutputImg1_38_EXMPLR ;
   OutputImg1(37) <= OutputImg1_37_EXMPLR ;
   OutputImg1(36) <= OutputImg1_36_EXMPLR ;
   OutputImg1(35) <= OutputImg1_35_EXMPLR ;
   OutputImg1(34) <= OutputImg1_34_EXMPLR ;
   OutputImg1(33) <= OutputImg1_33_EXMPLR ;
   OutputImg1(32) <= OutputImg1_32_EXMPLR ;
   OutputImg1(31) <= OutputImg1_31_EXMPLR ;
   OutputImg1(30) <= OutputImg1_30_EXMPLR ;
   OutputImg1(29) <= OutputImg1_29_EXMPLR ;
   OutputImg1(28) <= OutputImg1_28_EXMPLR ;
   OutputImg1(27) <= OutputImg1_27_EXMPLR ;
   OutputImg1(26) <= OutputImg1_26_EXMPLR ;
   OutputImg1(25) <= OutputImg1_25_EXMPLR ;
   OutputImg1(24) <= OutputImg1_24_EXMPLR ;
   OutputImg1(23) <= OutputImg1_23_EXMPLR ;
   OutputImg1(22) <= OutputImg1_22_EXMPLR ;
   OutputImg1(21) <= OutputImg1_21_EXMPLR ;
   OutputImg1(20) <= OutputImg1_20_EXMPLR ;
   OutputImg1(19) <= OutputImg1_19_EXMPLR ;
   OutputImg1(18) <= OutputImg1_18_EXMPLR ;
   OutputImg1(17) <= OutputImg1_17_EXMPLR ;
   OutputImg1(16) <= OutputImg1_16_EXMPLR ;
   OutputImg1(15) <= OutputImg1_15_EXMPLR ;
   OutputImg1(14) <= OutputImg1_14_EXMPLR ;
   OutputImg1(13) <= OutputImg1_13_EXMPLR ;
   OutputImg1(12) <= OutputImg1_12_EXMPLR ;
   OutputImg1(11) <= OutputImg1_11_EXMPLR ;
   OutputImg1(10) <= OutputImg1_10_EXMPLR ;
   OutputImg1(9) <= OutputImg1_9_EXMPLR ;
   OutputImg1(8) <= OutputImg1_8_EXMPLR ;
   OutputImg1(7) <= OutputImg1_7_EXMPLR ;
   OutputImg1(6) <= OutputImg1_6_EXMPLR ;
   OutputImg1(5) <= OutputImg1_5_EXMPLR ;
   OutputImg1(4) <= OutputImg1_4_EXMPLR ;
   OutputImg1(3) <= OutputImg1_3_EXMPLR ;
   OutputImg1(2) <= OutputImg1_2_EXMPLR ;
   OutputImg1(1) <= OutputImg1_1_EXMPLR ;
   OutputImg1(0) <= OutputImg1_0_EXMPLR ;
   OutputImg2(447) <= OutputImg2_447_EXMPLR ;
   OutputImg2(446) <= OutputImg2_446_EXMPLR ;
   OutputImg2(445) <= OutputImg2_445_EXMPLR ;
   OutputImg2(444) <= OutputImg2_444_EXMPLR ;
   OutputImg2(443) <= OutputImg2_443_EXMPLR ;
   OutputImg2(442) <= OutputImg2_442_EXMPLR ;
   OutputImg2(441) <= OutputImg2_441_EXMPLR ;
   OutputImg2(440) <= OutputImg2_440_EXMPLR ;
   OutputImg2(439) <= OutputImg2_439_EXMPLR ;
   OutputImg2(438) <= OutputImg2_438_EXMPLR ;
   OutputImg2(437) <= OutputImg2_437_EXMPLR ;
   OutputImg2(436) <= OutputImg2_436_EXMPLR ;
   OutputImg2(435) <= OutputImg2_435_EXMPLR ;
   OutputImg2(434) <= OutputImg2_434_EXMPLR ;
   OutputImg2(433) <= OutputImg2_433_EXMPLR ;
   OutputImg2(432) <= OutputImg2_432_EXMPLR ;
   OutputImg2(431) <= OutputImg2_431_EXMPLR ;
   OutputImg2(430) <= OutputImg2_430_EXMPLR ;
   OutputImg2(429) <= OutputImg2_429_EXMPLR ;
   OutputImg2(428) <= OutputImg2_428_EXMPLR ;
   OutputImg2(427) <= OutputImg2_427_EXMPLR ;
   OutputImg2(426) <= OutputImg2_426_EXMPLR ;
   OutputImg2(425) <= OutputImg2_425_EXMPLR ;
   OutputImg2(424) <= OutputImg2_424_EXMPLR ;
   OutputImg2(423) <= OutputImg2_423_EXMPLR ;
   OutputImg2(422) <= OutputImg2_422_EXMPLR ;
   OutputImg2(421) <= OutputImg2_421_EXMPLR ;
   OutputImg2(420) <= OutputImg2_420_EXMPLR ;
   OutputImg2(419) <= OutputImg2_419_EXMPLR ;
   OutputImg2(418) <= OutputImg2_418_EXMPLR ;
   OutputImg2(417) <= OutputImg2_417_EXMPLR ;
   OutputImg2(416) <= OutputImg2_416_EXMPLR ;
   OutputImg2(415) <= OutputImg2_415_EXMPLR ;
   OutputImg2(414) <= OutputImg2_414_EXMPLR ;
   OutputImg2(413) <= OutputImg2_413_EXMPLR ;
   OutputImg2(412) <= OutputImg2_412_EXMPLR ;
   OutputImg2(411) <= OutputImg2_411_EXMPLR ;
   OutputImg2(410) <= OutputImg2_410_EXMPLR ;
   OutputImg2(409) <= OutputImg2_409_EXMPLR ;
   OutputImg2(408) <= OutputImg2_408_EXMPLR ;
   OutputImg2(407) <= OutputImg2_407_EXMPLR ;
   OutputImg2(406) <= OutputImg2_406_EXMPLR ;
   OutputImg2(405) <= OutputImg2_405_EXMPLR ;
   OutputImg2(404) <= OutputImg2_404_EXMPLR ;
   OutputImg2(403) <= OutputImg2_403_EXMPLR ;
   OutputImg2(402) <= OutputImg2_402_EXMPLR ;
   OutputImg2(401) <= OutputImg2_401_EXMPLR ;
   OutputImg2(400) <= OutputImg2_400_EXMPLR ;
   OutputImg2(399) <= OutputImg2_399_EXMPLR ;
   OutputImg2(398) <= OutputImg2_398_EXMPLR ;
   OutputImg2(397) <= OutputImg2_397_EXMPLR ;
   OutputImg2(396) <= OutputImg2_396_EXMPLR ;
   OutputImg2(395) <= OutputImg2_395_EXMPLR ;
   OutputImg2(394) <= OutputImg2_394_EXMPLR ;
   OutputImg2(393) <= OutputImg2_393_EXMPLR ;
   OutputImg2(392) <= OutputImg2_392_EXMPLR ;
   OutputImg2(391) <= OutputImg2_391_EXMPLR ;
   OutputImg2(390) <= OutputImg2_390_EXMPLR ;
   OutputImg2(389) <= OutputImg2_389_EXMPLR ;
   OutputImg2(388) <= OutputImg2_388_EXMPLR ;
   OutputImg2(387) <= OutputImg2_387_EXMPLR ;
   OutputImg2(386) <= OutputImg2_386_EXMPLR ;
   OutputImg2(385) <= OutputImg2_385_EXMPLR ;
   OutputImg2(384) <= OutputImg2_384_EXMPLR ;
   OutputImg2(383) <= OutputImg2_383_EXMPLR ;
   OutputImg2(382) <= OutputImg2_382_EXMPLR ;
   OutputImg2(381) <= OutputImg2_381_EXMPLR ;
   OutputImg2(380) <= OutputImg2_380_EXMPLR ;
   OutputImg2(379) <= OutputImg2_379_EXMPLR ;
   OutputImg2(378) <= OutputImg2_378_EXMPLR ;
   OutputImg2(377) <= OutputImg2_377_EXMPLR ;
   OutputImg2(376) <= OutputImg2_376_EXMPLR ;
   OutputImg2(375) <= OutputImg2_375_EXMPLR ;
   OutputImg2(374) <= OutputImg2_374_EXMPLR ;
   OutputImg2(373) <= OutputImg2_373_EXMPLR ;
   OutputImg2(372) <= OutputImg2_372_EXMPLR ;
   OutputImg2(371) <= OutputImg2_371_EXMPLR ;
   OutputImg2(370) <= OutputImg2_370_EXMPLR ;
   OutputImg2(369) <= OutputImg2_369_EXMPLR ;
   OutputImg2(368) <= OutputImg2_368_EXMPLR ;
   OutputImg2(367) <= OutputImg2_367_EXMPLR ;
   OutputImg2(366) <= OutputImg2_366_EXMPLR ;
   OutputImg2(365) <= OutputImg2_365_EXMPLR ;
   OutputImg2(364) <= OutputImg2_364_EXMPLR ;
   OutputImg2(363) <= OutputImg2_363_EXMPLR ;
   OutputImg2(362) <= OutputImg2_362_EXMPLR ;
   OutputImg2(361) <= OutputImg2_361_EXMPLR ;
   OutputImg2(360) <= OutputImg2_360_EXMPLR ;
   OutputImg2(359) <= OutputImg2_359_EXMPLR ;
   OutputImg2(358) <= OutputImg2_358_EXMPLR ;
   OutputImg2(357) <= OutputImg2_357_EXMPLR ;
   OutputImg2(356) <= OutputImg2_356_EXMPLR ;
   OutputImg2(355) <= OutputImg2_355_EXMPLR ;
   OutputImg2(354) <= OutputImg2_354_EXMPLR ;
   OutputImg2(353) <= OutputImg2_353_EXMPLR ;
   OutputImg2(352) <= OutputImg2_352_EXMPLR ;
   OutputImg2(351) <= OutputImg2_351_EXMPLR ;
   OutputImg2(350) <= OutputImg2_350_EXMPLR ;
   OutputImg2(349) <= OutputImg2_349_EXMPLR ;
   OutputImg2(348) <= OutputImg2_348_EXMPLR ;
   OutputImg2(347) <= OutputImg2_347_EXMPLR ;
   OutputImg2(346) <= OutputImg2_346_EXMPLR ;
   OutputImg2(345) <= OutputImg2_345_EXMPLR ;
   OutputImg2(344) <= OutputImg2_344_EXMPLR ;
   OutputImg2(343) <= OutputImg2_343_EXMPLR ;
   OutputImg2(342) <= OutputImg2_342_EXMPLR ;
   OutputImg2(341) <= OutputImg2_341_EXMPLR ;
   OutputImg2(340) <= OutputImg2_340_EXMPLR ;
   OutputImg2(339) <= OutputImg2_339_EXMPLR ;
   OutputImg2(338) <= OutputImg2_338_EXMPLR ;
   OutputImg2(337) <= OutputImg2_337_EXMPLR ;
   OutputImg2(336) <= OutputImg2_336_EXMPLR ;
   OutputImg2(335) <= OutputImg2_335_EXMPLR ;
   OutputImg2(334) <= OutputImg2_334_EXMPLR ;
   OutputImg2(333) <= OutputImg2_333_EXMPLR ;
   OutputImg2(332) <= OutputImg2_332_EXMPLR ;
   OutputImg2(331) <= OutputImg2_331_EXMPLR ;
   OutputImg2(330) <= OutputImg2_330_EXMPLR ;
   OutputImg2(329) <= OutputImg2_329_EXMPLR ;
   OutputImg2(328) <= OutputImg2_328_EXMPLR ;
   OutputImg2(327) <= OutputImg2_327_EXMPLR ;
   OutputImg2(326) <= OutputImg2_326_EXMPLR ;
   OutputImg2(325) <= OutputImg2_325_EXMPLR ;
   OutputImg2(324) <= OutputImg2_324_EXMPLR ;
   OutputImg2(323) <= OutputImg2_323_EXMPLR ;
   OutputImg2(322) <= OutputImg2_322_EXMPLR ;
   OutputImg2(321) <= OutputImg2_321_EXMPLR ;
   OutputImg2(320) <= OutputImg2_320_EXMPLR ;
   OutputImg2(319) <= OutputImg2_319_EXMPLR ;
   OutputImg2(318) <= OutputImg2_318_EXMPLR ;
   OutputImg2(317) <= OutputImg2_317_EXMPLR ;
   OutputImg2(316) <= OutputImg2_316_EXMPLR ;
   OutputImg2(315) <= OutputImg2_315_EXMPLR ;
   OutputImg2(314) <= OutputImg2_314_EXMPLR ;
   OutputImg2(313) <= OutputImg2_313_EXMPLR ;
   OutputImg2(312) <= OutputImg2_312_EXMPLR ;
   OutputImg2(311) <= OutputImg2_311_EXMPLR ;
   OutputImg2(310) <= OutputImg2_310_EXMPLR ;
   OutputImg2(309) <= OutputImg2_309_EXMPLR ;
   OutputImg2(308) <= OutputImg2_308_EXMPLR ;
   OutputImg2(307) <= OutputImg2_307_EXMPLR ;
   OutputImg2(306) <= OutputImg2_306_EXMPLR ;
   OutputImg2(305) <= OutputImg2_305_EXMPLR ;
   OutputImg2(304) <= OutputImg2_304_EXMPLR ;
   OutputImg2(303) <= OutputImg2_303_EXMPLR ;
   OutputImg2(302) <= OutputImg2_302_EXMPLR ;
   OutputImg2(301) <= OutputImg2_301_EXMPLR ;
   OutputImg2(300) <= OutputImg2_300_EXMPLR ;
   OutputImg2(299) <= OutputImg2_299_EXMPLR ;
   OutputImg2(298) <= OutputImg2_298_EXMPLR ;
   OutputImg2(297) <= OutputImg2_297_EXMPLR ;
   OutputImg2(296) <= OutputImg2_296_EXMPLR ;
   OutputImg2(295) <= OutputImg2_295_EXMPLR ;
   OutputImg2(294) <= OutputImg2_294_EXMPLR ;
   OutputImg2(293) <= OutputImg2_293_EXMPLR ;
   OutputImg2(292) <= OutputImg2_292_EXMPLR ;
   OutputImg2(291) <= OutputImg2_291_EXMPLR ;
   OutputImg2(290) <= OutputImg2_290_EXMPLR ;
   OutputImg2(289) <= OutputImg2_289_EXMPLR ;
   OutputImg2(288) <= OutputImg2_288_EXMPLR ;
   OutputImg2(287) <= OutputImg2_287_EXMPLR ;
   OutputImg2(286) <= OutputImg2_286_EXMPLR ;
   OutputImg2(285) <= OutputImg2_285_EXMPLR ;
   OutputImg2(284) <= OutputImg2_284_EXMPLR ;
   OutputImg2(283) <= OutputImg2_283_EXMPLR ;
   OutputImg2(282) <= OutputImg2_282_EXMPLR ;
   OutputImg2(281) <= OutputImg2_281_EXMPLR ;
   OutputImg2(280) <= OutputImg2_280_EXMPLR ;
   OutputImg2(279) <= OutputImg2_279_EXMPLR ;
   OutputImg2(278) <= OutputImg2_278_EXMPLR ;
   OutputImg2(277) <= OutputImg2_277_EXMPLR ;
   OutputImg2(276) <= OutputImg2_276_EXMPLR ;
   OutputImg2(275) <= OutputImg2_275_EXMPLR ;
   OutputImg2(274) <= OutputImg2_274_EXMPLR ;
   OutputImg2(273) <= OutputImg2_273_EXMPLR ;
   OutputImg2(272) <= OutputImg2_272_EXMPLR ;
   OutputImg2(271) <= OutputImg2_271_EXMPLR ;
   OutputImg2(270) <= OutputImg2_270_EXMPLR ;
   OutputImg2(269) <= OutputImg2_269_EXMPLR ;
   OutputImg2(268) <= OutputImg2_268_EXMPLR ;
   OutputImg2(267) <= OutputImg2_267_EXMPLR ;
   OutputImg2(266) <= OutputImg2_266_EXMPLR ;
   OutputImg2(265) <= OutputImg2_265_EXMPLR ;
   OutputImg2(264) <= OutputImg2_264_EXMPLR ;
   OutputImg2(263) <= OutputImg2_263_EXMPLR ;
   OutputImg2(262) <= OutputImg2_262_EXMPLR ;
   OutputImg2(261) <= OutputImg2_261_EXMPLR ;
   OutputImg2(260) <= OutputImg2_260_EXMPLR ;
   OutputImg2(259) <= OutputImg2_259_EXMPLR ;
   OutputImg2(258) <= OutputImg2_258_EXMPLR ;
   OutputImg2(257) <= OutputImg2_257_EXMPLR ;
   OutputImg2(256) <= OutputImg2_256_EXMPLR ;
   OutputImg2(255) <= OutputImg2_255_EXMPLR ;
   OutputImg2(254) <= OutputImg2_254_EXMPLR ;
   OutputImg2(253) <= OutputImg2_253_EXMPLR ;
   OutputImg2(252) <= OutputImg2_252_EXMPLR ;
   OutputImg2(251) <= OutputImg2_251_EXMPLR ;
   OutputImg2(250) <= OutputImg2_250_EXMPLR ;
   OutputImg2(249) <= OutputImg2_249_EXMPLR ;
   OutputImg2(248) <= OutputImg2_248_EXMPLR ;
   OutputImg2(247) <= OutputImg2_247_EXMPLR ;
   OutputImg2(246) <= OutputImg2_246_EXMPLR ;
   OutputImg2(245) <= OutputImg2_245_EXMPLR ;
   OutputImg2(244) <= OutputImg2_244_EXMPLR ;
   OutputImg2(243) <= OutputImg2_243_EXMPLR ;
   OutputImg2(242) <= OutputImg2_242_EXMPLR ;
   OutputImg2(241) <= OutputImg2_241_EXMPLR ;
   OutputImg2(240) <= OutputImg2_240_EXMPLR ;
   OutputImg2(239) <= OutputImg2_239_EXMPLR ;
   OutputImg2(238) <= OutputImg2_238_EXMPLR ;
   OutputImg2(237) <= OutputImg2_237_EXMPLR ;
   OutputImg2(236) <= OutputImg2_236_EXMPLR ;
   OutputImg2(235) <= OutputImg2_235_EXMPLR ;
   OutputImg2(234) <= OutputImg2_234_EXMPLR ;
   OutputImg2(233) <= OutputImg2_233_EXMPLR ;
   OutputImg2(232) <= OutputImg2_232_EXMPLR ;
   OutputImg2(231) <= OutputImg2_231_EXMPLR ;
   OutputImg2(230) <= OutputImg2_230_EXMPLR ;
   OutputImg2(229) <= OutputImg2_229_EXMPLR ;
   OutputImg2(228) <= OutputImg2_228_EXMPLR ;
   OutputImg2(227) <= OutputImg2_227_EXMPLR ;
   OutputImg2(226) <= OutputImg2_226_EXMPLR ;
   OutputImg2(225) <= OutputImg2_225_EXMPLR ;
   OutputImg2(224) <= OutputImg2_224_EXMPLR ;
   OutputImg2(223) <= OutputImg2_223_EXMPLR ;
   OutputImg2(222) <= OutputImg2_222_EXMPLR ;
   OutputImg2(221) <= OutputImg2_221_EXMPLR ;
   OutputImg2(220) <= OutputImg2_220_EXMPLR ;
   OutputImg2(219) <= OutputImg2_219_EXMPLR ;
   OutputImg2(218) <= OutputImg2_218_EXMPLR ;
   OutputImg2(217) <= OutputImg2_217_EXMPLR ;
   OutputImg2(216) <= OutputImg2_216_EXMPLR ;
   OutputImg2(215) <= OutputImg2_215_EXMPLR ;
   OutputImg2(214) <= OutputImg2_214_EXMPLR ;
   OutputImg2(213) <= OutputImg2_213_EXMPLR ;
   OutputImg2(212) <= OutputImg2_212_EXMPLR ;
   OutputImg2(211) <= OutputImg2_211_EXMPLR ;
   OutputImg2(210) <= OutputImg2_210_EXMPLR ;
   OutputImg2(209) <= OutputImg2_209_EXMPLR ;
   OutputImg2(208) <= OutputImg2_208_EXMPLR ;
   OutputImg2(207) <= OutputImg2_207_EXMPLR ;
   OutputImg2(206) <= OutputImg2_206_EXMPLR ;
   OutputImg2(205) <= OutputImg2_205_EXMPLR ;
   OutputImg2(204) <= OutputImg2_204_EXMPLR ;
   OutputImg2(203) <= OutputImg2_203_EXMPLR ;
   OutputImg2(202) <= OutputImg2_202_EXMPLR ;
   OutputImg2(201) <= OutputImg2_201_EXMPLR ;
   OutputImg2(200) <= OutputImg2_200_EXMPLR ;
   OutputImg2(199) <= OutputImg2_199_EXMPLR ;
   OutputImg2(198) <= OutputImg2_198_EXMPLR ;
   OutputImg2(197) <= OutputImg2_197_EXMPLR ;
   OutputImg2(196) <= OutputImg2_196_EXMPLR ;
   OutputImg2(195) <= OutputImg2_195_EXMPLR ;
   OutputImg2(194) <= OutputImg2_194_EXMPLR ;
   OutputImg2(193) <= OutputImg2_193_EXMPLR ;
   OutputImg2(192) <= OutputImg2_192_EXMPLR ;
   OutputImg2(191) <= OutputImg2_191_EXMPLR ;
   OutputImg2(190) <= OutputImg2_190_EXMPLR ;
   OutputImg2(189) <= OutputImg2_189_EXMPLR ;
   OutputImg2(188) <= OutputImg2_188_EXMPLR ;
   OutputImg2(187) <= OutputImg2_187_EXMPLR ;
   OutputImg2(186) <= OutputImg2_186_EXMPLR ;
   OutputImg2(185) <= OutputImg2_185_EXMPLR ;
   OutputImg2(184) <= OutputImg2_184_EXMPLR ;
   OutputImg2(183) <= OutputImg2_183_EXMPLR ;
   OutputImg2(182) <= OutputImg2_182_EXMPLR ;
   OutputImg2(181) <= OutputImg2_181_EXMPLR ;
   OutputImg2(180) <= OutputImg2_180_EXMPLR ;
   OutputImg2(179) <= OutputImg2_179_EXMPLR ;
   OutputImg2(178) <= OutputImg2_178_EXMPLR ;
   OutputImg2(177) <= OutputImg2_177_EXMPLR ;
   OutputImg2(176) <= OutputImg2_176_EXMPLR ;
   OutputImg2(175) <= OutputImg2_175_EXMPLR ;
   OutputImg2(174) <= OutputImg2_174_EXMPLR ;
   OutputImg2(173) <= OutputImg2_173_EXMPLR ;
   OutputImg2(172) <= OutputImg2_172_EXMPLR ;
   OutputImg2(171) <= OutputImg2_171_EXMPLR ;
   OutputImg2(170) <= OutputImg2_170_EXMPLR ;
   OutputImg2(169) <= OutputImg2_169_EXMPLR ;
   OutputImg2(168) <= OutputImg2_168_EXMPLR ;
   OutputImg2(167) <= OutputImg2_167_EXMPLR ;
   OutputImg2(166) <= OutputImg2_166_EXMPLR ;
   OutputImg2(165) <= OutputImg2_165_EXMPLR ;
   OutputImg2(164) <= OutputImg2_164_EXMPLR ;
   OutputImg2(163) <= OutputImg2_163_EXMPLR ;
   OutputImg2(162) <= OutputImg2_162_EXMPLR ;
   OutputImg2(161) <= OutputImg2_161_EXMPLR ;
   OutputImg2(160) <= OutputImg2_160_EXMPLR ;
   OutputImg2(159) <= OutputImg2_159_EXMPLR ;
   OutputImg2(158) <= OutputImg2_158_EXMPLR ;
   OutputImg2(157) <= OutputImg2_157_EXMPLR ;
   OutputImg2(156) <= OutputImg2_156_EXMPLR ;
   OutputImg2(155) <= OutputImg2_155_EXMPLR ;
   OutputImg2(154) <= OutputImg2_154_EXMPLR ;
   OutputImg2(153) <= OutputImg2_153_EXMPLR ;
   OutputImg2(152) <= OutputImg2_152_EXMPLR ;
   OutputImg2(151) <= OutputImg2_151_EXMPLR ;
   OutputImg2(150) <= OutputImg2_150_EXMPLR ;
   OutputImg2(149) <= OutputImg2_149_EXMPLR ;
   OutputImg2(148) <= OutputImg2_148_EXMPLR ;
   OutputImg2(147) <= OutputImg2_147_EXMPLR ;
   OutputImg2(146) <= OutputImg2_146_EXMPLR ;
   OutputImg2(145) <= OutputImg2_145_EXMPLR ;
   OutputImg2(144) <= OutputImg2_144_EXMPLR ;
   OutputImg2(143) <= OutputImg2_143_EXMPLR ;
   OutputImg2(142) <= OutputImg2_142_EXMPLR ;
   OutputImg2(141) <= OutputImg2_141_EXMPLR ;
   OutputImg2(140) <= OutputImg2_140_EXMPLR ;
   OutputImg2(139) <= OutputImg2_139_EXMPLR ;
   OutputImg2(138) <= OutputImg2_138_EXMPLR ;
   OutputImg2(137) <= OutputImg2_137_EXMPLR ;
   OutputImg2(136) <= OutputImg2_136_EXMPLR ;
   OutputImg2(135) <= OutputImg2_135_EXMPLR ;
   OutputImg2(134) <= OutputImg2_134_EXMPLR ;
   OutputImg2(133) <= OutputImg2_133_EXMPLR ;
   OutputImg2(132) <= OutputImg2_132_EXMPLR ;
   OutputImg2(131) <= OutputImg2_131_EXMPLR ;
   OutputImg2(130) <= OutputImg2_130_EXMPLR ;
   OutputImg2(129) <= OutputImg2_129_EXMPLR ;
   OutputImg2(128) <= OutputImg2_128_EXMPLR ;
   OutputImg2(127) <= OutputImg2_127_EXMPLR ;
   OutputImg2(126) <= OutputImg2_126_EXMPLR ;
   OutputImg2(125) <= OutputImg2_125_EXMPLR ;
   OutputImg2(124) <= OutputImg2_124_EXMPLR ;
   OutputImg2(123) <= OutputImg2_123_EXMPLR ;
   OutputImg2(122) <= OutputImg2_122_EXMPLR ;
   OutputImg2(121) <= OutputImg2_121_EXMPLR ;
   OutputImg2(120) <= OutputImg2_120_EXMPLR ;
   OutputImg2(119) <= OutputImg2_119_EXMPLR ;
   OutputImg2(118) <= OutputImg2_118_EXMPLR ;
   OutputImg2(117) <= OutputImg2_117_EXMPLR ;
   OutputImg2(116) <= OutputImg2_116_EXMPLR ;
   OutputImg2(115) <= OutputImg2_115_EXMPLR ;
   OutputImg2(114) <= OutputImg2_114_EXMPLR ;
   OutputImg2(113) <= OutputImg2_113_EXMPLR ;
   OutputImg2(112) <= OutputImg2_112_EXMPLR ;
   OutputImg2(111) <= OutputImg2_111_EXMPLR ;
   OutputImg2(110) <= OutputImg2_110_EXMPLR ;
   OutputImg2(109) <= OutputImg2_109_EXMPLR ;
   OutputImg2(108) <= OutputImg2_108_EXMPLR ;
   OutputImg2(107) <= OutputImg2_107_EXMPLR ;
   OutputImg2(106) <= OutputImg2_106_EXMPLR ;
   OutputImg2(105) <= OutputImg2_105_EXMPLR ;
   OutputImg2(104) <= OutputImg2_104_EXMPLR ;
   OutputImg2(103) <= OutputImg2_103_EXMPLR ;
   OutputImg2(102) <= OutputImg2_102_EXMPLR ;
   OutputImg2(101) <= OutputImg2_101_EXMPLR ;
   OutputImg2(100) <= OutputImg2_100_EXMPLR ;
   OutputImg2(99) <= OutputImg2_99_EXMPLR ;
   OutputImg2(98) <= OutputImg2_98_EXMPLR ;
   OutputImg2(97) <= OutputImg2_97_EXMPLR ;
   OutputImg2(96) <= OutputImg2_96_EXMPLR ;
   OutputImg2(95) <= OutputImg2_95_EXMPLR ;
   OutputImg2(94) <= OutputImg2_94_EXMPLR ;
   OutputImg2(93) <= OutputImg2_93_EXMPLR ;
   OutputImg2(92) <= OutputImg2_92_EXMPLR ;
   OutputImg2(91) <= OutputImg2_91_EXMPLR ;
   OutputImg2(90) <= OutputImg2_90_EXMPLR ;
   OutputImg2(89) <= OutputImg2_89_EXMPLR ;
   OutputImg2(88) <= OutputImg2_88_EXMPLR ;
   OutputImg2(87) <= OutputImg2_87_EXMPLR ;
   OutputImg2(86) <= OutputImg2_86_EXMPLR ;
   OutputImg2(85) <= OutputImg2_85_EXMPLR ;
   OutputImg2(84) <= OutputImg2_84_EXMPLR ;
   OutputImg2(83) <= OutputImg2_83_EXMPLR ;
   OutputImg2(82) <= OutputImg2_82_EXMPLR ;
   OutputImg2(81) <= OutputImg2_81_EXMPLR ;
   OutputImg2(80) <= OutputImg2_80_EXMPLR ;
   OutputImg2(79) <= OutputImg2_79_EXMPLR ;
   OutputImg2(78) <= OutputImg2_78_EXMPLR ;
   OutputImg2(77) <= OutputImg2_77_EXMPLR ;
   OutputImg2(76) <= OutputImg2_76_EXMPLR ;
   OutputImg2(75) <= OutputImg2_75_EXMPLR ;
   OutputImg2(74) <= OutputImg2_74_EXMPLR ;
   OutputImg2(73) <= OutputImg2_73_EXMPLR ;
   OutputImg2(72) <= OutputImg2_72_EXMPLR ;
   OutputImg2(71) <= OutputImg2_71_EXMPLR ;
   OutputImg2(70) <= OutputImg2_70_EXMPLR ;
   OutputImg2(69) <= OutputImg2_69_EXMPLR ;
   OutputImg2(68) <= OutputImg2_68_EXMPLR ;
   OutputImg2(67) <= OutputImg2_67_EXMPLR ;
   OutputImg2(66) <= OutputImg2_66_EXMPLR ;
   OutputImg2(65) <= OutputImg2_65_EXMPLR ;
   OutputImg2(64) <= OutputImg2_64_EXMPLR ;
   OutputImg2(63) <= OutputImg2_63_EXMPLR ;
   OutputImg2(62) <= OutputImg2_62_EXMPLR ;
   OutputImg2(61) <= OutputImg2_61_EXMPLR ;
   OutputImg2(60) <= OutputImg2_60_EXMPLR ;
   OutputImg2(59) <= OutputImg2_59_EXMPLR ;
   OutputImg2(58) <= OutputImg2_58_EXMPLR ;
   OutputImg2(57) <= OutputImg2_57_EXMPLR ;
   OutputImg2(56) <= OutputImg2_56_EXMPLR ;
   OutputImg2(55) <= OutputImg2_55_EXMPLR ;
   OutputImg2(54) <= OutputImg2_54_EXMPLR ;
   OutputImg2(53) <= OutputImg2_53_EXMPLR ;
   OutputImg2(52) <= OutputImg2_52_EXMPLR ;
   OutputImg2(51) <= OutputImg2_51_EXMPLR ;
   OutputImg2(50) <= OutputImg2_50_EXMPLR ;
   OutputImg2(49) <= OutputImg2_49_EXMPLR ;
   OutputImg2(48) <= OutputImg2_48_EXMPLR ;
   OutputImg2(47) <= OutputImg2_47_EXMPLR ;
   OutputImg2(46) <= OutputImg2_46_EXMPLR ;
   OutputImg2(45) <= OutputImg2_45_EXMPLR ;
   OutputImg2(44) <= OutputImg2_44_EXMPLR ;
   OutputImg2(43) <= OutputImg2_43_EXMPLR ;
   OutputImg2(42) <= OutputImg2_42_EXMPLR ;
   OutputImg2(41) <= OutputImg2_41_EXMPLR ;
   OutputImg2(40) <= OutputImg2_40_EXMPLR ;
   OutputImg2(39) <= OutputImg2_39_EXMPLR ;
   OutputImg2(38) <= OutputImg2_38_EXMPLR ;
   OutputImg2(37) <= OutputImg2_37_EXMPLR ;
   OutputImg2(36) <= OutputImg2_36_EXMPLR ;
   OutputImg2(35) <= OutputImg2_35_EXMPLR ;
   OutputImg2(34) <= OutputImg2_34_EXMPLR ;
   OutputImg2(33) <= OutputImg2_33_EXMPLR ;
   OutputImg2(32) <= OutputImg2_32_EXMPLR ;
   OutputImg2(31) <= OutputImg2_31_EXMPLR ;
   OutputImg2(30) <= OutputImg2_30_EXMPLR ;
   OutputImg2(29) <= OutputImg2_29_EXMPLR ;
   OutputImg2(28) <= OutputImg2_28_EXMPLR ;
   OutputImg2(27) <= OutputImg2_27_EXMPLR ;
   OutputImg2(26) <= OutputImg2_26_EXMPLR ;
   OutputImg2(25) <= OutputImg2_25_EXMPLR ;
   OutputImg2(24) <= OutputImg2_24_EXMPLR ;
   OutputImg2(23) <= OutputImg2_23_EXMPLR ;
   OutputImg2(22) <= OutputImg2_22_EXMPLR ;
   OutputImg2(21) <= OutputImg2_21_EXMPLR ;
   OutputImg2(20) <= OutputImg2_20_EXMPLR ;
   OutputImg2(19) <= OutputImg2_19_EXMPLR ;
   OutputImg2(18) <= OutputImg2_18_EXMPLR ;
   OutputImg2(17) <= OutputImg2_17_EXMPLR ;
   OutputImg2(16) <= OutputImg2_16_EXMPLR ;
   OutputImg2(15) <= OutputImg2_15_EXMPLR ;
   OutputImg2(14) <= OutputImg2_14_EXMPLR ;
   OutputImg2(13) <= OutputImg2_13_EXMPLR ;
   OutputImg2(12) <= OutputImg2_12_EXMPLR ;
   OutputImg2(11) <= OutputImg2_11_EXMPLR ;
   OutputImg2(10) <= OutputImg2_10_EXMPLR ;
   OutputImg2(9) <= OutputImg2_9_EXMPLR ;
   OutputImg2(8) <= OutputImg2_8_EXMPLR ;
   OutputImg2(7) <= OutputImg2_7_EXMPLR ;
   OutputImg2(6) <= OutputImg2_6_EXMPLR ;
   OutputImg2(5) <= OutputImg2_5_EXMPLR ;
   OutputImg2(4) <= OutputImg2_4_EXMPLR ;
   OutputImg2(3) <= OutputImg2_3_EXMPLR ;
   OutputImg2(2) <= OutputImg2_2_EXMPLR ;
   OutputImg2(1) <= OutputImg2_1_EXMPLR ;
   OutputImg2(0) <= OutputImg2_0_EXMPLR ;
   OutputImg3(447) <= OutputImg3_447_EXMPLR ;
   OutputImg3(446) <= OutputImg3_446_EXMPLR ;
   OutputImg3(445) <= OutputImg3_445_EXMPLR ;
   OutputImg3(444) <= OutputImg3_444_EXMPLR ;
   OutputImg3(443) <= OutputImg3_443_EXMPLR ;
   OutputImg3(442) <= OutputImg3_442_EXMPLR ;
   OutputImg3(441) <= OutputImg3_441_EXMPLR ;
   OutputImg3(440) <= OutputImg3_440_EXMPLR ;
   OutputImg3(439) <= OutputImg3_439_EXMPLR ;
   OutputImg3(438) <= OutputImg3_438_EXMPLR ;
   OutputImg3(437) <= OutputImg3_437_EXMPLR ;
   OutputImg3(436) <= OutputImg3_436_EXMPLR ;
   OutputImg3(435) <= OutputImg3_435_EXMPLR ;
   OutputImg3(434) <= OutputImg3_434_EXMPLR ;
   OutputImg3(433) <= OutputImg3_433_EXMPLR ;
   OutputImg3(432) <= OutputImg3_432_EXMPLR ;
   OutputImg3(431) <= OutputImg3_431_EXMPLR ;
   OutputImg3(430) <= OutputImg3_430_EXMPLR ;
   OutputImg3(429) <= OutputImg3_429_EXMPLR ;
   OutputImg3(428) <= OutputImg3_428_EXMPLR ;
   OutputImg3(427) <= OutputImg3_427_EXMPLR ;
   OutputImg3(426) <= OutputImg3_426_EXMPLR ;
   OutputImg3(425) <= OutputImg3_425_EXMPLR ;
   OutputImg3(424) <= OutputImg3_424_EXMPLR ;
   OutputImg3(423) <= OutputImg3_423_EXMPLR ;
   OutputImg3(422) <= OutputImg3_422_EXMPLR ;
   OutputImg3(421) <= OutputImg3_421_EXMPLR ;
   OutputImg3(420) <= OutputImg3_420_EXMPLR ;
   OutputImg3(419) <= OutputImg3_419_EXMPLR ;
   OutputImg3(418) <= OutputImg3_418_EXMPLR ;
   OutputImg3(417) <= OutputImg3_417_EXMPLR ;
   OutputImg3(416) <= OutputImg3_416_EXMPLR ;
   OutputImg3(415) <= OutputImg3_415_EXMPLR ;
   OutputImg3(414) <= OutputImg3_414_EXMPLR ;
   OutputImg3(413) <= OutputImg3_413_EXMPLR ;
   OutputImg3(412) <= OutputImg3_412_EXMPLR ;
   OutputImg3(411) <= OutputImg3_411_EXMPLR ;
   OutputImg3(410) <= OutputImg3_410_EXMPLR ;
   OutputImg3(409) <= OutputImg3_409_EXMPLR ;
   OutputImg3(408) <= OutputImg3_408_EXMPLR ;
   OutputImg3(407) <= OutputImg3_407_EXMPLR ;
   OutputImg3(406) <= OutputImg3_406_EXMPLR ;
   OutputImg3(405) <= OutputImg3_405_EXMPLR ;
   OutputImg3(404) <= OutputImg3_404_EXMPLR ;
   OutputImg3(403) <= OutputImg3_403_EXMPLR ;
   OutputImg3(402) <= OutputImg3_402_EXMPLR ;
   OutputImg3(401) <= OutputImg3_401_EXMPLR ;
   OutputImg3(400) <= OutputImg3_400_EXMPLR ;
   OutputImg3(399) <= OutputImg3_399_EXMPLR ;
   OutputImg3(398) <= OutputImg3_398_EXMPLR ;
   OutputImg3(397) <= OutputImg3_397_EXMPLR ;
   OutputImg3(396) <= OutputImg3_396_EXMPLR ;
   OutputImg3(395) <= OutputImg3_395_EXMPLR ;
   OutputImg3(394) <= OutputImg3_394_EXMPLR ;
   OutputImg3(393) <= OutputImg3_393_EXMPLR ;
   OutputImg3(392) <= OutputImg3_392_EXMPLR ;
   OutputImg3(391) <= OutputImg3_391_EXMPLR ;
   OutputImg3(390) <= OutputImg3_390_EXMPLR ;
   OutputImg3(389) <= OutputImg3_389_EXMPLR ;
   OutputImg3(388) <= OutputImg3_388_EXMPLR ;
   OutputImg3(387) <= OutputImg3_387_EXMPLR ;
   OutputImg3(386) <= OutputImg3_386_EXMPLR ;
   OutputImg3(385) <= OutputImg3_385_EXMPLR ;
   OutputImg3(384) <= OutputImg3_384_EXMPLR ;
   OutputImg3(383) <= OutputImg3_383_EXMPLR ;
   OutputImg3(382) <= OutputImg3_382_EXMPLR ;
   OutputImg3(381) <= OutputImg3_381_EXMPLR ;
   OutputImg3(380) <= OutputImg3_380_EXMPLR ;
   OutputImg3(379) <= OutputImg3_379_EXMPLR ;
   OutputImg3(378) <= OutputImg3_378_EXMPLR ;
   OutputImg3(377) <= OutputImg3_377_EXMPLR ;
   OutputImg3(376) <= OutputImg3_376_EXMPLR ;
   OutputImg3(375) <= OutputImg3_375_EXMPLR ;
   OutputImg3(374) <= OutputImg3_374_EXMPLR ;
   OutputImg3(373) <= OutputImg3_373_EXMPLR ;
   OutputImg3(372) <= OutputImg3_372_EXMPLR ;
   OutputImg3(371) <= OutputImg3_371_EXMPLR ;
   OutputImg3(370) <= OutputImg3_370_EXMPLR ;
   OutputImg3(369) <= OutputImg3_369_EXMPLR ;
   OutputImg3(368) <= OutputImg3_368_EXMPLR ;
   OutputImg3(367) <= OutputImg3_367_EXMPLR ;
   OutputImg3(366) <= OutputImg3_366_EXMPLR ;
   OutputImg3(365) <= OutputImg3_365_EXMPLR ;
   OutputImg3(364) <= OutputImg3_364_EXMPLR ;
   OutputImg3(363) <= OutputImg3_363_EXMPLR ;
   OutputImg3(362) <= OutputImg3_362_EXMPLR ;
   OutputImg3(361) <= OutputImg3_361_EXMPLR ;
   OutputImg3(360) <= OutputImg3_360_EXMPLR ;
   OutputImg3(359) <= OutputImg3_359_EXMPLR ;
   OutputImg3(358) <= OutputImg3_358_EXMPLR ;
   OutputImg3(357) <= OutputImg3_357_EXMPLR ;
   OutputImg3(356) <= OutputImg3_356_EXMPLR ;
   OutputImg3(355) <= OutputImg3_355_EXMPLR ;
   OutputImg3(354) <= OutputImg3_354_EXMPLR ;
   OutputImg3(353) <= OutputImg3_353_EXMPLR ;
   OutputImg3(352) <= OutputImg3_352_EXMPLR ;
   OutputImg3(351) <= OutputImg3_351_EXMPLR ;
   OutputImg3(350) <= OutputImg3_350_EXMPLR ;
   OutputImg3(349) <= OutputImg3_349_EXMPLR ;
   OutputImg3(348) <= OutputImg3_348_EXMPLR ;
   OutputImg3(347) <= OutputImg3_347_EXMPLR ;
   OutputImg3(346) <= OutputImg3_346_EXMPLR ;
   OutputImg3(345) <= OutputImg3_345_EXMPLR ;
   OutputImg3(344) <= OutputImg3_344_EXMPLR ;
   OutputImg3(343) <= OutputImg3_343_EXMPLR ;
   OutputImg3(342) <= OutputImg3_342_EXMPLR ;
   OutputImg3(341) <= OutputImg3_341_EXMPLR ;
   OutputImg3(340) <= OutputImg3_340_EXMPLR ;
   OutputImg3(339) <= OutputImg3_339_EXMPLR ;
   OutputImg3(338) <= OutputImg3_338_EXMPLR ;
   OutputImg3(337) <= OutputImg3_337_EXMPLR ;
   OutputImg3(336) <= OutputImg3_336_EXMPLR ;
   OutputImg3(335) <= OutputImg3_335_EXMPLR ;
   OutputImg3(334) <= OutputImg3_334_EXMPLR ;
   OutputImg3(333) <= OutputImg3_333_EXMPLR ;
   OutputImg3(332) <= OutputImg3_332_EXMPLR ;
   OutputImg3(331) <= OutputImg3_331_EXMPLR ;
   OutputImg3(330) <= OutputImg3_330_EXMPLR ;
   OutputImg3(329) <= OutputImg3_329_EXMPLR ;
   OutputImg3(328) <= OutputImg3_328_EXMPLR ;
   OutputImg3(327) <= OutputImg3_327_EXMPLR ;
   OutputImg3(326) <= OutputImg3_326_EXMPLR ;
   OutputImg3(325) <= OutputImg3_325_EXMPLR ;
   OutputImg3(324) <= OutputImg3_324_EXMPLR ;
   OutputImg3(323) <= OutputImg3_323_EXMPLR ;
   OutputImg3(322) <= OutputImg3_322_EXMPLR ;
   OutputImg3(321) <= OutputImg3_321_EXMPLR ;
   OutputImg3(320) <= OutputImg3_320_EXMPLR ;
   OutputImg3(319) <= OutputImg3_319_EXMPLR ;
   OutputImg3(318) <= OutputImg3_318_EXMPLR ;
   OutputImg3(317) <= OutputImg3_317_EXMPLR ;
   OutputImg3(316) <= OutputImg3_316_EXMPLR ;
   OutputImg3(315) <= OutputImg3_315_EXMPLR ;
   OutputImg3(314) <= OutputImg3_314_EXMPLR ;
   OutputImg3(313) <= OutputImg3_313_EXMPLR ;
   OutputImg3(312) <= OutputImg3_312_EXMPLR ;
   OutputImg3(311) <= OutputImg3_311_EXMPLR ;
   OutputImg3(310) <= OutputImg3_310_EXMPLR ;
   OutputImg3(309) <= OutputImg3_309_EXMPLR ;
   OutputImg3(308) <= OutputImg3_308_EXMPLR ;
   OutputImg3(307) <= OutputImg3_307_EXMPLR ;
   OutputImg3(306) <= OutputImg3_306_EXMPLR ;
   OutputImg3(305) <= OutputImg3_305_EXMPLR ;
   OutputImg3(304) <= OutputImg3_304_EXMPLR ;
   OutputImg3(303) <= OutputImg3_303_EXMPLR ;
   OutputImg3(302) <= OutputImg3_302_EXMPLR ;
   OutputImg3(301) <= OutputImg3_301_EXMPLR ;
   OutputImg3(300) <= OutputImg3_300_EXMPLR ;
   OutputImg3(299) <= OutputImg3_299_EXMPLR ;
   OutputImg3(298) <= OutputImg3_298_EXMPLR ;
   OutputImg3(297) <= OutputImg3_297_EXMPLR ;
   OutputImg3(296) <= OutputImg3_296_EXMPLR ;
   OutputImg3(295) <= OutputImg3_295_EXMPLR ;
   OutputImg3(294) <= OutputImg3_294_EXMPLR ;
   OutputImg3(293) <= OutputImg3_293_EXMPLR ;
   OutputImg3(292) <= OutputImg3_292_EXMPLR ;
   OutputImg3(291) <= OutputImg3_291_EXMPLR ;
   OutputImg3(290) <= OutputImg3_290_EXMPLR ;
   OutputImg3(289) <= OutputImg3_289_EXMPLR ;
   OutputImg3(288) <= OutputImg3_288_EXMPLR ;
   OutputImg3(287) <= OutputImg3_287_EXMPLR ;
   OutputImg3(286) <= OutputImg3_286_EXMPLR ;
   OutputImg3(285) <= OutputImg3_285_EXMPLR ;
   OutputImg3(284) <= OutputImg3_284_EXMPLR ;
   OutputImg3(283) <= OutputImg3_283_EXMPLR ;
   OutputImg3(282) <= OutputImg3_282_EXMPLR ;
   OutputImg3(281) <= OutputImg3_281_EXMPLR ;
   OutputImg3(280) <= OutputImg3_280_EXMPLR ;
   OutputImg3(279) <= OutputImg3_279_EXMPLR ;
   OutputImg3(278) <= OutputImg3_278_EXMPLR ;
   OutputImg3(277) <= OutputImg3_277_EXMPLR ;
   OutputImg3(276) <= OutputImg3_276_EXMPLR ;
   OutputImg3(275) <= OutputImg3_275_EXMPLR ;
   OutputImg3(274) <= OutputImg3_274_EXMPLR ;
   OutputImg3(273) <= OutputImg3_273_EXMPLR ;
   OutputImg3(272) <= OutputImg3_272_EXMPLR ;
   OutputImg3(271) <= OutputImg3_271_EXMPLR ;
   OutputImg3(270) <= OutputImg3_270_EXMPLR ;
   OutputImg3(269) <= OutputImg3_269_EXMPLR ;
   OutputImg3(268) <= OutputImg3_268_EXMPLR ;
   OutputImg3(267) <= OutputImg3_267_EXMPLR ;
   OutputImg3(266) <= OutputImg3_266_EXMPLR ;
   OutputImg3(265) <= OutputImg3_265_EXMPLR ;
   OutputImg3(264) <= OutputImg3_264_EXMPLR ;
   OutputImg3(263) <= OutputImg3_263_EXMPLR ;
   OutputImg3(262) <= OutputImg3_262_EXMPLR ;
   OutputImg3(261) <= OutputImg3_261_EXMPLR ;
   OutputImg3(260) <= OutputImg3_260_EXMPLR ;
   OutputImg3(259) <= OutputImg3_259_EXMPLR ;
   OutputImg3(258) <= OutputImg3_258_EXMPLR ;
   OutputImg3(257) <= OutputImg3_257_EXMPLR ;
   OutputImg3(256) <= OutputImg3_256_EXMPLR ;
   OutputImg3(255) <= OutputImg3_255_EXMPLR ;
   OutputImg3(254) <= OutputImg3_254_EXMPLR ;
   OutputImg3(253) <= OutputImg3_253_EXMPLR ;
   OutputImg3(252) <= OutputImg3_252_EXMPLR ;
   OutputImg3(251) <= OutputImg3_251_EXMPLR ;
   OutputImg3(250) <= OutputImg3_250_EXMPLR ;
   OutputImg3(249) <= OutputImg3_249_EXMPLR ;
   OutputImg3(248) <= OutputImg3_248_EXMPLR ;
   OutputImg3(247) <= OutputImg3_247_EXMPLR ;
   OutputImg3(246) <= OutputImg3_246_EXMPLR ;
   OutputImg3(245) <= OutputImg3_245_EXMPLR ;
   OutputImg3(244) <= OutputImg3_244_EXMPLR ;
   OutputImg3(243) <= OutputImg3_243_EXMPLR ;
   OutputImg3(242) <= OutputImg3_242_EXMPLR ;
   OutputImg3(241) <= OutputImg3_241_EXMPLR ;
   OutputImg3(240) <= OutputImg3_240_EXMPLR ;
   OutputImg3(239) <= OutputImg3_239_EXMPLR ;
   OutputImg3(238) <= OutputImg3_238_EXMPLR ;
   OutputImg3(237) <= OutputImg3_237_EXMPLR ;
   OutputImg3(236) <= OutputImg3_236_EXMPLR ;
   OutputImg3(235) <= OutputImg3_235_EXMPLR ;
   OutputImg3(234) <= OutputImg3_234_EXMPLR ;
   OutputImg3(233) <= OutputImg3_233_EXMPLR ;
   OutputImg3(232) <= OutputImg3_232_EXMPLR ;
   OutputImg3(231) <= OutputImg3_231_EXMPLR ;
   OutputImg3(230) <= OutputImg3_230_EXMPLR ;
   OutputImg3(229) <= OutputImg3_229_EXMPLR ;
   OutputImg3(228) <= OutputImg3_228_EXMPLR ;
   OutputImg3(227) <= OutputImg3_227_EXMPLR ;
   OutputImg3(226) <= OutputImg3_226_EXMPLR ;
   OutputImg3(225) <= OutputImg3_225_EXMPLR ;
   OutputImg3(224) <= OutputImg3_224_EXMPLR ;
   OutputImg3(223) <= OutputImg3_223_EXMPLR ;
   OutputImg3(222) <= OutputImg3_222_EXMPLR ;
   OutputImg3(221) <= OutputImg3_221_EXMPLR ;
   OutputImg3(220) <= OutputImg3_220_EXMPLR ;
   OutputImg3(219) <= OutputImg3_219_EXMPLR ;
   OutputImg3(218) <= OutputImg3_218_EXMPLR ;
   OutputImg3(217) <= OutputImg3_217_EXMPLR ;
   OutputImg3(216) <= OutputImg3_216_EXMPLR ;
   OutputImg3(215) <= OutputImg3_215_EXMPLR ;
   OutputImg3(214) <= OutputImg3_214_EXMPLR ;
   OutputImg3(213) <= OutputImg3_213_EXMPLR ;
   OutputImg3(212) <= OutputImg3_212_EXMPLR ;
   OutputImg3(211) <= OutputImg3_211_EXMPLR ;
   OutputImg3(210) <= OutputImg3_210_EXMPLR ;
   OutputImg3(209) <= OutputImg3_209_EXMPLR ;
   OutputImg3(208) <= OutputImg3_208_EXMPLR ;
   OutputImg3(207) <= OutputImg3_207_EXMPLR ;
   OutputImg3(206) <= OutputImg3_206_EXMPLR ;
   OutputImg3(205) <= OutputImg3_205_EXMPLR ;
   OutputImg3(204) <= OutputImg3_204_EXMPLR ;
   OutputImg3(203) <= OutputImg3_203_EXMPLR ;
   OutputImg3(202) <= OutputImg3_202_EXMPLR ;
   OutputImg3(201) <= OutputImg3_201_EXMPLR ;
   OutputImg3(200) <= OutputImg3_200_EXMPLR ;
   OutputImg3(199) <= OutputImg3_199_EXMPLR ;
   OutputImg3(198) <= OutputImg3_198_EXMPLR ;
   OutputImg3(197) <= OutputImg3_197_EXMPLR ;
   OutputImg3(196) <= OutputImg3_196_EXMPLR ;
   OutputImg3(195) <= OutputImg3_195_EXMPLR ;
   OutputImg3(194) <= OutputImg3_194_EXMPLR ;
   OutputImg3(193) <= OutputImg3_193_EXMPLR ;
   OutputImg3(192) <= OutputImg3_192_EXMPLR ;
   OutputImg3(191) <= OutputImg3_191_EXMPLR ;
   OutputImg3(190) <= OutputImg3_190_EXMPLR ;
   OutputImg3(189) <= OutputImg3_189_EXMPLR ;
   OutputImg3(188) <= OutputImg3_188_EXMPLR ;
   OutputImg3(187) <= OutputImg3_187_EXMPLR ;
   OutputImg3(186) <= OutputImg3_186_EXMPLR ;
   OutputImg3(185) <= OutputImg3_185_EXMPLR ;
   OutputImg3(184) <= OutputImg3_184_EXMPLR ;
   OutputImg3(183) <= OutputImg3_183_EXMPLR ;
   OutputImg3(182) <= OutputImg3_182_EXMPLR ;
   OutputImg3(181) <= OutputImg3_181_EXMPLR ;
   OutputImg3(180) <= OutputImg3_180_EXMPLR ;
   OutputImg3(179) <= OutputImg3_179_EXMPLR ;
   OutputImg3(178) <= OutputImg3_178_EXMPLR ;
   OutputImg3(177) <= OutputImg3_177_EXMPLR ;
   OutputImg3(176) <= OutputImg3_176_EXMPLR ;
   OutputImg3(175) <= OutputImg3_175_EXMPLR ;
   OutputImg3(174) <= OutputImg3_174_EXMPLR ;
   OutputImg3(173) <= OutputImg3_173_EXMPLR ;
   OutputImg3(172) <= OutputImg3_172_EXMPLR ;
   OutputImg3(171) <= OutputImg3_171_EXMPLR ;
   OutputImg3(170) <= OutputImg3_170_EXMPLR ;
   OutputImg3(169) <= OutputImg3_169_EXMPLR ;
   OutputImg3(168) <= OutputImg3_168_EXMPLR ;
   OutputImg3(167) <= OutputImg3_167_EXMPLR ;
   OutputImg3(166) <= OutputImg3_166_EXMPLR ;
   OutputImg3(165) <= OutputImg3_165_EXMPLR ;
   OutputImg3(164) <= OutputImg3_164_EXMPLR ;
   OutputImg3(163) <= OutputImg3_163_EXMPLR ;
   OutputImg3(162) <= OutputImg3_162_EXMPLR ;
   OutputImg3(161) <= OutputImg3_161_EXMPLR ;
   OutputImg3(160) <= OutputImg3_160_EXMPLR ;
   OutputImg3(159) <= OutputImg3_159_EXMPLR ;
   OutputImg3(158) <= OutputImg3_158_EXMPLR ;
   OutputImg3(157) <= OutputImg3_157_EXMPLR ;
   OutputImg3(156) <= OutputImg3_156_EXMPLR ;
   OutputImg3(155) <= OutputImg3_155_EXMPLR ;
   OutputImg3(154) <= OutputImg3_154_EXMPLR ;
   OutputImg3(153) <= OutputImg3_153_EXMPLR ;
   OutputImg3(152) <= OutputImg3_152_EXMPLR ;
   OutputImg3(151) <= OutputImg3_151_EXMPLR ;
   OutputImg3(150) <= OutputImg3_150_EXMPLR ;
   OutputImg3(149) <= OutputImg3_149_EXMPLR ;
   OutputImg3(148) <= OutputImg3_148_EXMPLR ;
   OutputImg3(147) <= OutputImg3_147_EXMPLR ;
   OutputImg3(146) <= OutputImg3_146_EXMPLR ;
   OutputImg3(145) <= OutputImg3_145_EXMPLR ;
   OutputImg3(144) <= OutputImg3_144_EXMPLR ;
   OutputImg3(143) <= OutputImg3_143_EXMPLR ;
   OutputImg3(142) <= OutputImg3_142_EXMPLR ;
   OutputImg3(141) <= OutputImg3_141_EXMPLR ;
   OutputImg3(140) <= OutputImg3_140_EXMPLR ;
   OutputImg3(139) <= OutputImg3_139_EXMPLR ;
   OutputImg3(138) <= OutputImg3_138_EXMPLR ;
   OutputImg3(137) <= OutputImg3_137_EXMPLR ;
   OutputImg3(136) <= OutputImg3_136_EXMPLR ;
   OutputImg3(135) <= OutputImg3_135_EXMPLR ;
   OutputImg3(134) <= OutputImg3_134_EXMPLR ;
   OutputImg3(133) <= OutputImg3_133_EXMPLR ;
   OutputImg3(132) <= OutputImg3_132_EXMPLR ;
   OutputImg3(131) <= OutputImg3_131_EXMPLR ;
   OutputImg3(130) <= OutputImg3_130_EXMPLR ;
   OutputImg3(129) <= OutputImg3_129_EXMPLR ;
   OutputImg3(128) <= OutputImg3_128_EXMPLR ;
   OutputImg3(127) <= OutputImg3_127_EXMPLR ;
   OutputImg3(126) <= OutputImg3_126_EXMPLR ;
   OutputImg3(125) <= OutputImg3_125_EXMPLR ;
   OutputImg3(124) <= OutputImg3_124_EXMPLR ;
   OutputImg3(123) <= OutputImg3_123_EXMPLR ;
   OutputImg3(122) <= OutputImg3_122_EXMPLR ;
   OutputImg3(121) <= OutputImg3_121_EXMPLR ;
   OutputImg3(120) <= OutputImg3_120_EXMPLR ;
   OutputImg3(119) <= OutputImg3_119_EXMPLR ;
   OutputImg3(118) <= OutputImg3_118_EXMPLR ;
   OutputImg3(117) <= OutputImg3_117_EXMPLR ;
   OutputImg3(116) <= OutputImg3_116_EXMPLR ;
   OutputImg3(115) <= OutputImg3_115_EXMPLR ;
   OutputImg3(114) <= OutputImg3_114_EXMPLR ;
   OutputImg3(113) <= OutputImg3_113_EXMPLR ;
   OutputImg3(112) <= OutputImg3_112_EXMPLR ;
   OutputImg3(111) <= OutputImg3_111_EXMPLR ;
   OutputImg3(110) <= OutputImg3_110_EXMPLR ;
   OutputImg3(109) <= OutputImg3_109_EXMPLR ;
   OutputImg3(108) <= OutputImg3_108_EXMPLR ;
   OutputImg3(107) <= OutputImg3_107_EXMPLR ;
   OutputImg3(106) <= OutputImg3_106_EXMPLR ;
   OutputImg3(105) <= OutputImg3_105_EXMPLR ;
   OutputImg3(104) <= OutputImg3_104_EXMPLR ;
   OutputImg3(103) <= OutputImg3_103_EXMPLR ;
   OutputImg3(102) <= OutputImg3_102_EXMPLR ;
   OutputImg3(101) <= OutputImg3_101_EXMPLR ;
   OutputImg3(100) <= OutputImg3_100_EXMPLR ;
   OutputImg3(99) <= OutputImg3_99_EXMPLR ;
   OutputImg3(98) <= OutputImg3_98_EXMPLR ;
   OutputImg3(97) <= OutputImg3_97_EXMPLR ;
   OutputImg3(96) <= OutputImg3_96_EXMPLR ;
   OutputImg3(95) <= OutputImg3_95_EXMPLR ;
   OutputImg3(94) <= OutputImg3_94_EXMPLR ;
   OutputImg3(93) <= OutputImg3_93_EXMPLR ;
   OutputImg3(92) <= OutputImg3_92_EXMPLR ;
   OutputImg3(91) <= OutputImg3_91_EXMPLR ;
   OutputImg3(90) <= OutputImg3_90_EXMPLR ;
   OutputImg3(89) <= OutputImg3_89_EXMPLR ;
   OutputImg3(88) <= OutputImg3_88_EXMPLR ;
   OutputImg3(87) <= OutputImg3_87_EXMPLR ;
   OutputImg3(86) <= OutputImg3_86_EXMPLR ;
   OutputImg3(85) <= OutputImg3_85_EXMPLR ;
   OutputImg3(84) <= OutputImg3_84_EXMPLR ;
   OutputImg3(83) <= OutputImg3_83_EXMPLR ;
   OutputImg3(82) <= OutputImg3_82_EXMPLR ;
   OutputImg3(81) <= OutputImg3_81_EXMPLR ;
   OutputImg3(80) <= OutputImg3_80_EXMPLR ;
   OutputImg3(79) <= OutputImg3_79_EXMPLR ;
   OutputImg3(78) <= OutputImg3_78_EXMPLR ;
   OutputImg3(77) <= OutputImg3_77_EXMPLR ;
   OutputImg3(76) <= OutputImg3_76_EXMPLR ;
   OutputImg3(75) <= OutputImg3_75_EXMPLR ;
   OutputImg3(74) <= OutputImg3_74_EXMPLR ;
   OutputImg3(73) <= OutputImg3_73_EXMPLR ;
   OutputImg3(72) <= OutputImg3_72_EXMPLR ;
   OutputImg3(71) <= OutputImg3_71_EXMPLR ;
   OutputImg3(70) <= OutputImg3_70_EXMPLR ;
   OutputImg3(69) <= OutputImg3_69_EXMPLR ;
   OutputImg3(68) <= OutputImg3_68_EXMPLR ;
   OutputImg3(67) <= OutputImg3_67_EXMPLR ;
   OutputImg3(66) <= OutputImg3_66_EXMPLR ;
   OutputImg3(65) <= OutputImg3_65_EXMPLR ;
   OutputImg3(64) <= OutputImg3_64_EXMPLR ;
   OutputImg3(63) <= OutputImg3_63_EXMPLR ;
   OutputImg3(62) <= OutputImg3_62_EXMPLR ;
   OutputImg3(61) <= OutputImg3_61_EXMPLR ;
   OutputImg3(60) <= OutputImg3_60_EXMPLR ;
   OutputImg3(59) <= OutputImg3_59_EXMPLR ;
   OutputImg3(58) <= OutputImg3_58_EXMPLR ;
   OutputImg3(57) <= OutputImg3_57_EXMPLR ;
   OutputImg3(56) <= OutputImg3_56_EXMPLR ;
   OutputImg3(55) <= OutputImg3_55_EXMPLR ;
   OutputImg3(54) <= OutputImg3_54_EXMPLR ;
   OutputImg3(53) <= OutputImg3_53_EXMPLR ;
   OutputImg3(52) <= OutputImg3_52_EXMPLR ;
   OutputImg3(51) <= OutputImg3_51_EXMPLR ;
   OutputImg3(50) <= OutputImg3_50_EXMPLR ;
   OutputImg3(49) <= OutputImg3_49_EXMPLR ;
   OutputImg3(48) <= OutputImg3_48_EXMPLR ;
   OutputImg3(47) <= OutputImg3_47_EXMPLR ;
   OutputImg3(46) <= OutputImg3_46_EXMPLR ;
   OutputImg3(45) <= OutputImg3_45_EXMPLR ;
   OutputImg3(44) <= OutputImg3_44_EXMPLR ;
   OutputImg3(43) <= OutputImg3_43_EXMPLR ;
   OutputImg3(42) <= OutputImg3_42_EXMPLR ;
   OutputImg3(41) <= OutputImg3_41_EXMPLR ;
   OutputImg3(40) <= OutputImg3_40_EXMPLR ;
   OutputImg3(39) <= OutputImg3_39_EXMPLR ;
   OutputImg3(38) <= OutputImg3_38_EXMPLR ;
   OutputImg3(37) <= OutputImg3_37_EXMPLR ;
   OutputImg3(36) <= OutputImg3_36_EXMPLR ;
   OutputImg3(35) <= OutputImg3_35_EXMPLR ;
   OutputImg3(34) <= OutputImg3_34_EXMPLR ;
   OutputImg3(33) <= OutputImg3_33_EXMPLR ;
   OutputImg3(32) <= OutputImg3_32_EXMPLR ;
   OutputImg3(31) <= OutputImg3_31_EXMPLR ;
   OutputImg3(30) <= OutputImg3_30_EXMPLR ;
   OutputImg3(29) <= OutputImg3_29_EXMPLR ;
   OutputImg3(28) <= OutputImg3_28_EXMPLR ;
   OutputImg3(27) <= OutputImg3_27_EXMPLR ;
   OutputImg3(26) <= OutputImg3_26_EXMPLR ;
   OutputImg3(25) <= OutputImg3_25_EXMPLR ;
   OutputImg3(24) <= OutputImg3_24_EXMPLR ;
   OutputImg3(23) <= OutputImg3_23_EXMPLR ;
   OutputImg3(22) <= OutputImg3_22_EXMPLR ;
   OutputImg3(21) <= OutputImg3_21_EXMPLR ;
   OutputImg3(20) <= OutputImg3_20_EXMPLR ;
   OutputImg3(19) <= OutputImg3_19_EXMPLR ;
   OutputImg3(18) <= OutputImg3_18_EXMPLR ;
   OutputImg3(17) <= OutputImg3_17_EXMPLR ;
   OutputImg3(16) <= OutputImg3_16_EXMPLR ;
   OutputImg3(15) <= OutputImg3_15_EXMPLR ;
   OutputImg3(14) <= OutputImg3_14_EXMPLR ;
   OutputImg3(13) <= OutputImg3_13_EXMPLR ;
   OutputImg3(12) <= OutputImg3_12_EXMPLR ;
   OutputImg3(11) <= OutputImg3_11_EXMPLR ;
   OutputImg3(10) <= OutputImg3_10_EXMPLR ;
   OutputImg3(9) <= OutputImg3_9_EXMPLR ;
   OutputImg3(8) <= OutputImg3_8_EXMPLR ;
   OutputImg3(7) <= OutputImg3_7_EXMPLR ;
   OutputImg3(6) <= OutputImg3_6_EXMPLR ;
   OutputImg3(5) <= OutputImg3_5_EXMPLR ;
   OutputImg3(4) <= OutputImg3_4_EXMPLR ;
   OutputImg3(3) <= OutputImg3_3_EXMPLR ;
   OutputImg3(2) <= OutputImg3_2_EXMPLR ;
   OutputImg3(1) <= OutputImg3_1_EXMPLR ;
   OutputImg3(0) <= OutputImg3_0_EXMPLR ;
   OutputImg4(447) <= OutputImg4_447_EXMPLR ;
   OutputImg4(446) <= OutputImg4_446_EXMPLR ;
   OutputImg4(445) <= OutputImg4_445_EXMPLR ;
   OutputImg4(444) <= OutputImg4_444_EXMPLR ;
   OutputImg4(443) <= OutputImg4_443_EXMPLR ;
   OutputImg4(442) <= OutputImg4_442_EXMPLR ;
   OutputImg4(441) <= OutputImg4_441_EXMPLR ;
   OutputImg4(440) <= OutputImg4_440_EXMPLR ;
   OutputImg4(439) <= OutputImg4_439_EXMPLR ;
   OutputImg4(438) <= OutputImg4_438_EXMPLR ;
   OutputImg4(437) <= OutputImg4_437_EXMPLR ;
   OutputImg4(436) <= OutputImg4_436_EXMPLR ;
   OutputImg4(435) <= OutputImg4_435_EXMPLR ;
   OutputImg4(434) <= OutputImg4_434_EXMPLR ;
   OutputImg4(433) <= OutputImg4_433_EXMPLR ;
   OutputImg4(432) <= OutputImg4_432_EXMPLR ;
   OutputImg4(431) <= OutputImg4_431_EXMPLR ;
   OutputImg4(430) <= OutputImg4_430_EXMPLR ;
   OutputImg4(429) <= OutputImg4_429_EXMPLR ;
   OutputImg4(428) <= OutputImg4_428_EXMPLR ;
   OutputImg4(427) <= OutputImg4_427_EXMPLR ;
   OutputImg4(426) <= OutputImg4_426_EXMPLR ;
   OutputImg4(425) <= OutputImg4_425_EXMPLR ;
   OutputImg4(424) <= OutputImg4_424_EXMPLR ;
   OutputImg4(423) <= OutputImg4_423_EXMPLR ;
   OutputImg4(422) <= OutputImg4_422_EXMPLR ;
   OutputImg4(421) <= OutputImg4_421_EXMPLR ;
   OutputImg4(420) <= OutputImg4_420_EXMPLR ;
   OutputImg4(419) <= OutputImg4_419_EXMPLR ;
   OutputImg4(418) <= OutputImg4_418_EXMPLR ;
   OutputImg4(417) <= OutputImg4_417_EXMPLR ;
   OutputImg4(416) <= OutputImg4_416_EXMPLR ;
   OutputImg4(415) <= OutputImg4_415_EXMPLR ;
   OutputImg4(414) <= OutputImg4_414_EXMPLR ;
   OutputImg4(413) <= OutputImg4_413_EXMPLR ;
   OutputImg4(412) <= OutputImg4_412_EXMPLR ;
   OutputImg4(411) <= OutputImg4_411_EXMPLR ;
   OutputImg4(410) <= OutputImg4_410_EXMPLR ;
   OutputImg4(409) <= OutputImg4_409_EXMPLR ;
   OutputImg4(408) <= OutputImg4_408_EXMPLR ;
   OutputImg4(407) <= OutputImg4_407_EXMPLR ;
   OutputImg4(406) <= OutputImg4_406_EXMPLR ;
   OutputImg4(405) <= OutputImg4_405_EXMPLR ;
   OutputImg4(404) <= OutputImg4_404_EXMPLR ;
   OutputImg4(403) <= OutputImg4_403_EXMPLR ;
   OutputImg4(402) <= OutputImg4_402_EXMPLR ;
   OutputImg4(401) <= OutputImg4_401_EXMPLR ;
   OutputImg4(400) <= OutputImg4_400_EXMPLR ;
   OutputImg4(399) <= OutputImg4_399_EXMPLR ;
   OutputImg4(398) <= OutputImg4_398_EXMPLR ;
   OutputImg4(397) <= OutputImg4_397_EXMPLR ;
   OutputImg4(396) <= OutputImg4_396_EXMPLR ;
   OutputImg4(395) <= OutputImg4_395_EXMPLR ;
   OutputImg4(394) <= OutputImg4_394_EXMPLR ;
   OutputImg4(393) <= OutputImg4_393_EXMPLR ;
   OutputImg4(392) <= OutputImg4_392_EXMPLR ;
   OutputImg4(391) <= OutputImg4_391_EXMPLR ;
   OutputImg4(390) <= OutputImg4_390_EXMPLR ;
   OutputImg4(389) <= OutputImg4_389_EXMPLR ;
   OutputImg4(388) <= OutputImg4_388_EXMPLR ;
   OutputImg4(387) <= OutputImg4_387_EXMPLR ;
   OutputImg4(386) <= OutputImg4_386_EXMPLR ;
   OutputImg4(385) <= OutputImg4_385_EXMPLR ;
   OutputImg4(384) <= OutputImg4_384_EXMPLR ;
   OutputImg4(383) <= OutputImg4_383_EXMPLR ;
   OutputImg4(382) <= OutputImg4_382_EXMPLR ;
   OutputImg4(381) <= OutputImg4_381_EXMPLR ;
   OutputImg4(380) <= OutputImg4_380_EXMPLR ;
   OutputImg4(379) <= OutputImg4_379_EXMPLR ;
   OutputImg4(378) <= OutputImg4_378_EXMPLR ;
   OutputImg4(377) <= OutputImg4_377_EXMPLR ;
   OutputImg4(376) <= OutputImg4_376_EXMPLR ;
   OutputImg4(375) <= OutputImg4_375_EXMPLR ;
   OutputImg4(374) <= OutputImg4_374_EXMPLR ;
   OutputImg4(373) <= OutputImg4_373_EXMPLR ;
   OutputImg4(372) <= OutputImg4_372_EXMPLR ;
   OutputImg4(371) <= OutputImg4_371_EXMPLR ;
   OutputImg4(370) <= OutputImg4_370_EXMPLR ;
   OutputImg4(369) <= OutputImg4_369_EXMPLR ;
   OutputImg4(368) <= OutputImg4_368_EXMPLR ;
   OutputImg4(367) <= OutputImg4_367_EXMPLR ;
   OutputImg4(366) <= OutputImg4_366_EXMPLR ;
   OutputImg4(365) <= OutputImg4_365_EXMPLR ;
   OutputImg4(364) <= OutputImg4_364_EXMPLR ;
   OutputImg4(363) <= OutputImg4_363_EXMPLR ;
   OutputImg4(362) <= OutputImg4_362_EXMPLR ;
   OutputImg4(361) <= OutputImg4_361_EXMPLR ;
   OutputImg4(360) <= OutputImg4_360_EXMPLR ;
   OutputImg4(359) <= OutputImg4_359_EXMPLR ;
   OutputImg4(358) <= OutputImg4_358_EXMPLR ;
   OutputImg4(357) <= OutputImg4_357_EXMPLR ;
   OutputImg4(356) <= OutputImg4_356_EXMPLR ;
   OutputImg4(355) <= OutputImg4_355_EXMPLR ;
   OutputImg4(354) <= OutputImg4_354_EXMPLR ;
   OutputImg4(353) <= OutputImg4_353_EXMPLR ;
   OutputImg4(352) <= OutputImg4_352_EXMPLR ;
   OutputImg4(351) <= OutputImg4_351_EXMPLR ;
   OutputImg4(350) <= OutputImg4_350_EXMPLR ;
   OutputImg4(349) <= OutputImg4_349_EXMPLR ;
   OutputImg4(348) <= OutputImg4_348_EXMPLR ;
   OutputImg4(347) <= OutputImg4_347_EXMPLR ;
   OutputImg4(346) <= OutputImg4_346_EXMPLR ;
   OutputImg4(345) <= OutputImg4_345_EXMPLR ;
   OutputImg4(344) <= OutputImg4_344_EXMPLR ;
   OutputImg4(343) <= OutputImg4_343_EXMPLR ;
   OutputImg4(342) <= OutputImg4_342_EXMPLR ;
   OutputImg4(341) <= OutputImg4_341_EXMPLR ;
   OutputImg4(340) <= OutputImg4_340_EXMPLR ;
   OutputImg4(339) <= OutputImg4_339_EXMPLR ;
   OutputImg4(338) <= OutputImg4_338_EXMPLR ;
   OutputImg4(337) <= OutputImg4_337_EXMPLR ;
   OutputImg4(336) <= OutputImg4_336_EXMPLR ;
   OutputImg4(335) <= OutputImg4_335_EXMPLR ;
   OutputImg4(334) <= OutputImg4_334_EXMPLR ;
   OutputImg4(333) <= OutputImg4_333_EXMPLR ;
   OutputImg4(332) <= OutputImg4_332_EXMPLR ;
   OutputImg4(331) <= OutputImg4_331_EXMPLR ;
   OutputImg4(330) <= OutputImg4_330_EXMPLR ;
   OutputImg4(329) <= OutputImg4_329_EXMPLR ;
   OutputImg4(328) <= OutputImg4_328_EXMPLR ;
   OutputImg4(327) <= OutputImg4_327_EXMPLR ;
   OutputImg4(326) <= OutputImg4_326_EXMPLR ;
   OutputImg4(325) <= OutputImg4_325_EXMPLR ;
   OutputImg4(324) <= OutputImg4_324_EXMPLR ;
   OutputImg4(323) <= OutputImg4_323_EXMPLR ;
   OutputImg4(322) <= OutputImg4_322_EXMPLR ;
   OutputImg4(321) <= OutputImg4_321_EXMPLR ;
   OutputImg4(320) <= OutputImg4_320_EXMPLR ;
   OutputImg4(319) <= OutputImg4_319_EXMPLR ;
   OutputImg4(318) <= OutputImg4_318_EXMPLR ;
   OutputImg4(317) <= OutputImg4_317_EXMPLR ;
   OutputImg4(316) <= OutputImg4_316_EXMPLR ;
   OutputImg4(315) <= OutputImg4_315_EXMPLR ;
   OutputImg4(314) <= OutputImg4_314_EXMPLR ;
   OutputImg4(313) <= OutputImg4_313_EXMPLR ;
   OutputImg4(312) <= OutputImg4_312_EXMPLR ;
   OutputImg4(311) <= OutputImg4_311_EXMPLR ;
   OutputImg4(310) <= OutputImg4_310_EXMPLR ;
   OutputImg4(309) <= OutputImg4_309_EXMPLR ;
   OutputImg4(308) <= OutputImg4_308_EXMPLR ;
   OutputImg4(307) <= OutputImg4_307_EXMPLR ;
   OutputImg4(306) <= OutputImg4_306_EXMPLR ;
   OutputImg4(305) <= OutputImg4_305_EXMPLR ;
   OutputImg4(304) <= OutputImg4_304_EXMPLR ;
   OutputImg4(303) <= OutputImg4_303_EXMPLR ;
   OutputImg4(302) <= OutputImg4_302_EXMPLR ;
   OutputImg4(301) <= OutputImg4_301_EXMPLR ;
   OutputImg4(300) <= OutputImg4_300_EXMPLR ;
   OutputImg4(299) <= OutputImg4_299_EXMPLR ;
   OutputImg4(298) <= OutputImg4_298_EXMPLR ;
   OutputImg4(297) <= OutputImg4_297_EXMPLR ;
   OutputImg4(296) <= OutputImg4_296_EXMPLR ;
   OutputImg4(295) <= OutputImg4_295_EXMPLR ;
   OutputImg4(294) <= OutputImg4_294_EXMPLR ;
   OutputImg4(293) <= OutputImg4_293_EXMPLR ;
   OutputImg4(292) <= OutputImg4_292_EXMPLR ;
   OutputImg4(291) <= OutputImg4_291_EXMPLR ;
   OutputImg4(290) <= OutputImg4_290_EXMPLR ;
   OutputImg4(289) <= OutputImg4_289_EXMPLR ;
   OutputImg4(288) <= OutputImg4_288_EXMPLR ;
   OutputImg4(287) <= OutputImg4_287_EXMPLR ;
   OutputImg4(286) <= OutputImg4_286_EXMPLR ;
   OutputImg4(285) <= OutputImg4_285_EXMPLR ;
   OutputImg4(284) <= OutputImg4_284_EXMPLR ;
   OutputImg4(283) <= OutputImg4_283_EXMPLR ;
   OutputImg4(282) <= OutputImg4_282_EXMPLR ;
   OutputImg4(281) <= OutputImg4_281_EXMPLR ;
   OutputImg4(280) <= OutputImg4_280_EXMPLR ;
   OutputImg4(279) <= OutputImg4_279_EXMPLR ;
   OutputImg4(278) <= OutputImg4_278_EXMPLR ;
   OutputImg4(277) <= OutputImg4_277_EXMPLR ;
   OutputImg4(276) <= OutputImg4_276_EXMPLR ;
   OutputImg4(275) <= OutputImg4_275_EXMPLR ;
   OutputImg4(274) <= OutputImg4_274_EXMPLR ;
   OutputImg4(273) <= OutputImg4_273_EXMPLR ;
   OutputImg4(272) <= OutputImg4_272_EXMPLR ;
   OutputImg4(271) <= OutputImg4_271_EXMPLR ;
   OutputImg4(270) <= OutputImg4_270_EXMPLR ;
   OutputImg4(269) <= OutputImg4_269_EXMPLR ;
   OutputImg4(268) <= OutputImg4_268_EXMPLR ;
   OutputImg4(267) <= OutputImg4_267_EXMPLR ;
   OutputImg4(266) <= OutputImg4_266_EXMPLR ;
   OutputImg4(265) <= OutputImg4_265_EXMPLR ;
   OutputImg4(264) <= OutputImg4_264_EXMPLR ;
   OutputImg4(263) <= OutputImg4_263_EXMPLR ;
   OutputImg4(262) <= OutputImg4_262_EXMPLR ;
   OutputImg4(261) <= OutputImg4_261_EXMPLR ;
   OutputImg4(260) <= OutputImg4_260_EXMPLR ;
   OutputImg4(259) <= OutputImg4_259_EXMPLR ;
   OutputImg4(258) <= OutputImg4_258_EXMPLR ;
   OutputImg4(257) <= OutputImg4_257_EXMPLR ;
   OutputImg4(256) <= OutputImg4_256_EXMPLR ;
   OutputImg4(255) <= OutputImg4_255_EXMPLR ;
   OutputImg4(254) <= OutputImg4_254_EXMPLR ;
   OutputImg4(253) <= OutputImg4_253_EXMPLR ;
   OutputImg4(252) <= OutputImg4_252_EXMPLR ;
   OutputImg4(251) <= OutputImg4_251_EXMPLR ;
   OutputImg4(250) <= OutputImg4_250_EXMPLR ;
   OutputImg4(249) <= OutputImg4_249_EXMPLR ;
   OutputImg4(248) <= OutputImg4_248_EXMPLR ;
   OutputImg4(247) <= OutputImg4_247_EXMPLR ;
   OutputImg4(246) <= OutputImg4_246_EXMPLR ;
   OutputImg4(245) <= OutputImg4_245_EXMPLR ;
   OutputImg4(244) <= OutputImg4_244_EXMPLR ;
   OutputImg4(243) <= OutputImg4_243_EXMPLR ;
   OutputImg4(242) <= OutputImg4_242_EXMPLR ;
   OutputImg4(241) <= OutputImg4_241_EXMPLR ;
   OutputImg4(240) <= OutputImg4_240_EXMPLR ;
   OutputImg4(239) <= OutputImg4_239_EXMPLR ;
   OutputImg4(238) <= OutputImg4_238_EXMPLR ;
   OutputImg4(237) <= OutputImg4_237_EXMPLR ;
   OutputImg4(236) <= OutputImg4_236_EXMPLR ;
   OutputImg4(235) <= OutputImg4_235_EXMPLR ;
   OutputImg4(234) <= OutputImg4_234_EXMPLR ;
   OutputImg4(233) <= OutputImg4_233_EXMPLR ;
   OutputImg4(232) <= OutputImg4_232_EXMPLR ;
   OutputImg4(231) <= OutputImg4_231_EXMPLR ;
   OutputImg4(230) <= OutputImg4_230_EXMPLR ;
   OutputImg4(229) <= OutputImg4_229_EXMPLR ;
   OutputImg4(228) <= OutputImg4_228_EXMPLR ;
   OutputImg4(227) <= OutputImg4_227_EXMPLR ;
   OutputImg4(226) <= OutputImg4_226_EXMPLR ;
   OutputImg4(225) <= OutputImg4_225_EXMPLR ;
   OutputImg4(224) <= OutputImg4_224_EXMPLR ;
   OutputImg4(223) <= OutputImg4_223_EXMPLR ;
   OutputImg4(222) <= OutputImg4_222_EXMPLR ;
   OutputImg4(221) <= OutputImg4_221_EXMPLR ;
   OutputImg4(220) <= OutputImg4_220_EXMPLR ;
   OutputImg4(219) <= OutputImg4_219_EXMPLR ;
   OutputImg4(218) <= OutputImg4_218_EXMPLR ;
   OutputImg4(217) <= OutputImg4_217_EXMPLR ;
   OutputImg4(216) <= OutputImg4_216_EXMPLR ;
   OutputImg4(215) <= OutputImg4_215_EXMPLR ;
   OutputImg4(214) <= OutputImg4_214_EXMPLR ;
   OutputImg4(213) <= OutputImg4_213_EXMPLR ;
   OutputImg4(212) <= OutputImg4_212_EXMPLR ;
   OutputImg4(211) <= OutputImg4_211_EXMPLR ;
   OutputImg4(210) <= OutputImg4_210_EXMPLR ;
   OutputImg4(209) <= OutputImg4_209_EXMPLR ;
   OutputImg4(208) <= OutputImg4_208_EXMPLR ;
   OutputImg4(207) <= OutputImg4_207_EXMPLR ;
   OutputImg4(206) <= OutputImg4_206_EXMPLR ;
   OutputImg4(205) <= OutputImg4_205_EXMPLR ;
   OutputImg4(204) <= OutputImg4_204_EXMPLR ;
   OutputImg4(203) <= OutputImg4_203_EXMPLR ;
   OutputImg4(202) <= OutputImg4_202_EXMPLR ;
   OutputImg4(201) <= OutputImg4_201_EXMPLR ;
   OutputImg4(200) <= OutputImg4_200_EXMPLR ;
   OutputImg4(199) <= OutputImg4_199_EXMPLR ;
   OutputImg4(198) <= OutputImg4_198_EXMPLR ;
   OutputImg4(197) <= OutputImg4_197_EXMPLR ;
   OutputImg4(196) <= OutputImg4_196_EXMPLR ;
   OutputImg4(195) <= OutputImg4_195_EXMPLR ;
   OutputImg4(194) <= OutputImg4_194_EXMPLR ;
   OutputImg4(193) <= OutputImg4_193_EXMPLR ;
   OutputImg4(192) <= OutputImg4_192_EXMPLR ;
   OutputImg4(191) <= OutputImg4_191_EXMPLR ;
   OutputImg4(190) <= OutputImg4_190_EXMPLR ;
   OutputImg4(189) <= OutputImg4_189_EXMPLR ;
   OutputImg4(188) <= OutputImg4_188_EXMPLR ;
   OutputImg4(187) <= OutputImg4_187_EXMPLR ;
   OutputImg4(186) <= OutputImg4_186_EXMPLR ;
   OutputImg4(185) <= OutputImg4_185_EXMPLR ;
   OutputImg4(184) <= OutputImg4_184_EXMPLR ;
   OutputImg4(183) <= OutputImg4_183_EXMPLR ;
   OutputImg4(182) <= OutputImg4_182_EXMPLR ;
   OutputImg4(181) <= OutputImg4_181_EXMPLR ;
   OutputImg4(180) <= OutputImg4_180_EXMPLR ;
   OutputImg4(179) <= OutputImg4_179_EXMPLR ;
   OutputImg4(178) <= OutputImg4_178_EXMPLR ;
   OutputImg4(177) <= OutputImg4_177_EXMPLR ;
   OutputImg4(176) <= OutputImg4_176_EXMPLR ;
   OutputImg4(175) <= OutputImg4_175_EXMPLR ;
   OutputImg4(174) <= OutputImg4_174_EXMPLR ;
   OutputImg4(173) <= OutputImg4_173_EXMPLR ;
   OutputImg4(172) <= OutputImg4_172_EXMPLR ;
   OutputImg4(171) <= OutputImg4_171_EXMPLR ;
   OutputImg4(170) <= OutputImg4_170_EXMPLR ;
   OutputImg4(169) <= OutputImg4_169_EXMPLR ;
   OutputImg4(168) <= OutputImg4_168_EXMPLR ;
   OutputImg4(167) <= OutputImg4_167_EXMPLR ;
   OutputImg4(166) <= OutputImg4_166_EXMPLR ;
   OutputImg4(165) <= OutputImg4_165_EXMPLR ;
   OutputImg4(164) <= OutputImg4_164_EXMPLR ;
   OutputImg4(163) <= OutputImg4_163_EXMPLR ;
   OutputImg4(162) <= OutputImg4_162_EXMPLR ;
   OutputImg4(161) <= OutputImg4_161_EXMPLR ;
   OutputImg4(160) <= OutputImg4_160_EXMPLR ;
   OutputImg4(159) <= OutputImg4_159_EXMPLR ;
   OutputImg4(158) <= OutputImg4_158_EXMPLR ;
   OutputImg4(157) <= OutputImg4_157_EXMPLR ;
   OutputImg4(156) <= OutputImg4_156_EXMPLR ;
   OutputImg4(155) <= OutputImg4_155_EXMPLR ;
   OutputImg4(154) <= OutputImg4_154_EXMPLR ;
   OutputImg4(153) <= OutputImg4_153_EXMPLR ;
   OutputImg4(152) <= OutputImg4_152_EXMPLR ;
   OutputImg4(151) <= OutputImg4_151_EXMPLR ;
   OutputImg4(150) <= OutputImg4_150_EXMPLR ;
   OutputImg4(149) <= OutputImg4_149_EXMPLR ;
   OutputImg4(148) <= OutputImg4_148_EXMPLR ;
   OutputImg4(147) <= OutputImg4_147_EXMPLR ;
   OutputImg4(146) <= OutputImg4_146_EXMPLR ;
   OutputImg4(145) <= OutputImg4_145_EXMPLR ;
   OutputImg4(144) <= OutputImg4_144_EXMPLR ;
   OutputImg4(143) <= OutputImg4_143_EXMPLR ;
   OutputImg4(142) <= OutputImg4_142_EXMPLR ;
   OutputImg4(141) <= OutputImg4_141_EXMPLR ;
   OutputImg4(140) <= OutputImg4_140_EXMPLR ;
   OutputImg4(139) <= OutputImg4_139_EXMPLR ;
   OutputImg4(138) <= OutputImg4_138_EXMPLR ;
   OutputImg4(137) <= OutputImg4_137_EXMPLR ;
   OutputImg4(136) <= OutputImg4_136_EXMPLR ;
   OutputImg4(135) <= OutputImg4_135_EXMPLR ;
   OutputImg4(134) <= OutputImg4_134_EXMPLR ;
   OutputImg4(133) <= OutputImg4_133_EXMPLR ;
   OutputImg4(132) <= OutputImg4_132_EXMPLR ;
   OutputImg4(131) <= OutputImg4_131_EXMPLR ;
   OutputImg4(130) <= OutputImg4_130_EXMPLR ;
   OutputImg4(129) <= OutputImg4_129_EXMPLR ;
   OutputImg4(128) <= OutputImg4_128_EXMPLR ;
   OutputImg4(127) <= OutputImg4_127_EXMPLR ;
   OutputImg4(126) <= OutputImg4_126_EXMPLR ;
   OutputImg4(125) <= OutputImg4_125_EXMPLR ;
   OutputImg4(124) <= OutputImg4_124_EXMPLR ;
   OutputImg4(123) <= OutputImg4_123_EXMPLR ;
   OutputImg4(122) <= OutputImg4_122_EXMPLR ;
   OutputImg4(121) <= OutputImg4_121_EXMPLR ;
   OutputImg4(120) <= OutputImg4_120_EXMPLR ;
   OutputImg4(119) <= OutputImg4_119_EXMPLR ;
   OutputImg4(118) <= OutputImg4_118_EXMPLR ;
   OutputImg4(117) <= OutputImg4_117_EXMPLR ;
   OutputImg4(116) <= OutputImg4_116_EXMPLR ;
   OutputImg4(115) <= OutputImg4_115_EXMPLR ;
   OutputImg4(114) <= OutputImg4_114_EXMPLR ;
   OutputImg4(113) <= OutputImg4_113_EXMPLR ;
   OutputImg4(112) <= OutputImg4_112_EXMPLR ;
   OutputImg4(111) <= OutputImg4_111_EXMPLR ;
   OutputImg4(110) <= OutputImg4_110_EXMPLR ;
   OutputImg4(109) <= OutputImg4_109_EXMPLR ;
   OutputImg4(108) <= OutputImg4_108_EXMPLR ;
   OutputImg4(107) <= OutputImg4_107_EXMPLR ;
   OutputImg4(106) <= OutputImg4_106_EXMPLR ;
   OutputImg4(105) <= OutputImg4_105_EXMPLR ;
   OutputImg4(104) <= OutputImg4_104_EXMPLR ;
   OutputImg4(103) <= OutputImg4_103_EXMPLR ;
   OutputImg4(102) <= OutputImg4_102_EXMPLR ;
   OutputImg4(101) <= OutputImg4_101_EXMPLR ;
   OutputImg4(100) <= OutputImg4_100_EXMPLR ;
   OutputImg4(99) <= OutputImg4_99_EXMPLR ;
   OutputImg4(98) <= OutputImg4_98_EXMPLR ;
   OutputImg4(97) <= OutputImg4_97_EXMPLR ;
   OutputImg4(96) <= OutputImg4_96_EXMPLR ;
   OutputImg4(95) <= OutputImg4_95_EXMPLR ;
   OutputImg4(94) <= OutputImg4_94_EXMPLR ;
   OutputImg4(93) <= OutputImg4_93_EXMPLR ;
   OutputImg4(92) <= OutputImg4_92_EXMPLR ;
   OutputImg4(91) <= OutputImg4_91_EXMPLR ;
   OutputImg4(90) <= OutputImg4_90_EXMPLR ;
   OutputImg4(89) <= OutputImg4_89_EXMPLR ;
   OutputImg4(88) <= OutputImg4_88_EXMPLR ;
   OutputImg4(87) <= OutputImg4_87_EXMPLR ;
   OutputImg4(86) <= OutputImg4_86_EXMPLR ;
   OutputImg4(85) <= OutputImg4_85_EXMPLR ;
   OutputImg4(84) <= OutputImg4_84_EXMPLR ;
   OutputImg4(83) <= OutputImg4_83_EXMPLR ;
   OutputImg4(82) <= OutputImg4_82_EXMPLR ;
   OutputImg4(81) <= OutputImg4_81_EXMPLR ;
   OutputImg4(80) <= OutputImg4_80_EXMPLR ;
   OutputImg4(79) <= OutputImg4_79_EXMPLR ;
   OutputImg4(78) <= OutputImg4_78_EXMPLR ;
   OutputImg4(77) <= OutputImg4_77_EXMPLR ;
   OutputImg4(76) <= OutputImg4_76_EXMPLR ;
   OutputImg4(75) <= OutputImg4_75_EXMPLR ;
   OutputImg4(74) <= OutputImg4_74_EXMPLR ;
   OutputImg4(73) <= OutputImg4_73_EXMPLR ;
   OutputImg4(72) <= OutputImg4_72_EXMPLR ;
   OutputImg4(71) <= OutputImg4_71_EXMPLR ;
   OutputImg4(70) <= OutputImg4_70_EXMPLR ;
   OutputImg4(69) <= OutputImg4_69_EXMPLR ;
   OutputImg4(68) <= OutputImg4_68_EXMPLR ;
   OutputImg4(67) <= OutputImg4_67_EXMPLR ;
   OutputImg4(66) <= OutputImg4_66_EXMPLR ;
   OutputImg4(65) <= OutputImg4_65_EXMPLR ;
   OutputImg4(64) <= OutputImg4_64_EXMPLR ;
   OutputImg4(63) <= OutputImg4_63_EXMPLR ;
   OutputImg4(62) <= OutputImg4_62_EXMPLR ;
   OutputImg4(61) <= OutputImg4_61_EXMPLR ;
   OutputImg4(60) <= OutputImg4_60_EXMPLR ;
   OutputImg4(59) <= OutputImg4_59_EXMPLR ;
   OutputImg4(58) <= OutputImg4_58_EXMPLR ;
   OutputImg4(57) <= OutputImg4_57_EXMPLR ;
   OutputImg4(56) <= OutputImg4_56_EXMPLR ;
   OutputImg4(55) <= OutputImg4_55_EXMPLR ;
   OutputImg4(54) <= OutputImg4_54_EXMPLR ;
   OutputImg4(53) <= OutputImg4_53_EXMPLR ;
   OutputImg4(52) <= OutputImg4_52_EXMPLR ;
   OutputImg4(51) <= OutputImg4_51_EXMPLR ;
   OutputImg4(50) <= OutputImg4_50_EXMPLR ;
   OutputImg4(49) <= OutputImg4_49_EXMPLR ;
   OutputImg4(48) <= OutputImg4_48_EXMPLR ;
   OutputImg4(47) <= OutputImg4_47_EXMPLR ;
   OutputImg4(46) <= OutputImg4_46_EXMPLR ;
   OutputImg4(45) <= OutputImg4_45_EXMPLR ;
   OutputImg4(44) <= OutputImg4_44_EXMPLR ;
   OutputImg4(43) <= OutputImg4_43_EXMPLR ;
   OutputImg4(42) <= OutputImg4_42_EXMPLR ;
   OutputImg4(41) <= OutputImg4_41_EXMPLR ;
   OutputImg4(40) <= OutputImg4_40_EXMPLR ;
   OutputImg4(39) <= OutputImg4_39_EXMPLR ;
   OutputImg4(38) <= OutputImg4_38_EXMPLR ;
   OutputImg4(37) <= OutputImg4_37_EXMPLR ;
   OutputImg4(36) <= OutputImg4_36_EXMPLR ;
   OutputImg4(35) <= OutputImg4_35_EXMPLR ;
   OutputImg4(34) <= OutputImg4_34_EXMPLR ;
   OutputImg4(33) <= OutputImg4_33_EXMPLR ;
   OutputImg4(32) <= OutputImg4_32_EXMPLR ;
   OutputImg4(31) <= OutputImg4_31_EXMPLR ;
   OutputImg4(30) <= OutputImg4_30_EXMPLR ;
   OutputImg4(29) <= OutputImg4_29_EXMPLR ;
   OutputImg4(28) <= OutputImg4_28_EXMPLR ;
   OutputImg4(27) <= OutputImg4_27_EXMPLR ;
   OutputImg4(26) <= OutputImg4_26_EXMPLR ;
   OutputImg4(25) <= OutputImg4_25_EXMPLR ;
   OutputImg4(24) <= OutputImg4_24_EXMPLR ;
   OutputImg4(23) <= OutputImg4_23_EXMPLR ;
   OutputImg4(22) <= OutputImg4_22_EXMPLR ;
   OutputImg4(21) <= OutputImg4_21_EXMPLR ;
   OutputImg4(20) <= OutputImg4_20_EXMPLR ;
   OutputImg4(19) <= OutputImg4_19_EXMPLR ;
   OutputImg4(18) <= OutputImg4_18_EXMPLR ;
   OutputImg4(17) <= OutputImg4_17_EXMPLR ;
   OutputImg4(16) <= OutputImg4_16_EXMPLR ;
   OutputImg4(15) <= OutputImg4_15_EXMPLR ;
   OutputImg4(14) <= OutputImg4_14_EXMPLR ;
   OutputImg4(13) <= OutputImg4_13_EXMPLR ;
   OutputImg4(12) <= OutputImg4_12_EXMPLR ;
   OutputImg4(11) <= OutputImg4_11_EXMPLR ;
   OutputImg4(10) <= OutputImg4_10_EXMPLR ;
   OutputImg4(9) <= OutputImg4_9_EXMPLR ;
   OutputImg4(8) <= OutputImg4_8_EXMPLR ;
   OutputImg4(7) <= OutputImg4_7_EXMPLR ;
   OutputImg4(6) <= OutputImg4_6_EXMPLR ;
   OutputImg4(5) <= OutputImg4_5_EXMPLR ;
   OutputImg4(4) <= OutputImg4_4_EXMPLR ;
   OutputImg4(3) <= OutputImg4_3_EXMPLR ;
   OutputImg4(2) <= OutputImg4_2_EXMPLR ;
   OutputImg4(1) <= OutputImg4_1_EXMPLR ;
   OutputImg4(0) <= OutputImg4_0_EXMPLR ;
   OutputImg5(447) <= OutputImg5_447_EXMPLR ;
   OutputImg5(446) <= OutputImg5_446_EXMPLR ;
   OutputImg5(445) <= OutputImg5_445_EXMPLR ;
   OutputImg5(444) <= OutputImg5_444_EXMPLR ;
   OutputImg5(443) <= OutputImg5_443_EXMPLR ;
   OutputImg5(442) <= OutputImg5_442_EXMPLR ;
   OutputImg5(441) <= OutputImg5_441_EXMPLR ;
   OutputImg5(440) <= OutputImg5_440_EXMPLR ;
   OutputImg5(439) <= OutputImg5_439_EXMPLR ;
   OutputImg5(438) <= OutputImg5_438_EXMPLR ;
   OutputImg5(437) <= OutputImg5_437_EXMPLR ;
   OutputImg5(436) <= OutputImg5_436_EXMPLR ;
   OutputImg5(435) <= OutputImg5_435_EXMPLR ;
   OutputImg5(434) <= OutputImg5_434_EXMPLR ;
   OutputImg5(433) <= OutputImg5_433_EXMPLR ;
   OutputImg5(432) <= OutputImg5_432_EXMPLR ;
   OutputImg5(431) <= OutputImg5_431_EXMPLR ;
   OutputImg5(430) <= OutputImg5_430_EXMPLR ;
   OutputImg5(429) <= OutputImg5_429_EXMPLR ;
   OutputImg5(428) <= OutputImg5_428_EXMPLR ;
   OutputImg5(427) <= OutputImg5_427_EXMPLR ;
   OutputImg5(426) <= OutputImg5_426_EXMPLR ;
   OutputImg5(425) <= OutputImg5_425_EXMPLR ;
   OutputImg5(424) <= OutputImg5_424_EXMPLR ;
   OutputImg5(423) <= OutputImg5_423_EXMPLR ;
   OutputImg5(422) <= OutputImg5_422_EXMPLR ;
   OutputImg5(421) <= OutputImg5_421_EXMPLR ;
   OutputImg5(420) <= OutputImg5_420_EXMPLR ;
   OutputImg5(419) <= OutputImg5_419_EXMPLR ;
   OutputImg5(418) <= OutputImg5_418_EXMPLR ;
   OutputImg5(417) <= OutputImg5_417_EXMPLR ;
   OutputImg5(416) <= OutputImg5_416_EXMPLR ;
   OutputImg5(415) <= OutputImg5_415_EXMPLR ;
   OutputImg5(414) <= OutputImg5_414_EXMPLR ;
   OutputImg5(413) <= OutputImg5_413_EXMPLR ;
   OutputImg5(412) <= OutputImg5_412_EXMPLR ;
   OutputImg5(411) <= OutputImg5_411_EXMPLR ;
   OutputImg5(410) <= OutputImg5_410_EXMPLR ;
   OutputImg5(409) <= OutputImg5_409_EXMPLR ;
   OutputImg5(408) <= OutputImg5_408_EXMPLR ;
   OutputImg5(407) <= OutputImg5_407_EXMPLR ;
   OutputImg5(406) <= OutputImg5_406_EXMPLR ;
   OutputImg5(405) <= OutputImg5_405_EXMPLR ;
   OutputImg5(404) <= OutputImg5_404_EXMPLR ;
   OutputImg5(403) <= OutputImg5_403_EXMPLR ;
   OutputImg5(402) <= OutputImg5_402_EXMPLR ;
   OutputImg5(401) <= OutputImg5_401_EXMPLR ;
   OutputImg5(400) <= OutputImg5_400_EXMPLR ;
   OutputImg5(399) <= OutputImg5_399_EXMPLR ;
   OutputImg5(398) <= OutputImg5_398_EXMPLR ;
   OutputImg5(397) <= OutputImg5_397_EXMPLR ;
   OutputImg5(396) <= OutputImg5_396_EXMPLR ;
   OutputImg5(395) <= OutputImg5_395_EXMPLR ;
   OutputImg5(394) <= OutputImg5_394_EXMPLR ;
   OutputImg5(393) <= OutputImg5_393_EXMPLR ;
   OutputImg5(392) <= OutputImg5_392_EXMPLR ;
   OutputImg5(391) <= OutputImg5_391_EXMPLR ;
   OutputImg5(390) <= OutputImg5_390_EXMPLR ;
   OutputImg5(389) <= OutputImg5_389_EXMPLR ;
   OutputImg5(388) <= OutputImg5_388_EXMPLR ;
   OutputImg5(387) <= OutputImg5_387_EXMPLR ;
   OutputImg5(386) <= OutputImg5_386_EXMPLR ;
   OutputImg5(385) <= OutputImg5_385_EXMPLR ;
   OutputImg5(384) <= OutputImg5_384_EXMPLR ;
   OutputImg5(383) <= OutputImg5_383_EXMPLR ;
   OutputImg5(382) <= OutputImg5_382_EXMPLR ;
   OutputImg5(381) <= OutputImg5_381_EXMPLR ;
   OutputImg5(380) <= OutputImg5_380_EXMPLR ;
   OutputImg5(379) <= OutputImg5_379_EXMPLR ;
   OutputImg5(378) <= OutputImg5_378_EXMPLR ;
   OutputImg5(377) <= OutputImg5_377_EXMPLR ;
   OutputImg5(376) <= OutputImg5_376_EXMPLR ;
   OutputImg5(375) <= OutputImg5_375_EXMPLR ;
   OutputImg5(374) <= OutputImg5_374_EXMPLR ;
   OutputImg5(373) <= OutputImg5_373_EXMPLR ;
   OutputImg5(372) <= OutputImg5_372_EXMPLR ;
   OutputImg5(371) <= OutputImg5_371_EXMPLR ;
   OutputImg5(370) <= OutputImg5_370_EXMPLR ;
   OutputImg5(369) <= OutputImg5_369_EXMPLR ;
   OutputImg5(368) <= OutputImg5_368_EXMPLR ;
   OutputImg5(367) <= OutputImg5_367_EXMPLR ;
   OutputImg5(366) <= OutputImg5_366_EXMPLR ;
   OutputImg5(365) <= OutputImg5_365_EXMPLR ;
   OutputImg5(364) <= OutputImg5_364_EXMPLR ;
   OutputImg5(363) <= OutputImg5_363_EXMPLR ;
   OutputImg5(362) <= OutputImg5_362_EXMPLR ;
   OutputImg5(361) <= OutputImg5_361_EXMPLR ;
   OutputImg5(360) <= OutputImg5_360_EXMPLR ;
   OutputImg5(359) <= OutputImg5_359_EXMPLR ;
   OutputImg5(358) <= OutputImg5_358_EXMPLR ;
   OutputImg5(357) <= OutputImg5_357_EXMPLR ;
   OutputImg5(356) <= OutputImg5_356_EXMPLR ;
   OutputImg5(355) <= OutputImg5_355_EXMPLR ;
   OutputImg5(354) <= OutputImg5_354_EXMPLR ;
   OutputImg5(353) <= OutputImg5_353_EXMPLR ;
   OutputImg5(352) <= OutputImg5_352_EXMPLR ;
   OutputImg5(351) <= OutputImg5_351_EXMPLR ;
   OutputImg5(350) <= OutputImg5_350_EXMPLR ;
   OutputImg5(349) <= OutputImg5_349_EXMPLR ;
   OutputImg5(348) <= OutputImg5_348_EXMPLR ;
   OutputImg5(347) <= OutputImg5_347_EXMPLR ;
   OutputImg5(346) <= OutputImg5_346_EXMPLR ;
   OutputImg5(345) <= OutputImg5_345_EXMPLR ;
   OutputImg5(344) <= OutputImg5_344_EXMPLR ;
   OutputImg5(343) <= OutputImg5_343_EXMPLR ;
   OutputImg5(342) <= OutputImg5_342_EXMPLR ;
   OutputImg5(341) <= OutputImg5_341_EXMPLR ;
   OutputImg5(340) <= OutputImg5_340_EXMPLR ;
   OutputImg5(339) <= OutputImg5_339_EXMPLR ;
   OutputImg5(338) <= OutputImg5_338_EXMPLR ;
   OutputImg5(337) <= OutputImg5_337_EXMPLR ;
   OutputImg5(336) <= OutputImg5_336_EXMPLR ;
   OutputImg5(335) <= OutputImg5_335_EXMPLR ;
   OutputImg5(334) <= OutputImg5_334_EXMPLR ;
   OutputImg5(333) <= OutputImg5_333_EXMPLR ;
   OutputImg5(332) <= OutputImg5_332_EXMPLR ;
   OutputImg5(331) <= OutputImg5_331_EXMPLR ;
   OutputImg5(330) <= OutputImg5_330_EXMPLR ;
   OutputImg5(329) <= OutputImg5_329_EXMPLR ;
   OutputImg5(328) <= OutputImg5_328_EXMPLR ;
   OutputImg5(327) <= OutputImg5_327_EXMPLR ;
   OutputImg5(326) <= OutputImg5_326_EXMPLR ;
   OutputImg5(325) <= OutputImg5_325_EXMPLR ;
   OutputImg5(324) <= OutputImg5_324_EXMPLR ;
   OutputImg5(323) <= OutputImg5_323_EXMPLR ;
   OutputImg5(322) <= OutputImg5_322_EXMPLR ;
   OutputImg5(321) <= OutputImg5_321_EXMPLR ;
   OutputImg5(320) <= OutputImg5_320_EXMPLR ;
   OutputImg5(319) <= OutputImg5_319_EXMPLR ;
   OutputImg5(318) <= OutputImg5_318_EXMPLR ;
   OutputImg5(317) <= OutputImg5_317_EXMPLR ;
   OutputImg5(316) <= OutputImg5_316_EXMPLR ;
   OutputImg5(315) <= OutputImg5_315_EXMPLR ;
   OutputImg5(314) <= OutputImg5_314_EXMPLR ;
   OutputImg5(313) <= OutputImg5_313_EXMPLR ;
   OutputImg5(312) <= OutputImg5_312_EXMPLR ;
   OutputImg5(311) <= OutputImg5_311_EXMPLR ;
   OutputImg5(310) <= OutputImg5_310_EXMPLR ;
   OutputImg5(309) <= OutputImg5_309_EXMPLR ;
   OutputImg5(308) <= OutputImg5_308_EXMPLR ;
   OutputImg5(307) <= OutputImg5_307_EXMPLR ;
   OutputImg5(306) <= OutputImg5_306_EXMPLR ;
   OutputImg5(305) <= OutputImg5_305_EXMPLR ;
   OutputImg5(304) <= OutputImg5_304_EXMPLR ;
   OutputImg5(303) <= OutputImg5_303_EXMPLR ;
   OutputImg5(302) <= OutputImg5_302_EXMPLR ;
   OutputImg5(301) <= OutputImg5_301_EXMPLR ;
   OutputImg5(300) <= OutputImg5_300_EXMPLR ;
   OutputImg5(299) <= OutputImg5_299_EXMPLR ;
   OutputImg5(298) <= OutputImg5_298_EXMPLR ;
   OutputImg5(297) <= OutputImg5_297_EXMPLR ;
   OutputImg5(296) <= OutputImg5_296_EXMPLR ;
   OutputImg5(295) <= OutputImg5_295_EXMPLR ;
   OutputImg5(294) <= OutputImg5_294_EXMPLR ;
   OutputImg5(293) <= OutputImg5_293_EXMPLR ;
   OutputImg5(292) <= OutputImg5_292_EXMPLR ;
   OutputImg5(291) <= OutputImg5_291_EXMPLR ;
   OutputImg5(290) <= OutputImg5_290_EXMPLR ;
   OutputImg5(289) <= OutputImg5_289_EXMPLR ;
   OutputImg5(288) <= OutputImg5_288_EXMPLR ;
   OutputImg5(287) <= OutputImg5_287_EXMPLR ;
   OutputImg5(286) <= OutputImg5_286_EXMPLR ;
   OutputImg5(285) <= OutputImg5_285_EXMPLR ;
   OutputImg5(284) <= OutputImg5_284_EXMPLR ;
   OutputImg5(283) <= OutputImg5_283_EXMPLR ;
   OutputImg5(282) <= OutputImg5_282_EXMPLR ;
   OutputImg5(281) <= OutputImg5_281_EXMPLR ;
   OutputImg5(280) <= OutputImg5_280_EXMPLR ;
   OutputImg5(279) <= OutputImg5_279_EXMPLR ;
   OutputImg5(278) <= OutputImg5_278_EXMPLR ;
   OutputImg5(277) <= OutputImg5_277_EXMPLR ;
   OutputImg5(276) <= OutputImg5_276_EXMPLR ;
   OutputImg5(275) <= OutputImg5_275_EXMPLR ;
   OutputImg5(274) <= OutputImg5_274_EXMPLR ;
   OutputImg5(273) <= OutputImg5_273_EXMPLR ;
   OutputImg5(272) <= OutputImg5_272_EXMPLR ;
   OutputImg5(271) <= OutputImg5_271_EXMPLR ;
   OutputImg5(270) <= OutputImg5_270_EXMPLR ;
   OutputImg5(269) <= OutputImg5_269_EXMPLR ;
   OutputImg5(268) <= OutputImg5_268_EXMPLR ;
   OutputImg5(267) <= OutputImg5_267_EXMPLR ;
   OutputImg5(266) <= OutputImg5_266_EXMPLR ;
   OutputImg5(265) <= OutputImg5_265_EXMPLR ;
   OutputImg5(264) <= OutputImg5_264_EXMPLR ;
   OutputImg5(263) <= OutputImg5_263_EXMPLR ;
   OutputImg5(262) <= OutputImg5_262_EXMPLR ;
   OutputImg5(261) <= OutputImg5_261_EXMPLR ;
   OutputImg5(260) <= OutputImg5_260_EXMPLR ;
   OutputImg5(259) <= OutputImg5_259_EXMPLR ;
   OutputImg5(258) <= OutputImg5_258_EXMPLR ;
   OutputImg5(257) <= OutputImg5_257_EXMPLR ;
   OutputImg5(256) <= OutputImg5_256_EXMPLR ;
   OutputImg5(255) <= OutputImg5_255_EXMPLR ;
   OutputImg5(254) <= OutputImg5_254_EXMPLR ;
   OutputImg5(253) <= OutputImg5_253_EXMPLR ;
   OutputImg5(252) <= OutputImg5_252_EXMPLR ;
   OutputImg5(251) <= OutputImg5_251_EXMPLR ;
   OutputImg5(250) <= OutputImg5_250_EXMPLR ;
   OutputImg5(249) <= OutputImg5_249_EXMPLR ;
   OutputImg5(248) <= OutputImg5_248_EXMPLR ;
   OutputImg5(247) <= OutputImg5_247_EXMPLR ;
   OutputImg5(246) <= OutputImg5_246_EXMPLR ;
   OutputImg5(245) <= OutputImg5_245_EXMPLR ;
   OutputImg5(244) <= OutputImg5_244_EXMPLR ;
   OutputImg5(243) <= OutputImg5_243_EXMPLR ;
   OutputImg5(242) <= OutputImg5_242_EXMPLR ;
   OutputImg5(241) <= OutputImg5_241_EXMPLR ;
   OutputImg5(240) <= OutputImg5_240_EXMPLR ;
   OutputImg5(239) <= OutputImg5_239_EXMPLR ;
   OutputImg5(238) <= OutputImg5_238_EXMPLR ;
   OutputImg5(237) <= OutputImg5_237_EXMPLR ;
   OutputImg5(236) <= OutputImg5_236_EXMPLR ;
   OutputImg5(235) <= OutputImg5_235_EXMPLR ;
   OutputImg5(234) <= OutputImg5_234_EXMPLR ;
   OutputImg5(233) <= OutputImg5_233_EXMPLR ;
   OutputImg5(232) <= OutputImg5_232_EXMPLR ;
   OutputImg5(231) <= OutputImg5_231_EXMPLR ;
   OutputImg5(230) <= OutputImg5_230_EXMPLR ;
   OutputImg5(229) <= OutputImg5_229_EXMPLR ;
   OutputImg5(228) <= OutputImg5_228_EXMPLR ;
   OutputImg5(227) <= OutputImg5_227_EXMPLR ;
   OutputImg5(226) <= OutputImg5_226_EXMPLR ;
   OutputImg5(225) <= OutputImg5_225_EXMPLR ;
   OutputImg5(224) <= OutputImg5_224_EXMPLR ;
   OutputImg5(223) <= OutputImg5_223_EXMPLR ;
   OutputImg5(222) <= OutputImg5_222_EXMPLR ;
   OutputImg5(221) <= OutputImg5_221_EXMPLR ;
   OutputImg5(220) <= OutputImg5_220_EXMPLR ;
   OutputImg5(219) <= OutputImg5_219_EXMPLR ;
   OutputImg5(218) <= OutputImg5_218_EXMPLR ;
   OutputImg5(217) <= OutputImg5_217_EXMPLR ;
   OutputImg5(216) <= OutputImg5_216_EXMPLR ;
   OutputImg5(215) <= OutputImg5_215_EXMPLR ;
   OutputImg5(214) <= OutputImg5_214_EXMPLR ;
   OutputImg5(213) <= OutputImg5_213_EXMPLR ;
   OutputImg5(212) <= OutputImg5_212_EXMPLR ;
   OutputImg5(211) <= OutputImg5_211_EXMPLR ;
   OutputImg5(210) <= OutputImg5_210_EXMPLR ;
   OutputImg5(209) <= OutputImg5_209_EXMPLR ;
   OutputImg5(208) <= OutputImg5_208_EXMPLR ;
   OutputImg5(207) <= OutputImg5_207_EXMPLR ;
   OutputImg5(206) <= OutputImg5_206_EXMPLR ;
   OutputImg5(205) <= OutputImg5_205_EXMPLR ;
   OutputImg5(204) <= OutputImg5_204_EXMPLR ;
   OutputImg5(203) <= OutputImg5_203_EXMPLR ;
   OutputImg5(202) <= OutputImg5_202_EXMPLR ;
   OutputImg5(201) <= OutputImg5_201_EXMPLR ;
   OutputImg5(200) <= OutputImg5_200_EXMPLR ;
   OutputImg5(199) <= OutputImg5_199_EXMPLR ;
   OutputImg5(198) <= OutputImg5_198_EXMPLR ;
   OutputImg5(197) <= OutputImg5_197_EXMPLR ;
   OutputImg5(196) <= OutputImg5_196_EXMPLR ;
   OutputImg5(195) <= OutputImg5_195_EXMPLR ;
   OutputImg5(194) <= OutputImg5_194_EXMPLR ;
   OutputImg5(193) <= OutputImg5_193_EXMPLR ;
   OutputImg5(192) <= OutputImg5_192_EXMPLR ;
   OutputImg5(191) <= OutputImg5_191_EXMPLR ;
   OutputImg5(190) <= OutputImg5_190_EXMPLR ;
   OutputImg5(189) <= OutputImg5_189_EXMPLR ;
   OutputImg5(188) <= OutputImg5_188_EXMPLR ;
   OutputImg5(187) <= OutputImg5_187_EXMPLR ;
   OutputImg5(186) <= OutputImg5_186_EXMPLR ;
   OutputImg5(185) <= OutputImg5_185_EXMPLR ;
   OutputImg5(184) <= OutputImg5_184_EXMPLR ;
   OutputImg5(183) <= OutputImg5_183_EXMPLR ;
   OutputImg5(182) <= OutputImg5_182_EXMPLR ;
   OutputImg5(181) <= OutputImg5_181_EXMPLR ;
   OutputImg5(180) <= OutputImg5_180_EXMPLR ;
   OutputImg5(179) <= OutputImg5_179_EXMPLR ;
   OutputImg5(178) <= OutputImg5_178_EXMPLR ;
   OutputImg5(177) <= OutputImg5_177_EXMPLR ;
   OutputImg5(176) <= OutputImg5_176_EXMPLR ;
   OutputImg5(175) <= OutputImg5_175_EXMPLR ;
   OutputImg5(174) <= OutputImg5_174_EXMPLR ;
   OutputImg5(173) <= OutputImg5_173_EXMPLR ;
   OutputImg5(172) <= OutputImg5_172_EXMPLR ;
   OutputImg5(171) <= OutputImg5_171_EXMPLR ;
   OutputImg5(170) <= OutputImg5_170_EXMPLR ;
   OutputImg5(169) <= OutputImg5_169_EXMPLR ;
   OutputImg5(168) <= OutputImg5_168_EXMPLR ;
   OutputImg5(167) <= OutputImg5_167_EXMPLR ;
   OutputImg5(166) <= OutputImg5_166_EXMPLR ;
   OutputImg5(165) <= OutputImg5_165_EXMPLR ;
   OutputImg5(164) <= OutputImg5_164_EXMPLR ;
   OutputImg5(163) <= OutputImg5_163_EXMPLR ;
   OutputImg5(162) <= OutputImg5_162_EXMPLR ;
   OutputImg5(161) <= OutputImg5_161_EXMPLR ;
   OutputImg5(160) <= OutputImg5_160_EXMPLR ;
   OutputImg5(159) <= OutputImg5_159_EXMPLR ;
   OutputImg5(158) <= OutputImg5_158_EXMPLR ;
   OutputImg5(157) <= OutputImg5_157_EXMPLR ;
   OutputImg5(156) <= OutputImg5_156_EXMPLR ;
   OutputImg5(155) <= OutputImg5_155_EXMPLR ;
   OutputImg5(154) <= OutputImg5_154_EXMPLR ;
   OutputImg5(153) <= OutputImg5_153_EXMPLR ;
   OutputImg5(152) <= OutputImg5_152_EXMPLR ;
   OutputImg5(151) <= OutputImg5_151_EXMPLR ;
   OutputImg5(150) <= OutputImg5_150_EXMPLR ;
   OutputImg5(149) <= OutputImg5_149_EXMPLR ;
   OutputImg5(148) <= OutputImg5_148_EXMPLR ;
   OutputImg5(147) <= OutputImg5_147_EXMPLR ;
   OutputImg5(146) <= OutputImg5_146_EXMPLR ;
   OutputImg5(145) <= OutputImg5_145_EXMPLR ;
   OutputImg5(144) <= OutputImg5_144_EXMPLR ;
   OutputImg5(143) <= OutputImg5_143_EXMPLR ;
   OutputImg5(142) <= OutputImg5_142_EXMPLR ;
   OutputImg5(141) <= OutputImg5_141_EXMPLR ;
   OutputImg5(140) <= OutputImg5_140_EXMPLR ;
   OutputImg5(139) <= OutputImg5_139_EXMPLR ;
   OutputImg5(138) <= OutputImg5_138_EXMPLR ;
   OutputImg5(137) <= OutputImg5_137_EXMPLR ;
   OutputImg5(136) <= OutputImg5_136_EXMPLR ;
   OutputImg5(135) <= OutputImg5_135_EXMPLR ;
   OutputImg5(134) <= OutputImg5_134_EXMPLR ;
   OutputImg5(133) <= OutputImg5_133_EXMPLR ;
   OutputImg5(132) <= OutputImg5_132_EXMPLR ;
   OutputImg5(131) <= OutputImg5_131_EXMPLR ;
   OutputImg5(130) <= OutputImg5_130_EXMPLR ;
   OutputImg5(129) <= OutputImg5_129_EXMPLR ;
   OutputImg5(128) <= OutputImg5_128_EXMPLR ;
   OutputImg5(127) <= OutputImg5_127_EXMPLR ;
   OutputImg5(126) <= OutputImg5_126_EXMPLR ;
   OutputImg5(125) <= OutputImg5_125_EXMPLR ;
   OutputImg5(124) <= OutputImg5_124_EXMPLR ;
   OutputImg5(123) <= OutputImg5_123_EXMPLR ;
   OutputImg5(122) <= OutputImg5_122_EXMPLR ;
   OutputImg5(121) <= OutputImg5_121_EXMPLR ;
   OutputImg5(120) <= OutputImg5_120_EXMPLR ;
   OutputImg5(119) <= OutputImg5_119_EXMPLR ;
   OutputImg5(118) <= OutputImg5_118_EXMPLR ;
   OutputImg5(117) <= OutputImg5_117_EXMPLR ;
   OutputImg5(116) <= OutputImg5_116_EXMPLR ;
   OutputImg5(115) <= OutputImg5_115_EXMPLR ;
   OutputImg5(114) <= OutputImg5_114_EXMPLR ;
   OutputImg5(113) <= OutputImg5_113_EXMPLR ;
   OutputImg5(112) <= OutputImg5_112_EXMPLR ;
   OutputImg5(111) <= OutputImg5_111_EXMPLR ;
   OutputImg5(110) <= OutputImg5_110_EXMPLR ;
   OutputImg5(109) <= OutputImg5_109_EXMPLR ;
   OutputImg5(108) <= OutputImg5_108_EXMPLR ;
   OutputImg5(107) <= OutputImg5_107_EXMPLR ;
   OutputImg5(106) <= OutputImg5_106_EXMPLR ;
   OutputImg5(105) <= OutputImg5_105_EXMPLR ;
   OutputImg5(104) <= OutputImg5_104_EXMPLR ;
   OutputImg5(103) <= OutputImg5_103_EXMPLR ;
   OutputImg5(102) <= OutputImg5_102_EXMPLR ;
   OutputImg5(101) <= OutputImg5_101_EXMPLR ;
   OutputImg5(100) <= OutputImg5_100_EXMPLR ;
   OutputImg5(99) <= OutputImg5_99_EXMPLR ;
   OutputImg5(98) <= OutputImg5_98_EXMPLR ;
   OutputImg5(97) <= OutputImg5_97_EXMPLR ;
   OutputImg5(96) <= OutputImg5_96_EXMPLR ;
   OutputImg5(95) <= OutputImg5_95_EXMPLR ;
   OutputImg5(94) <= OutputImg5_94_EXMPLR ;
   OutputImg5(93) <= OutputImg5_93_EXMPLR ;
   OutputImg5(92) <= OutputImg5_92_EXMPLR ;
   OutputImg5(91) <= OutputImg5_91_EXMPLR ;
   OutputImg5(90) <= OutputImg5_90_EXMPLR ;
   OutputImg5(89) <= OutputImg5_89_EXMPLR ;
   OutputImg5(88) <= OutputImg5_88_EXMPLR ;
   OutputImg5(87) <= OutputImg5_87_EXMPLR ;
   OutputImg5(86) <= OutputImg5_86_EXMPLR ;
   OutputImg5(85) <= OutputImg5_85_EXMPLR ;
   OutputImg5(84) <= OutputImg5_84_EXMPLR ;
   OutputImg5(83) <= OutputImg5_83_EXMPLR ;
   OutputImg5(82) <= OutputImg5_82_EXMPLR ;
   OutputImg5(81) <= OutputImg5_81_EXMPLR ;
   OutputImg5(80) <= OutputImg5_80_EXMPLR ;
   OutputImg5(79) <= OutputImg5_79_EXMPLR ;
   OutputImg5(78) <= OutputImg5_78_EXMPLR ;
   OutputImg5(77) <= OutputImg5_77_EXMPLR ;
   OutputImg5(76) <= OutputImg5_76_EXMPLR ;
   OutputImg5(75) <= OutputImg5_75_EXMPLR ;
   OutputImg5(74) <= OutputImg5_74_EXMPLR ;
   OutputImg5(73) <= OutputImg5_73_EXMPLR ;
   OutputImg5(72) <= OutputImg5_72_EXMPLR ;
   OutputImg5(71) <= OutputImg5_71_EXMPLR ;
   OutputImg5(70) <= OutputImg5_70_EXMPLR ;
   OutputImg5(69) <= OutputImg5_69_EXMPLR ;
   OutputImg5(68) <= OutputImg5_68_EXMPLR ;
   OutputImg5(67) <= OutputImg5_67_EXMPLR ;
   OutputImg5(66) <= OutputImg5_66_EXMPLR ;
   OutputImg5(65) <= OutputImg5_65_EXMPLR ;
   OutputImg5(64) <= OutputImg5_64_EXMPLR ;
   OutputImg5(63) <= OutputImg5_63_EXMPLR ;
   OutputImg5(62) <= OutputImg5_62_EXMPLR ;
   OutputImg5(61) <= OutputImg5_61_EXMPLR ;
   OutputImg5(60) <= OutputImg5_60_EXMPLR ;
   OutputImg5(59) <= OutputImg5_59_EXMPLR ;
   OutputImg5(58) <= OutputImg5_58_EXMPLR ;
   OutputImg5(57) <= OutputImg5_57_EXMPLR ;
   OutputImg5(56) <= OutputImg5_56_EXMPLR ;
   OutputImg5(55) <= OutputImg5_55_EXMPLR ;
   OutputImg5(54) <= OutputImg5_54_EXMPLR ;
   OutputImg5(53) <= OutputImg5_53_EXMPLR ;
   OutputImg5(52) <= OutputImg5_52_EXMPLR ;
   OutputImg5(51) <= OutputImg5_51_EXMPLR ;
   OutputImg5(50) <= OutputImg5_50_EXMPLR ;
   OutputImg5(49) <= OutputImg5_49_EXMPLR ;
   OutputImg5(48) <= OutputImg5_48_EXMPLR ;
   OutputImg5(47) <= OutputImg5_47_EXMPLR ;
   OutputImg5(46) <= OutputImg5_46_EXMPLR ;
   OutputImg5(45) <= OutputImg5_45_EXMPLR ;
   OutputImg5(44) <= OutputImg5_44_EXMPLR ;
   OutputImg5(43) <= OutputImg5_43_EXMPLR ;
   OutputImg5(42) <= OutputImg5_42_EXMPLR ;
   OutputImg5(41) <= OutputImg5_41_EXMPLR ;
   OutputImg5(40) <= OutputImg5_40_EXMPLR ;
   OutputImg5(39) <= OutputImg5_39_EXMPLR ;
   OutputImg5(38) <= OutputImg5_38_EXMPLR ;
   OutputImg5(37) <= OutputImg5_37_EXMPLR ;
   OutputImg5(36) <= OutputImg5_36_EXMPLR ;
   OutputImg5(35) <= OutputImg5_35_EXMPLR ;
   OutputImg5(34) <= OutputImg5_34_EXMPLR ;
   OutputImg5(33) <= OutputImg5_33_EXMPLR ;
   OutputImg5(32) <= OutputImg5_32_EXMPLR ;
   OutputImg5(31) <= OutputImg5_31_EXMPLR ;
   OutputImg5(30) <= OutputImg5_30_EXMPLR ;
   OutputImg5(29) <= OutputImg5_29_EXMPLR ;
   OutputImg5(28) <= OutputImg5_28_EXMPLR ;
   OutputImg5(27) <= OutputImg5_27_EXMPLR ;
   OutputImg5(26) <= OutputImg5_26_EXMPLR ;
   OutputImg5(25) <= OutputImg5_25_EXMPLR ;
   OutputImg5(24) <= OutputImg5_24_EXMPLR ;
   OutputImg5(23) <= OutputImg5_23_EXMPLR ;
   OutputImg5(22) <= OutputImg5_22_EXMPLR ;
   OutputImg5(21) <= OutputImg5_21_EXMPLR ;
   OutputImg5(20) <= OutputImg5_20_EXMPLR ;
   OutputImg5(19) <= OutputImg5_19_EXMPLR ;
   OutputImg5(18) <= OutputImg5_18_EXMPLR ;
   OutputImg5(17) <= OutputImg5_17_EXMPLR ;
   OutputImg5(16) <= OutputImg5_16_EXMPLR ;
   OutputImg5(15) <= OutputImg5_15_EXMPLR ;
   OutputImg5(14) <= OutputImg5_14_EXMPLR ;
   OutputImg5(13) <= OutputImg5_13_EXMPLR ;
   OutputImg5(12) <= OutputImg5_12_EXMPLR ;
   OutputImg5(11) <= OutputImg5_11_EXMPLR ;
   OutputImg5(10) <= OutputImg5_10_EXMPLR ;
   OutputImg5(9) <= OutputImg5_9_EXMPLR ;
   OutputImg5(8) <= OutputImg5_8_EXMPLR ;
   OutputImg5(7) <= OutputImg5_7_EXMPLR ;
   OutputImg5(6) <= OutputImg5_6_EXMPLR ;
   OutputImg5(5) <= OutputImg5_5_EXMPLR ;
   OutputImg5(4) <= OutputImg5_4_EXMPLR ;
   OutputImg5(3) <= OutputImg5_3_EXMPLR ;
   OutputImg5(2) <= OutputImg5_2_EXMPLR ;
   OutputImg5(1) <= OutputImg5_1_EXMPLR ;
   OutputImg5(0) <= OutputImg5_0_EXMPLR ;
   ImgCounterOuput(2) <= ImgCounterOuput_2_EXMPLR ;
   ImgCounterOuput(1) <= ImgCounterOuput_1_EXMPLR ;
   ImgCounterOuput(0) <= ImgCounterOuput_0_EXMPLR ;
   ImgIndic(0) <= ImgIndic_0_EXMPLR ;
   ImgEn(5) <= ImgEn_5_EXMPLR ;
   ImgEn(4) <= ImgEn_4_EXMPLR ;
   ImgEn(3) <= ImgEn_3_EXMPLR ;
   ImgEn(2) <= ImgEn_2_EXMPLR ;
   ImgEn(1) <= ImgEn_1_EXMPLR ;
   ImgEn(0) <= ImgEn_0_EXMPLR ;
   adder0 : my_nadder_16 port map ( a(15)=>firstOperand_15, a(14)=>
      firstOperand_15, a(13)=>firstOperand_15, a(12)=>ImgAddress(12), a(11)
      =>ImgAddress(11), a(10)=>ImgAddress(10), a(9)=>ImgAddress(9), a(8)=>
      ImgAddress(8), a(7)=>ImgAddress(7), a(6)=>ImgAddress(6), a(5)=>
      ImgAddress(5), a(4)=>ImgAddress(4), a(3)=>ImgAddress(3), a(2)=>
      ImgAddress(2), a(1)=>ImgAddress(1), a(0)=>ImgAddress(0), b(15)=>
      ImgWidth(15), b(14)=>ImgWidth(14), b(13)=>ImgWidth(13), b(12)=>
      ImgWidth(12), b(11)=>ImgWidth(11), b(10)=>ImgWidth(10), b(9)=>
      ImgWidth(9), b(8)=>ImgWidth(8), b(7)=>ImgWidth(7), b(6)=>ImgWidth(6), 
      b(5)=>ImgWidth(5), b(4)=>ImgWidth(4), b(3)=>ImgWidth(3), b(2)=>
      ImgWidth(2), b(1)=>ImgWidth(1), b(0)=>ImgWidth(0), cin=>
      firstOperand_15, s(15)=>DANGLING(0), s(14)=>DANGLING(1), s(13)=>
      DANGLING(2), s(12)=>newAdd16_12, s(11)=>newAdd16_11, s(10)=>
      newAdd16_10, s(9)=>newAdd16_9, s(8)=>newAdd16_8, s(7)=>newAdd16_7, 
      s(6)=>newAdd16_6, s(5)=>newAdd16_5, s(4)=>newAdd16_4, s(3)=>newAdd16_3, 
      s(2)=>newAdd16_2, s(1)=>newAdd16_1, s(0)=>newAdd16_0, cout=>DANGLING(3
      ));
   triStateAdd : triStateBuffer_13 port map ( D(12)=>newAdd16_12, D(11)=>
      newAdd16_11, D(10)=>newAdd16_10, D(9)=>newAdd16_9, D(8)=>newAdd16_8, 
      D(7)=>newAdd16_7, D(6)=>newAdd16_6, D(5)=>newAdd16_5, D(4)=>newAdd16_4, 
      D(3)=>newAdd16_3, D(2)=>newAdd16_2, D(1)=>newAdd16_1, D(0)=>newAdd16_0, 
      EN=>TriAddEn, F(12)=>UpdatedAddress(12), F(11)=>UpdatedAddress(11), 
      F(10)=>UpdatedAddress(10), F(9)=>UpdatedAddress(9), F(8)=>
      UpdatedAddress(8), F(7)=>UpdatedAddress(7), F(6)=>UpdatedAddress(6), 
      F(5)=>UpdatedAddress(5), F(4)=>UpdatedAddress(4), F(3)=>
      UpdatedAddress(3), F(2)=>UpdatedAddress(2), F(1)=>UpdatedAddress(1), 
      F(0)=>UpdatedAddress(0));
   TriStateAddToDma : triStateBuffer_13 port map ( D(12)=>ImgAddress(12), 
      D(11)=>ImgAddress(11), D(10)=>ImgAddress(10), D(9)=>ImgAddress(9), 
      D(8)=>ImgAddress(8), D(7)=>ImgAddress(7), D(6)=>ImgAddress(6), D(5)=>
      ImgAddress(5), D(4)=>ImgAddress(4), D(3)=>ImgAddress(3), D(2)=>
      ImgAddress(2), D(1)=>ImgAddress(1), D(0)=>ImgAddress(0), EN=>TriAddEn, 
      F(12)=>ImgAddToDma(12), F(11)=>ImgAddToDma(11), F(10)=>ImgAddToDma(10), 
      F(9)=>ImgAddToDma(9), F(8)=>ImgAddToDma(8), F(7)=>ImgAddToDma(7), F(6)
      =>ImgAddToDma(6), F(5)=>ImgAddToDma(5), F(4)=>ImgAddToDma(4), F(3)=>
      ImgAddToDma(3), F(2)=>ImgAddToDma(2), F(1)=>ImgAddToDma(1), F(0)=>
      ImgAddToDma(0));
   DDF0 : nBitRegister_1 port map ( D(0)=>NOT_ImgIndic_0, CLK=>DFFCLK, RST=>
      IndRst, EN=>PWR, Q(0)=>ImgIndic_0_EXMPLR);
   RegCounter0 : Counter_3 port map ( enable=>cEnable, reset=>cReset, clk=>
      nx23828, load=>firstOperand_15, output(2)=>ImgCounterOuput_2_EXMPLR, 
      output(1)=>ImgCounterOuput_1_EXMPLR, output(0)=>
      ImgCounterOuput_0_EXMPLR, input(2)=>firstOperand_15, input(1)=>
      firstOperand_15, input(0)=>PWR);
   dec : Decoder port map ( input(2)=>ImgCounterOuput_2_EXMPLR, input(1)=>
      ImgCounterOuput_1_EXMPLR, input(0)=>ImgCounterOuput_0_EXMPLR, 
      output(5)=>DecOutput_5, output(4)=>DecOutput_4, output(3)=>DecOutput_3, 
      output(2)=>DecOutput_2, output(1)=>DecOutput_1, output(0)=>DecOutput_0
   );
   TriImgReg : triStateBuffer_6 port map ( D(5)=>DecOutput_5, D(4)=>
      DecOutput_4, D(3)=>DecOutput_3, D(2)=>DecOutput_2, D(1)=>DecOutput_1, 
      D(0)=>DecOutput_0, EN=>TriImgRegEn, F(5)=>ImgEn_5_EXMPLR, F(4)=>
      ImgEn_4_EXMPLR, F(3)=>ImgEn_3_EXMPLR, F(2)=>ImgEn_2_EXMPLR, F(1)=>
      ImgEn_1_EXMPLR, F(0)=>ImgEn_0_EXMPLR);
   loop3_0_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_31_EXMPLR, D(14)=>OutputImg0_30_EXMPLR, D(13)=>
      OutputImg0_29_EXMPLR, D(12)=>OutputImg0_28_EXMPLR, D(11)=>
      OutputImg0_27_EXMPLR, D(10)=>OutputImg0_26_EXMPLR, D(9)=>
      OutputImg0_25_EXMPLR, D(8)=>OutputImg0_24_EXMPLR, D(7)=>
      OutputImg0_23_EXMPLR, D(6)=>OutputImg0_22_EXMPLR, D(5)=>
      OutputImg0_21_EXMPLR, D(4)=>OutputImg0_20_EXMPLR, D(3)=>
      OutputImg0_19_EXMPLR, D(2)=>OutputImg0_18_EXMPLR, D(1)=>
      OutputImg0_17_EXMPLR, D(0)=>OutputImg0_16_EXMPLR, EN=>nx23666, F(15)=>
      ImgReg0IN_15, F(14)=>ImgReg0IN_14, F(13)=>ImgReg0IN_13, F(12)=>
      ImgReg0IN_12, F(11)=>ImgReg0IN_11, F(10)=>ImgReg0IN_10, F(9)=>
      ImgReg0IN_9, F(8)=>ImgReg0IN_8, F(7)=>ImgReg0IN_7, F(6)=>ImgReg0IN_6, 
      F(5)=>ImgReg0IN_5, F(4)=>ImgReg0IN_4, F(3)=>ImgReg0IN_3, F(2)=>
      ImgReg0IN_2, F(1)=>ImgReg0IN_1, F(0)=>ImgReg0IN_0);
   loop3_0_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_31_EXMPLR, D(14)=>OutputImg1_30_EXMPLR, D(13)=>
      OutputImg1_29_EXMPLR, D(12)=>OutputImg1_28_EXMPLR, D(11)=>
      OutputImg1_27_EXMPLR, D(10)=>OutputImg1_26_EXMPLR, D(9)=>
      OutputImg1_25_EXMPLR, D(8)=>OutputImg1_24_EXMPLR, D(7)=>
      OutputImg1_23_EXMPLR, D(6)=>OutputImg1_22_EXMPLR, D(5)=>
      OutputImg1_21_EXMPLR, D(4)=>OutputImg1_20_EXMPLR, D(3)=>
      OutputImg1_19_EXMPLR, D(2)=>OutputImg1_18_EXMPLR, D(1)=>
      OutputImg1_17_EXMPLR, D(0)=>OutputImg1_16_EXMPLR, EN=>nx23666, F(15)=>
      ImgReg1IN_15, F(14)=>ImgReg1IN_14, F(13)=>ImgReg1IN_13, F(12)=>
      ImgReg1IN_12, F(11)=>ImgReg1IN_11, F(10)=>ImgReg1IN_10, F(9)=>
      ImgReg1IN_9, F(8)=>ImgReg1IN_8, F(7)=>ImgReg1IN_7, F(6)=>ImgReg1IN_6, 
      F(5)=>ImgReg1IN_5, F(4)=>ImgReg1IN_4, F(3)=>ImgReg1IN_3, F(2)=>
      ImgReg1IN_2, F(1)=>ImgReg1IN_1, F(0)=>ImgReg1IN_0);
   loop3_0_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_31_EXMPLR, D(14)=>OutputImg2_30_EXMPLR, D(13)=>
      OutputImg2_29_EXMPLR, D(12)=>OutputImg2_28_EXMPLR, D(11)=>
      OutputImg2_27_EXMPLR, D(10)=>OutputImg2_26_EXMPLR, D(9)=>
      OutputImg2_25_EXMPLR, D(8)=>OutputImg2_24_EXMPLR, D(7)=>
      OutputImg2_23_EXMPLR, D(6)=>OutputImg2_22_EXMPLR, D(5)=>
      OutputImg2_21_EXMPLR, D(4)=>OutputImg2_20_EXMPLR, D(3)=>
      OutputImg2_19_EXMPLR, D(2)=>OutputImg2_18_EXMPLR, D(1)=>
      OutputImg2_17_EXMPLR, D(0)=>OutputImg2_16_EXMPLR, EN=>nx23666, F(15)=>
      ImgReg2IN_15, F(14)=>ImgReg2IN_14, F(13)=>ImgReg2IN_13, F(12)=>
      ImgReg2IN_12, F(11)=>ImgReg2IN_11, F(10)=>ImgReg2IN_10, F(9)=>
      ImgReg2IN_9, F(8)=>ImgReg2IN_8, F(7)=>ImgReg2IN_7, F(6)=>ImgReg2IN_6, 
      F(5)=>ImgReg2IN_5, F(4)=>ImgReg2IN_4, F(3)=>ImgReg2IN_3, F(2)=>
      ImgReg2IN_2, F(1)=>ImgReg2IN_1, F(0)=>ImgReg2IN_0);
   loop3_0_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_31_EXMPLR, D(14)=>OutputImg3_30_EXMPLR, D(13)=>
      OutputImg3_29_EXMPLR, D(12)=>OutputImg3_28_EXMPLR, D(11)=>
      OutputImg3_27_EXMPLR, D(10)=>OutputImg3_26_EXMPLR, D(9)=>
      OutputImg3_25_EXMPLR, D(8)=>OutputImg3_24_EXMPLR, D(7)=>
      OutputImg3_23_EXMPLR, D(6)=>OutputImg3_22_EXMPLR, D(5)=>
      OutputImg3_21_EXMPLR, D(4)=>OutputImg3_20_EXMPLR, D(3)=>
      OutputImg3_19_EXMPLR, D(2)=>OutputImg3_18_EXMPLR, D(1)=>
      OutputImg3_17_EXMPLR, D(0)=>OutputImg3_16_EXMPLR, EN=>nx23666, F(15)=>
      ImgReg3IN_15, F(14)=>ImgReg3IN_14, F(13)=>ImgReg3IN_13, F(12)=>
      ImgReg3IN_12, F(11)=>ImgReg3IN_11, F(10)=>ImgReg3IN_10, F(9)=>
      ImgReg3IN_9, F(8)=>ImgReg3IN_8, F(7)=>ImgReg3IN_7, F(6)=>ImgReg3IN_6, 
      F(5)=>ImgReg3IN_5, F(4)=>ImgReg3IN_4, F(3)=>ImgReg3IN_3, F(2)=>
      ImgReg3IN_2, F(1)=>ImgReg3IN_1, F(0)=>ImgReg3IN_0);
   loop3_0_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_31_EXMPLR, D(14)=>OutputImg4_30_EXMPLR, D(13)=>
      OutputImg4_29_EXMPLR, D(12)=>OutputImg4_28_EXMPLR, D(11)=>
      OutputImg4_27_EXMPLR, D(10)=>OutputImg4_26_EXMPLR, D(9)=>
      OutputImg4_25_EXMPLR, D(8)=>OutputImg4_24_EXMPLR, D(7)=>
      OutputImg4_23_EXMPLR, D(6)=>OutputImg4_22_EXMPLR, D(5)=>
      OutputImg4_21_EXMPLR, D(4)=>OutputImg4_20_EXMPLR, D(3)=>
      OutputImg4_19_EXMPLR, D(2)=>OutputImg4_18_EXMPLR, D(1)=>
      OutputImg4_17_EXMPLR, D(0)=>OutputImg4_16_EXMPLR, EN=>nx23666, F(15)=>
      ImgReg4IN_15, F(14)=>ImgReg4IN_14, F(13)=>ImgReg4IN_13, F(12)=>
      ImgReg4IN_12, F(11)=>ImgReg4IN_11, F(10)=>ImgReg4IN_10, F(9)=>
      ImgReg4IN_9, F(8)=>ImgReg4IN_8, F(7)=>ImgReg4IN_7, F(6)=>ImgReg4IN_6, 
      F(5)=>ImgReg4IN_5, F(4)=>ImgReg4IN_4, F(3)=>ImgReg4IN_3, F(2)=>
      ImgReg4IN_2, F(1)=>ImgReg4IN_1, F(0)=>ImgReg4IN_0);
   loop3_0_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_31_EXMPLR, D(14)=>OutputImg5_30_EXMPLR, D(13)=>
      OutputImg5_29_EXMPLR, D(12)=>OutputImg5_28_EXMPLR, D(11)=>
      OutputImg5_27_EXMPLR, D(10)=>OutputImg5_26_EXMPLR, D(9)=>
      OutputImg5_25_EXMPLR, D(8)=>OutputImg5_24_EXMPLR, D(7)=>
      OutputImg5_23_EXMPLR, D(6)=>OutputImg5_22_EXMPLR, D(5)=>
      OutputImg5_21_EXMPLR, D(4)=>OutputImg5_20_EXMPLR, D(3)=>
      OutputImg5_19_EXMPLR, D(2)=>OutputImg5_18_EXMPLR, D(1)=>
      OutputImg5_17_EXMPLR, D(0)=>OutputImg5_16_EXMPLR, EN=>nx23666, F(15)=>
      ImgReg5IN_15, F(14)=>ImgReg5IN_14, F(13)=>ImgReg5IN_13, F(12)=>
      ImgReg5IN_12, F(11)=>ImgReg5IN_11, F(10)=>ImgReg5IN_10, F(9)=>
      ImgReg5IN_9, F(8)=>ImgReg5IN_8, F(7)=>ImgReg5IN_7, F(6)=>ImgReg5IN_6, 
      F(5)=>ImgReg5IN_5, F(4)=>ImgReg5IN_4, F(3)=>ImgReg5IN_3, F(2)=>
      ImgReg5IN_2, F(1)=>ImgReg5IN_1, F(0)=>ImgReg5IN_0);
   loop3_0_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(15), D(14)
      =>DATA(14), D(13)=>DATA(13), D(12)=>DATA(12), D(11)=>DATA(11), D(10)=>
      DATA(10), D(9)=>DATA(9), D(8)=>DATA(8), D(7)=>DATA(7), D(6)=>DATA(6), 
      D(5)=>DATA(5), D(4)=>DATA(4), D(3)=>DATA(3), D(2)=>DATA(2), D(1)=>
      DATA(1), D(0)=>DATA(0), EN=>nx23654, F(15)=>ImgReg0IN_15, F(14)=>
      ImgReg0IN_14, F(13)=>ImgReg0IN_13, F(12)=>ImgReg0IN_12, F(11)=>
      ImgReg0IN_11, F(10)=>ImgReg0IN_10, F(9)=>ImgReg0IN_9, F(8)=>
      ImgReg0IN_8, F(7)=>ImgReg0IN_7, F(6)=>ImgReg0IN_6, F(5)=>ImgReg0IN_5, 
      F(4)=>ImgReg0IN_4, F(3)=>ImgReg0IN_3, F(2)=>ImgReg0IN_2, F(1)=>
      ImgReg0IN_1, F(0)=>ImgReg0IN_0);
   loop3_0_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(15), D(14)
      =>DATA(14), D(13)=>DATA(13), D(12)=>DATA(12), D(11)=>DATA(11), D(10)=>
      DATA(10), D(9)=>DATA(9), D(8)=>DATA(8), D(7)=>DATA(7), D(6)=>DATA(6), 
      D(5)=>DATA(5), D(4)=>DATA(4), D(3)=>DATA(3), D(2)=>DATA(2), D(1)=>
      DATA(1), D(0)=>DATA(0), EN=>nx23642, F(15)=>ImgReg1IN_15, F(14)=>
      ImgReg1IN_14, F(13)=>ImgReg1IN_13, F(12)=>ImgReg1IN_12, F(11)=>
      ImgReg1IN_11, F(10)=>ImgReg1IN_10, F(9)=>ImgReg1IN_9, F(8)=>
      ImgReg1IN_8, F(7)=>ImgReg1IN_7, F(6)=>ImgReg1IN_6, F(5)=>ImgReg1IN_5, 
      F(4)=>ImgReg1IN_4, F(3)=>ImgReg1IN_3, F(2)=>ImgReg1IN_2, F(1)=>
      ImgReg1IN_1, F(0)=>ImgReg1IN_0);
   loop3_0_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(15), D(14)
      =>DATA(14), D(13)=>DATA(13), D(12)=>DATA(12), D(11)=>DATA(11), D(10)=>
      DATA(10), D(9)=>DATA(9), D(8)=>DATA(8), D(7)=>DATA(7), D(6)=>DATA(6), 
      D(5)=>DATA(5), D(4)=>DATA(4), D(3)=>DATA(3), D(2)=>DATA(2), D(1)=>
      DATA(1), D(0)=>DATA(0), EN=>nx23630, F(15)=>ImgReg2IN_15, F(14)=>
      ImgReg2IN_14, F(13)=>ImgReg2IN_13, F(12)=>ImgReg2IN_12, F(11)=>
      ImgReg2IN_11, F(10)=>ImgReg2IN_10, F(9)=>ImgReg2IN_9, F(8)=>
      ImgReg2IN_8, F(7)=>ImgReg2IN_7, F(6)=>ImgReg2IN_6, F(5)=>ImgReg2IN_5, 
      F(4)=>ImgReg2IN_4, F(3)=>ImgReg2IN_3, F(2)=>ImgReg2IN_2, F(1)=>
      ImgReg2IN_1, F(0)=>ImgReg2IN_0);
   loop3_0_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(15), D(14)
      =>DATA(14), D(13)=>DATA(13), D(12)=>DATA(12), D(11)=>DATA(11), D(10)=>
      DATA(10), D(9)=>DATA(9), D(8)=>DATA(8), D(7)=>DATA(7), D(6)=>DATA(6), 
      D(5)=>DATA(5), D(4)=>DATA(4), D(3)=>DATA(3), D(2)=>DATA(2), D(1)=>
      DATA(1), D(0)=>DATA(0), EN=>nx23618, F(15)=>ImgReg3IN_15, F(14)=>
      ImgReg3IN_14, F(13)=>ImgReg3IN_13, F(12)=>ImgReg3IN_12, F(11)=>
      ImgReg3IN_11, F(10)=>ImgReg3IN_10, F(9)=>ImgReg3IN_9, F(8)=>
      ImgReg3IN_8, F(7)=>ImgReg3IN_7, F(6)=>ImgReg3IN_6, F(5)=>ImgReg3IN_5, 
      F(4)=>ImgReg3IN_4, F(3)=>ImgReg3IN_3, F(2)=>ImgReg3IN_2, F(1)=>
      ImgReg3IN_1, F(0)=>ImgReg3IN_0);
   loop3_0_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(15), D(14)
      =>DATA(14), D(13)=>DATA(13), D(12)=>DATA(12), D(11)=>DATA(11), D(10)=>
      DATA(10), D(9)=>DATA(9), D(8)=>DATA(8), D(7)=>DATA(7), D(6)=>DATA(6), 
      D(5)=>DATA(5), D(4)=>DATA(4), D(3)=>DATA(3), D(2)=>DATA(2), D(1)=>
      DATA(1), D(0)=>DATA(0), EN=>nx23606, F(15)=>ImgReg4IN_15, F(14)=>
      ImgReg4IN_14, F(13)=>ImgReg4IN_13, F(12)=>ImgReg4IN_12, F(11)=>
      ImgReg4IN_11, F(10)=>ImgReg4IN_10, F(9)=>ImgReg4IN_9, F(8)=>
      ImgReg4IN_8, F(7)=>ImgReg4IN_7, F(6)=>ImgReg4IN_6, F(5)=>ImgReg4IN_5, 
      F(4)=>ImgReg4IN_4, F(3)=>ImgReg4IN_3, F(2)=>ImgReg4IN_2, F(1)=>
      ImgReg4IN_1, F(0)=>ImgReg4IN_0);
   loop3_0_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(15), D(14)
      =>DATA(14), D(13)=>DATA(13), D(12)=>DATA(12), D(11)=>DATA(11), D(10)=>
      DATA(10), D(9)=>DATA(9), D(8)=>DATA(8), D(7)=>DATA(7), D(6)=>DATA(6), 
      D(5)=>DATA(5), D(4)=>DATA(4), D(3)=>DATA(3), D(2)=>DATA(2), D(1)=>
      DATA(1), D(0)=>DATA(0), EN=>nx23594, F(15)=>ImgReg5IN_15, F(14)=>
      ImgReg5IN_14, F(13)=>ImgReg5IN_13, F(12)=>ImgReg5IN_12, F(11)=>
      ImgReg5IN_11, F(10)=>ImgReg5IN_10, F(9)=>ImgReg5IN_9, F(8)=>
      ImgReg5IN_8, F(7)=>ImgReg5IN_7, F(6)=>ImgReg5IN_6, F(5)=>ImgReg5IN_5, 
      F(4)=>ImgReg5IN_4, F(3)=>ImgReg5IN_3, F(2)=>ImgReg5IN_2, F(1)=>
      ImgReg5IN_1, F(0)=>ImgReg5IN_0);
   loop3_0_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_15_EXMPLR, D(14)=>OutputImg1_14_EXMPLR, D(13)=>
      OutputImg1_13_EXMPLR, D(12)=>OutputImg1_12_EXMPLR, D(11)=>
      OutputImg1_11_EXMPLR, D(10)=>OutputImg1_10_EXMPLR, D(9)=>
      OutputImg1_9_EXMPLR, D(8)=>OutputImg1_8_EXMPLR, D(7)=>
      OutputImg1_7_EXMPLR, D(6)=>OutputImg1_6_EXMPLR, D(5)=>
      OutputImg1_5_EXMPLR, D(4)=>OutputImg1_4_EXMPLR, D(3)=>
      OutputImg1_3_EXMPLR, D(2)=>OutputImg1_2_EXMPLR, D(1)=>
      OutputImg1_1_EXMPLR, D(0)=>OutputImg1_0_EXMPLR, EN=>nx23786, F(15)=>
      ImgReg0IN_15, F(14)=>ImgReg0IN_14, F(13)=>ImgReg0IN_13, F(12)=>
      ImgReg0IN_12, F(11)=>ImgReg0IN_11, F(10)=>ImgReg0IN_10, F(9)=>
      ImgReg0IN_9, F(8)=>ImgReg0IN_8, F(7)=>ImgReg0IN_7, F(6)=>ImgReg0IN_6, 
      F(5)=>ImgReg0IN_5, F(4)=>ImgReg0IN_4, F(3)=>ImgReg0IN_3, F(2)=>
      ImgReg0IN_2, F(1)=>ImgReg0IN_1, F(0)=>ImgReg0IN_0);
   loop3_0_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_15_EXMPLR, D(14)=>OutputImg2_14_EXMPLR, D(13)=>
      OutputImg2_13_EXMPLR, D(12)=>OutputImg2_12_EXMPLR, D(11)=>
      OutputImg2_11_EXMPLR, D(10)=>OutputImg2_10_EXMPLR, D(9)=>
      OutputImg2_9_EXMPLR, D(8)=>OutputImg2_8_EXMPLR, D(7)=>
      OutputImg2_7_EXMPLR, D(6)=>OutputImg2_6_EXMPLR, D(5)=>
      OutputImg2_5_EXMPLR, D(4)=>OutputImg2_4_EXMPLR, D(3)=>
      OutputImg2_3_EXMPLR, D(2)=>OutputImg2_2_EXMPLR, D(1)=>
      OutputImg2_1_EXMPLR, D(0)=>OutputImg2_0_EXMPLR, EN=>nx23786, F(15)=>
      ImgReg1IN_15, F(14)=>ImgReg1IN_14, F(13)=>ImgReg1IN_13, F(12)=>
      ImgReg1IN_12, F(11)=>ImgReg1IN_11, F(10)=>ImgReg1IN_10, F(9)=>
      ImgReg1IN_9, F(8)=>ImgReg1IN_8, F(7)=>ImgReg1IN_7, F(6)=>ImgReg1IN_6, 
      F(5)=>ImgReg1IN_5, F(4)=>ImgReg1IN_4, F(3)=>ImgReg1IN_3, F(2)=>
      ImgReg1IN_2, F(1)=>ImgReg1IN_1, F(0)=>ImgReg1IN_0);
   loop3_0_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_15_EXMPLR, D(14)=>OutputImg3_14_EXMPLR, D(13)=>
      OutputImg3_13_EXMPLR, D(12)=>OutputImg3_12_EXMPLR, D(11)=>
      OutputImg3_11_EXMPLR, D(10)=>OutputImg3_10_EXMPLR, D(9)=>
      OutputImg3_9_EXMPLR, D(8)=>OutputImg3_8_EXMPLR, D(7)=>
      OutputImg3_7_EXMPLR, D(6)=>OutputImg3_6_EXMPLR, D(5)=>
      OutputImg3_5_EXMPLR, D(4)=>OutputImg3_4_EXMPLR, D(3)=>
      OutputImg3_3_EXMPLR, D(2)=>OutputImg3_2_EXMPLR, D(1)=>
      OutputImg3_1_EXMPLR, D(0)=>OutputImg3_0_EXMPLR, EN=>nx23786, F(15)=>
      ImgReg2IN_15, F(14)=>ImgReg2IN_14, F(13)=>ImgReg2IN_13, F(12)=>
      ImgReg2IN_12, F(11)=>ImgReg2IN_11, F(10)=>ImgReg2IN_10, F(9)=>
      ImgReg2IN_9, F(8)=>ImgReg2IN_8, F(7)=>ImgReg2IN_7, F(6)=>ImgReg2IN_6, 
      F(5)=>ImgReg2IN_5, F(4)=>ImgReg2IN_4, F(3)=>ImgReg2IN_3, F(2)=>
      ImgReg2IN_2, F(1)=>ImgReg2IN_1, F(0)=>ImgReg2IN_0);
   loop3_0_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_15_EXMPLR, D(14)=>OutputImg4_14_EXMPLR, D(13)=>
      OutputImg4_13_EXMPLR, D(12)=>OutputImg4_12_EXMPLR, D(11)=>
      OutputImg4_11_EXMPLR, D(10)=>OutputImg4_10_EXMPLR, D(9)=>
      OutputImg4_9_EXMPLR, D(8)=>OutputImg4_8_EXMPLR, D(7)=>
      OutputImg4_7_EXMPLR, D(6)=>OutputImg4_6_EXMPLR, D(5)=>
      OutputImg4_5_EXMPLR, D(4)=>OutputImg4_4_EXMPLR, D(3)=>
      OutputImg4_3_EXMPLR, D(2)=>OutputImg4_2_EXMPLR, D(1)=>
      OutputImg4_1_EXMPLR, D(0)=>OutputImg4_0_EXMPLR, EN=>nx23786, F(15)=>
      ImgReg3IN_15, F(14)=>ImgReg3IN_14, F(13)=>ImgReg3IN_13, F(12)=>
      ImgReg3IN_12, F(11)=>ImgReg3IN_11, F(10)=>ImgReg3IN_10, F(9)=>
      ImgReg3IN_9, F(8)=>ImgReg3IN_8, F(7)=>ImgReg3IN_7, F(6)=>ImgReg3IN_6, 
      F(5)=>ImgReg3IN_5, F(4)=>ImgReg3IN_4, F(3)=>ImgReg3IN_3, F(2)=>
      ImgReg3IN_2, F(1)=>ImgReg3IN_1, F(0)=>ImgReg3IN_0);
   loop3_0_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_15_EXMPLR, D(14)=>OutputImg5_14_EXMPLR, D(13)=>
      OutputImg5_13_EXMPLR, D(12)=>OutputImg5_12_EXMPLR, D(11)=>
      OutputImg5_11_EXMPLR, D(10)=>OutputImg5_10_EXMPLR, D(9)=>
      OutputImg5_9_EXMPLR, D(8)=>OutputImg5_8_EXMPLR, D(7)=>
      OutputImg5_7_EXMPLR, D(6)=>OutputImg5_6_EXMPLR, D(5)=>
      OutputImg5_5_EXMPLR, D(4)=>OutputImg5_4_EXMPLR, D(3)=>
      OutputImg5_3_EXMPLR, D(2)=>OutputImg5_2_EXMPLR, D(1)=>
      OutputImg5_1_EXMPLR, D(0)=>OutputImg5_0_EXMPLR, EN=>nx23786, F(15)=>
      ImgReg4IN_15, F(14)=>ImgReg4IN_14, F(13)=>ImgReg4IN_13, F(12)=>
      ImgReg4IN_12, F(11)=>ImgReg4IN_11, F(10)=>ImgReg4IN_10, F(9)=>
      ImgReg4IN_9, F(8)=>ImgReg4IN_8, F(7)=>ImgReg4IN_7, F(6)=>ImgReg4IN_6, 
      F(5)=>ImgReg4IN_5, F(4)=>ImgReg4IN_4, F(3)=>ImgReg4IN_3, F(2)=>
      ImgReg4IN_2, F(1)=>ImgReg4IN_1, F(0)=>ImgReg4IN_0);
   loop3_0_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_15, D(14)=>
      ImgReg0IN_14, D(13)=>ImgReg0IN_13, D(12)=>ImgReg0IN_12, D(11)=>
      ImgReg0IN_11, D(10)=>ImgReg0IN_10, D(9)=>ImgReg0IN_9, D(8)=>
      ImgReg0IN_8, D(7)=>ImgReg0IN_7, D(6)=>ImgReg0IN_6, D(5)=>ImgReg0IN_5, 
      D(4)=>ImgReg0IN_4, D(3)=>ImgReg0IN_3, D(2)=>ImgReg0IN_2, D(1)=>
      ImgReg0IN_1, D(0)=>ImgReg0IN_0, CLK=>nx23828, RST=>RST, EN=>nx23718, 
      Q(15)=>OutputImg0_15_EXMPLR, Q(14)=>OutputImg0_14_EXMPLR, Q(13)=>
      OutputImg0_13_EXMPLR, Q(12)=>OutputImg0_12_EXMPLR, Q(11)=>
      OutputImg0_11_EXMPLR, Q(10)=>OutputImg0_10_EXMPLR, Q(9)=>
      OutputImg0_9_EXMPLR, Q(8)=>OutputImg0_8_EXMPLR, Q(7)=>
      OutputImg0_7_EXMPLR, Q(6)=>OutputImg0_6_EXMPLR, Q(5)=>
      OutputImg0_5_EXMPLR, Q(4)=>OutputImg0_4_EXMPLR, Q(3)=>
      OutputImg0_3_EXMPLR, Q(2)=>OutputImg0_2_EXMPLR, Q(1)=>
      OutputImg0_1_EXMPLR, Q(0)=>OutputImg0_0_EXMPLR);
   loop3_0_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_15, D(14)=>
      ImgReg1IN_14, D(13)=>ImgReg1IN_13, D(12)=>ImgReg1IN_12, D(11)=>
      ImgReg1IN_11, D(10)=>ImgReg1IN_10, D(9)=>ImgReg1IN_9, D(8)=>
      ImgReg1IN_8, D(7)=>ImgReg1IN_7, D(6)=>ImgReg1IN_6, D(5)=>ImgReg1IN_5, 
      D(4)=>ImgReg1IN_4, D(3)=>ImgReg1IN_3, D(2)=>ImgReg1IN_2, D(1)=>
      ImgReg1IN_1, D(0)=>ImgReg1IN_0, CLK=>nx23830, RST=>RST, EN=>nx23728, 
      Q(15)=>OutputImg1_15_EXMPLR, Q(14)=>OutputImg1_14_EXMPLR, Q(13)=>
      OutputImg1_13_EXMPLR, Q(12)=>OutputImg1_12_EXMPLR, Q(11)=>
      OutputImg1_11_EXMPLR, Q(10)=>OutputImg1_10_EXMPLR, Q(9)=>
      OutputImg1_9_EXMPLR, Q(8)=>OutputImg1_8_EXMPLR, Q(7)=>
      OutputImg1_7_EXMPLR, Q(6)=>OutputImg1_6_EXMPLR, Q(5)=>
      OutputImg1_5_EXMPLR, Q(4)=>OutputImg1_4_EXMPLR, Q(3)=>
      OutputImg1_3_EXMPLR, Q(2)=>OutputImg1_2_EXMPLR, Q(1)=>
      OutputImg1_1_EXMPLR, Q(0)=>OutputImg1_0_EXMPLR);
   loop3_0_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_15, D(14)=>
      ImgReg2IN_14, D(13)=>ImgReg2IN_13, D(12)=>ImgReg2IN_12, D(11)=>
      ImgReg2IN_11, D(10)=>ImgReg2IN_10, D(9)=>ImgReg2IN_9, D(8)=>
      ImgReg2IN_8, D(7)=>ImgReg2IN_7, D(6)=>ImgReg2IN_6, D(5)=>ImgReg2IN_5, 
      D(4)=>ImgReg2IN_4, D(3)=>ImgReg2IN_3, D(2)=>ImgReg2IN_2, D(1)=>
      ImgReg2IN_1, D(0)=>ImgReg2IN_0, CLK=>nx23830, RST=>RST, EN=>nx23738, 
      Q(15)=>OutputImg2_15_EXMPLR, Q(14)=>OutputImg2_14_EXMPLR, Q(13)=>
      OutputImg2_13_EXMPLR, Q(12)=>OutputImg2_12_EXMPLR, Q(11)=>
      OutputImg2_11_EXMPLR, Q(10)=>OutputImg2_10_EXMPLR, Q(9)=>
      OutputImg2_9_EXMPLR, Q(8)=>OutputImg2_8_EXMPLR, Q(7)=>
      OutputImg2_7_EXMPLR, Q(6)=>OutputImg2_6_EXMPLR, Q(5)=>
      OutputImg2_5_EXMPLR, Q(4)=>OutputImg2_4_EXMPLR, Q(3)=>
      OutputImg2_3_EXMPLR, Q(2)=>OutputImg2_2_EXMPLR, Q(1)=>
      OutputImg2_1_EXMPLR, Q(0)=>OutputImg2_0_EXMPLR);
   loop3_0_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_15, D(14)=>
      ImgReg3IN_14, D(13)=>ImgReg3IN_13, D(12)=>ImgReg3IN_12, D(11)=>
      ImgReg3IN_11, D(10)=>ImgReg3IN_10, D(9)=>ImgReg3IN_9, D(8)=>
      ImgReg3IN_8, D(7)=>ImgReg3IN_7, D(6)=>ImgReg3IN_6, D(5)=>ImgReg3IN_5, 
      D(4)=>ImgReg3IN_4, D(3)=>ImgReg3IN_3, D(2)=>ImgReg3IN_2, D(1)=>
      ImgReg3IN_1, D(0)=>ImgReg3IN_0, CLK=>nx23832, RST=>RST, EN=>nx23748, 
      Q(15)=>OutputImg3_15_EXMPLR, Q(14)=>OutputImg3_14_EXMPLR, Q(13)=>
      OutputImg3_13_EXMPLR, Q(12)=>OutputImg3_12_EXMPLR, Q(11)=>
      OutputImg3_11_EXMPLR, Q(10)=>OutputImg3_10_EXMPLR, Q(9)=>
      OutputImg3_9_EXMPLR, Q(8)=>OutputImg3_8_EXMPLR, Q(7)=>
      OutputImg3_7_EXMPLR, Q(6)=>OutputImg3_6_EXMPLR, Q(5)=>
      OutputImg3_5_EXMPLR, Q(4)=>OutputImg3_4_EXMPLR, Q(3)=>
      OutputImg3_3_EXMPLR, Q(2)=>OutputImg3_2_EXMPLR, Q(1)=>
      OutputImg3_1_EXMPLR, Q(0)=>OutputImg3_0_EXMPLR);
   loop3_0_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_15, D(14)=>
      ImgReg4IN_14, D(13)=>ImgReg4IN_13, D(12)=>ImgReg4IN_12, D(11)=>
      ImgReg4IN_11, D(10)=>ImgReg4IN_10, D(9)=>ImgReg4IN_9, D(8)=>
      ImgReg4IN_8, D(7)=>ImgReg4IN_7, D(6)=>ImgReg4IN_6, D(5)=>ImgReg4IN_5, 
      D(4)=>ImgReg4IN_4, D(3)=>ImgReg4IN_3, D(2)=>ImgReg4IN_2, D(1)=>
      ImgReg4IN_1, D(0)=>ImgReg4IN_0, CLK=>nx23832, RST=>RST, EN=>nx23758, 
      Q(15)=>OutputImg4_15_EXMPLR, Q(14)=>OutputImg4_14_EXMPLR, Q(13)=>
      OutputImg4_13_EXMPLR, Q(12)=>OutputImg4_12_EXMPLR, Q(11)=>
      OutputImg4_11_EXMPLR, Q(10)=>OutputImg4_10_EXMPLR, Q(9)=>
      OutputImg4_9_EXMPLR, Q(8)=>OutputImg4_8_EXMPLR, Q(7)=>
      OutputImg4_7_EXMPLR, Q(6)=>OutputImg4_6_EXMPLR, Q(5)=>
      OutputImg4_5_EXMPLR, Q(4)=>OutputImg4_4_EXMPLR, Q(3)=>
      OutputImg4_3_EXMPLR, Q(2)=>OutputImg4_2_EXMPLR, Q(1)=>
      OutputImg4_1_EXMPLR, Q(0)=>OutputImg4_0_EXMPLR);
   loop3_0_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_15, D(14)=>
      ImgReg5IN_14, D(13)=>ImgReg5IN_13, D(12)=>ImgReg5IN_12, D(11)=>
      ImgReg5IN_11, D(10)=>ImgReg5IN_10, D(9)=>ImgReg5IN_9, D(8)=>
      ImgReg5IN_8, D(7)=>ImgReg5IN_7, D(6)=>ImgReg5IN_6, D(5)=>ImgReg5IN_5, 
      D(4)=>ImgReg5IN_4, D(3)=>ImgReg5IN_3, D(2)=>ImgReg5IN_2, D(1)=>
      ImgReg5IN_1, D(0)=>ImgReg5IN_0, CLK=>nx23834, RST=>RST, EN=>nx23768, 
      Q(15)=>OutputImg5_15_EXMPLR, Q(14)=>OutputImg5_14_EXMPLR, Q(13)=>
      OutputImg5_13_EXMPLR, Q(12)=>OutputImg5_12_EXMPLR, Q(11)=>
      OutputImg5_11_EXMPLR, Q(10)=>OutputImg5_10_EXMPLR, Q(9)=>
      OutputImg5_9_EXMPLR, Q(8)=>OutputImg5_8_EXMPLR, Q(7)=>
      OutputImg5_7_EXMPLR, Q(6)=>OutputImg5_6_EXMPLR, Q(5)=>
      OutputImg5_5_EXMPLR, Q(4)=>OutputImg5_4_EXMPLR, Q(3)=>
      OutputImg5_3_EXMPLR, Q(2)=>OutputImg5_2_EXMPLR, Q(1)=>
      OutputImg5_1_EXMPLR, Q(0)=>OutputImg5_0_EXMPLR);
   loop3_1_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_47_EXMPLR, D(14)=>OutputImg0_46_EXMPLR, D(13)=>
      OutputImg0_45_EXMPLR, D(12)=>OutputImg0_44_EXMPLR, D(11)=>
      OutputImg0_43_EXMPLR, D(10)=>OutputImg0_42_EXMPLR, D(9)=>
      OutputImg0_41_EXMPLR, D(8)=>OutputImg0_40_EXMPLR, D(7)=>
      OutputImg0_39_EXMPLR, D(6)=>OutputImg0_38_EXMPLR, D(5)=>
      OutputImg0_37_EXMPLR, D(4)=>OutputImg0_36_EXMPLR, D(3)=>
      OutputImg0_35_EXMPLR, D(2)=>OutputImg0_34_EXMPLR, D(1)=>
      OutputImg0_33_EXMPLR, D(0)=>OutputImg0_32_EXMPLR, EN=>nx23666, F(15)=>
      ImgReg0IN_31, F(14)=>ImgReg0IN_30, F(13)=>ImgReg0IN_29, F(12)=>
      ImgReg0IN_28, F(11)=>ImgReg0IN_27, F(10)=>ImgReg0IN_26, F(9)=>
      ImgReg0IN_25, F(8)=>ImgReg0IN_24, F(7)=>ImgReg0IN_23, F(6)=>
      ImgReg0IN_22, F(5)=>ImgReg0IN_21, F(4)=>ImgReg0IN_20, F(3)=>
      ImgReg0IN_19, F(2)=>ImgReg0IN_18, F(1)=>ImgReg0IN_17, F(0)=>
      ImgReg0IN_16);
   loop3_1_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_47_EXMPLR, D(14)=>OutputImg1_46_EXMPLR, D(13)=>
      OutputImg1_45_EXMPLR, D(12)=>OutputImg1_44_EXMPLR, D(11)=>
      OutputImg1_43_EXMPLR, D(10)=>OutputImg1_42_EXMPLR, D(9)=>
      OutputImg1_41_EXMPLR, D(8)=>OutputImg1_40_EXMPLR, D(7)=>
      OutputImg1_39_EXMPLR, D(6)=>OutputImg1_38_EXMPLR, D(5)=>
      OutputImg1_37_EXMPLR, D(4)=>OutputImg1_36_EXMPLR, D(3)=>
      OutputImg1_35_EXMPLR, D(2)=>OutputImg1_34_EXMPLR, D(1)=>
      OutputImg1_33_EXMPLR, D(0)=>OutputImg1_32_EXMPLR, EN=>nx23668, F(15)=>
      ImgReg1IN_31, F(14)=>ImgReg1IN_30, F(13)=>ImgReg1IN_29, F(12)=>
      ImgReg1IN_28, F(11)=>ImgReg1IN_27, F(10)=>ImgReg1IN_26, F(9)=>
      ImgReg1IN_25, F(8)=>ImgReg1IN_24, F(7)=>ImgReg1IN_23, F(6)=>
      ImgReg1IN_22, F(5)=>ImgReg1IN_21, F(4)=>ImgReg1IN_20, F(3)=>
      ImgReg1IN_19, F(2)=>ImgReg1IN_18, F(1)=>ImgReg1IN_17, F(0)=>
      ImgReg1IN_16);
   loop3_1_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_47_EXMPLR, D(14)=>OutputImg2_46_EXMPLR, D(13)=>
      OutputImg2_45_EXMPLR, D(12)=>OutputImg2_44_EXMPLR, D(11)=>
      OutputImg2_43_EXMPLR, D(10)=>OutputImg2_42_EXMPLR, D(9)=>
      OutputImg2_41_EXMPLR, D(8)=>OutputImg2_40_EXMPLR, D(7)=>
      OutputImg2_39_EXMPLR, D(6)=>OutputImg2_38_EXMPLR, D(5)=>
      OutputImg2_37_EXMPLR, D(4)=>OutputImg2_36_EXMPLR, D(3)=>
      OutputImg2_35_EXMPLR, D(2)=>OutputImg2_34_EXMPLR, D(1)=>
      OutputImg2_33_EXMPLR, D(0)=>OutputImg2_32_EXMPLR, EN=>nx23668, F(15)=>
      ImgReg2IN_31, F(14)=>ImgReg2IN_30, F(13)=>ImgReg2IN_29, F(12)=>
      ImgReg2IN_28, F(11)=>ImgReg2IN_27, F(10)=>ImgReg2IN_26, F(9)=>
      ImgReg2IN_25, F(8)=>ImgReg2IN_24, F(7)=>ImgReg2IN_23, F(6)=>
      ImgReg2IN_22, F(5)=>ImgReg2IN_21, F(4)=>ImgReg2IN_20, F(3)=>
      ImgReg2IN_19, F(2)=>ImgReg2IN_18, F(1)=>ImgReg2IN_17, F(0)=>
      ImgReg2IN_16);
   loop3_1_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_47_EXMPLR, D(14)=>OutputImg3_46_EXMPLR, D(13)=>
      OutputImg3_45_EXMPLR, D(12)=>OutputImg3_44_EXMPLR, D(11)=>
      OutputImg3_43_EXMPLR, D(10)=>OutputImg3_42_EXMPLR, D(9)=>
      OutputImg3_41_EXMPLR, D(8)=>OutputImg3_40_EXMPLR, D(7)=>
      OutputImg3_39_EXMPLR, D(6)=>OutputImg3_38_EXMPLR, D(5)=>
      OutputImg3_37_EXMPLR, D(4)=>OutputImg3_36_EXMPLR, D(3)=>
      OutputImg3_35_EXMPLR, D(2)=>OutputImg3_34_EXMPLR, D(1)=>
      OutputImg3_33_EXMPLR, D(0)=>OutputImg3_32_EXMPLR, EN=>nx23668, F(15)=>
      ImgReg3IN_31, F(14)=>ImgReg3IN_30, F(13)=>ImgReg3IN_29, F(12)=>
      ImgReg3IN_28, F(11)=>ImgReg3IN_27, F(10)=>ImgReg3IN_26, F(9)=>
      ImgReg3IN_25, F(8)=>ImgReg3IN_24, F(7)=>ImgReg3IN_23, F(6)=>
      ImgReg3IN_22, F(5)=>ImgReg3IN_21, F(4)=>ImgReg3IN_20, F(3)=>
      ImgReg3IN_19, F(2)=>ImgReg3IN_18, F(1)=>ImgReg3IN_17, F(0)=>
      ImgReg3IN_16);
   loop3_1_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_47_EXMPLR, D(14)=>OutputImg4_46_EXMPLR, D(13)=>
      OutputImg4_45_EXMPLR, D(12)=>OutputImg4_44_EXMPLR, D(11)=>
      OutputImg4_43_EXMPLR, D(10)=>OutputImg4_42_EXMPLR, D(9)=>
      OutputImg4_41_EXMPLR, D(8)=>OutputImg4_40_EXMPLR, D(7)=>
      OutputImg4_39_EXMPLR, D(6)=>OutputImg4_38_EXMPLR, D(5)=>
      OutputImg4_37_EXMPLR, D(4)=>OutputImg4_36_EXMPLR, D(3)=>
      OutputImg4_35_EXMPLR, D(2)=>OutputImg4_34_EXMPLR, D(1)=>
      OutputImg4_33_EXMPLR, D(0)=>OutputImg4_32_EXMPLR, EN=>nx23668, F(15)=>
      ImgReg4IN_31, F(14)=>ImgReg4IN_30, F(13)=>ImgReg4IN_29, F(12)=>
      ImgReg4IN_28, F(11)=>ImgReg4IN_27, F(10)=>ImgReg4IN_26, F(9)=>
      ImgReg4IN_25, F(8)=>ImgReg4IN_24, F(7)=>ImgReg4IN_23, F(6)=>
      ImgReg4IN_22, F(5)=>ImgReg4IN_21, F(4)=>ImgReg4IN_20, F(3)=>
      ImgReg4IN_19, F(2)=>ImgReg4IN_18, F(1)=>ImgReg4IN_17, F(0)=>
      ImgReg4IN_16);
   loop3_1_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_47_EXMPLR, D(14)=>OutputImg5_46_EXMPLR, D(13)=>
      OutputImg5_45_EXMPLR, D(12)=>OutputImg5_44_EXMPLR, D(11)=>
      OutputImg5_43_EXMPLR, D(10)=>OutputImg5_42_EXMPLR, D(9)=>
      OutputImg5_41_EXMPLR, D(8)=>OutputImg5_40_EXMPLR, D(7)=>
      OutputImg5_39_EXMPLR, D(6)=>OutputImg5_38_EXMPLR, D(5)=>
      OutputImg5_37_EXMPLR, D(4)=>OutputImg5_36_EXMPLR, D(3)=>
      OutputImg5_35_EXMPLR, D(2)=>OutputImg5_34_EXMPLR, D(1)=>
      OutputImg5_33_EXMPLR, D(0)=>OutputImg5_32_EXMPLR, EN=>nx23668, F(15)=>
      ImgReg5IN_31, F(14)=>ImgReg5IN_30, F(13)=>ImgReg5IN_29, F(12)=>
      ImgReg5IN_28, F(11)=>ImgReg5IN_27, F(10)=>ImgReg5IN_26, F(9)=>
      ImgReg5IN_25, F(8)=>ImgReg5IN_24, F(7)=>ImgReg5IN_23, F(6)=>
      ImgReg5IN_22, F(5)=>ImgReg5IN_21, F(4)=>ImgReg5IN_20, F(3)=>
      ImgReg5IN_19, F(2)=>ImgReg5IN_18, F(1)=>ImgReg5IN_17, F(0)=>
      ImgReg5IN_16);
   loop3_1_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(31), D(14)
      =>DATA(30), D(13)=>DATA(29), D(12)=>DATA(28), D(11)=>DATA(27), D(10)=>
      DATA(26), D(9)=>DATA(25), D(8)=>DATA(24), D(7)=>DATA(23), D(6)=>
      DATA(22), D(5)=>DATA(21), D(4)=>DATA(20), D(3)=>DATA(19), D(2)=>
      DATA(18), D(1)=>DATA(17), D(0)=>DATA(16), EN=>nx23654, F(15)=>
      ImgReg0IN_31, F(14)=>ImgReg0IN_30, F(13)=>ImgReg0IN_29, F(12)=>
      ImgReg0IN_28, F(11)=>ImgReg0IN_27, F(10)=>ImgReg0IN_26, F(9)=>
      ImgReg0IN_25, F(8)=>ImgReg0IN_24, F(7)=>ImgReg0IN_23, F(6)=>
      ImgReg0IN_22, F(5)=>ImgReg0IN_21, F(4)=>ImgReg0IN_20, F(3)=>
      ImgReg0IN_19, F(2)=>ImgReg0IN_18, F(1)=>ImgReg0IN_17, F(0)=>
      ImgReg0IN_16);
   loop3_1_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(31), D(14)
      =>DATA(30), D(13)=>DATA(29), D(12)=>DATA(28), D(11)=>DATA(27), D(10)=>
      DATA(26), D(9)=>DATA(25), D(8)=>DATA(24), D(7)=>DATA(23), D(6)=>
      DATA(22), D(5)=>DATA(21), D(4)=>DATA(20), D(3)=>DATA(19), D(2)=>
      DATA(18), D(1)=>DATA(17), D(0)=>DATA(16), EN=>nx23642, F(15)=>
      ImgReg1IN_31, F(14)=>ImgReg1IN_30, F(13)=>ImgReg1IN_29, F(12)=>
      ImgReg1IN_28, F(11)=>ImgReg1IN_27, F(10)=>ImgReg1IN_26, F(9)=>
      ImgReg1IN_25, F(8)=>ImgReg1IN_24, F(7)=>ImgReg1IN_23, F(6)=>
      ImgReg1IN_22, F(5)=>ImgReg1IN_21, F(4)=>ImgReg1IN_20, F(3)=>
      ImgReg1IN_19, F(2)=>ImgReg1IN_18, F(1)=>ImgReg1IN_17, F(0)=>
      ImgReg1IN_16);
   loop3_1_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(31), D(14)
      =>DATA(30), D(13)=>DATA(29), D(12)=>DATA(28), D(11)=>DATA(27), D(10)=>
      DATA(26), D(9)=>DATA(25), D(8)=>DATA(24), D(7)=>DATA(23), D(6)=>
      DATA(22), D(5)=>DATA(21), D(4)=>DATA(20), D(3)=>DATA(19), D(2)=>
      DATA(18), D(1)=>DATA(17), D(0)=>DATA(16), EN=>nx23630, F(15)=>
      ImgReg2IN_31, F(14)=>ImgReg2IN_30, F(13)=>ImgReg2IN_29, F(12)=>
      ImgReg2IN_28, F(11)=>ImgReg2IN_27, F(10)=>ImgReg2IN_26, F(9)=>
      ImgReg2IN_25, F(8)=>ImgReg2IN_24, F(7)=>ImgReg2IN_23, F(6)=>
      ImgReg2IN_22, F(5)=>ImgReg2IN_21, F(4)=>ImgReg2IN_20, F(3)=>
      ImgReg2IN_19, F(2)=>ImgReg2IN_18, F(1)=>ImgReg2IN_17, F(0)=>
      ImgReg2IN_16);
   loop3_1_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(31), D(14)
      =>DATA(30), D(13)=>DATA(29), D(12)=>DATA(28), D(11)=>DATA(27), D(10)=>
      DATA(26), D(9)=>DATA(25), D(8)=>DATA(24), D(7)=>DATA(23), D(6)=>
      DATA(22), D(5)=>DATA(21), D(4)=>DATA(20), D(3)=>DATA(19), D(2)=>
      DATA(18), D(1)=>DATA(17), D(0)=>DATA(16), EN=>nx23618, F(15)=>
      ImgReg3IN_31, F(14)=>ImgReg3IN_30, F(13)=>ImgReg3IN_29, F(12)=>
      ImgReg3IN_28, F(11)=>ImgReg3IN_27, F(10)=>ImgReg3IN_26, F(9)=>
      ImgReg3IN_25, F(8)=>ImgReg3IN_24, F(7)=>ImgReg3IN_23, F(6)=>
      ImgReg3IN_22, F(5)=>ImgReg3IN_21, F(4)=>ImgReg3IN_20, F(3)=>
      ImgReg3IN_19, F(2)=>ImgReg3IN_18, F(1)=>ImgReg3IN_17, F(0)=>
      ImgReg3IN_16);
   loop3_1_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(31), D(14)
      =>DATA(30), D(13)=>DATA(29), D(12)=>DATA(28), D(11)=>DATA(27), D(10)=>
      DATA(26), D(9)=>DATA(25), D(8)=>DATA(24), D(7)=>DATA(23), D(6)=>
      DATA(22), D(5)=>DATA(21), D(4)=>DATA(20), D(3)=>DATA(19), D(2)=>
      DATA(18), D(1)=>DATA(17), D(0)=>DATA(16), EN=>nx23606, F(15)=>
      ImgReg4IN_31, F(14)=>ImgReg4IN_30, F(13)=>ImgReg4IN_29, F(12)=>
      ImgReg4IN_28, F(11)=>ImgReg4IN_27, F(10)=>ImgReg4IN_26, F(9)=>
      ImgReg4IN_25, F(8)=>ImgReg4IN_24, F(7)=>ImgReg4IN_23, F(6)=>
      ImgReg4IN_22, F(5)=>ImgReg4IN_21, F(4)=>ImgReg4IN_20, F(3)=>
      ImgReg4IN_19, F(2)=>ImgReg4IN_18, F(1)=>ImgReg4IN_17, F(0)=>
      ImgReg4IN_16);
   loop3_1_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(31), D(14)
      =>DATA(30), D(13)=>DATA(29), D(12)=>DATA(28), D(11)=>DATA(27), D(10)=>
      DATA(26), D(9)=>DATA(25), D(8)=>DATA(24), D(7)=>DATA(23), D(6)=>
      DATA(22), D(5)=>DATA(21), D(4)=>DATA(20), D(3)=>DATA(19), D(2)=>
      DATA(18), D(1)=>DATA(17), D(0)=>DATA(16), EN=>nx23594, F(15)=>
      ImgReg5IN_31, F(14)=>ImgReg5IN_30, F(13)=>ImgReg5IN_29, F(12)=>
      ImgReg5IN_28, F(11)=>ImgReg5IN_27, F(10)=>ImgReg5IN_26, F(9)=>
      ImgReg5IN_25, F(8)=>ImgReg5IN_24, F(7)=>ImgReg5IN_23, F(6)=>
      ImgReg5IN_22, F(5)=>ImgReg5IN_21, F(4)=>ImgReg5IN_20, F(3)=>
      ImgReg5IN_19, F(2)=>ImgReg5IN_18, F(1)=>ImgReg5IN_17, F(0)=>
      ImgReg5IN_16);
   loop3_1_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_31_EXMPLR, D(14)=>OutputImg1_30_EXMPLR, D(13)=>
      OutputImg1_29_EXMPLR, D(12)=>OutputImg1_28_EXMPLR, D(11)=>
      OutputImg1_27_EXMPLR, D(10)=>OutputImg1_26_EXMPLR, D(9)=>
      OutputImg1_25_EXMPLR, D(8)=>OutputImg1_24_EXMPLR, D(7)=>
      OutputImg1_23_EXMPLR, D(6)=>OutputImg1_22_EXMPLR, D(5)=>
      OutputImg1_21_EXMPLR, D(4)=>OutputImg1_20_EXMPLR, D(3)=>
      OutputImg1_19_EXMPLR, D(2)=>OutputImg1_18_EXMPLR, D(1)=>
      OutputImg1_17_EXMPLR, D(0)=>OutputImg1_16_EXMPLR, EN=>nx23786, F(15)=>
      ImgReg0IN_31, F(14)=>ImgReg0IN_30, F(13)=>ImgReg0IN_29, F(12)=>
      ImgReg0IN_28, F(11)=>ImgReg0IN_27, F(10)=>ImgReg0IN_26, F(9)=>
      ImgReg0IN_25, F(8)=>ImgReg0IN_24, F(7)=>ImgReg0IN_23, F(6)=>
      ImgReg0IN_22, F(5)=>ImgReg0IN_21, F(4)=>ImgReg0IN_20, F(3)=>
      ImgReg0IN_19, F(2)=>ImgReg0IN_18, F(1)=>ImgReg0IN_17, F(0)=>
      ImgReg0IN_16);
   loop3_1_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_31_EXMPLR, D(14)=>OutputImg2_30_EXMPLR, D(13)=>
      OutputImg2_29_EXMPLR, D(12)=>OutputImg2_28_EXMPLR, D(11)=>
      OutputImg2_27_EXMPLR, D(10)=>OutputImg2_26_EXMPLR, D(9)=>
      OutputImg2_25_EXMPLR, D(8)=>OutputImg2_24_EXMPLR, D(7)=>
      OutputImg2_23_EXMPLR, D(6)=>OutputImg2_22_EXMPLR, D(5)=>
      OutputImg2_21_EXMPLR, D(4)=>OutputImg2_20_EXMPLR, D(3)=>
      OutputImg2_19_EXMPLR, D(2)=>OutputImg2_18_EXMPLR, D(1)=>
      OutputImg2_17_EXMPLR, D(0)=>OutputImg2_16_EXMPLR, EN=>nx23786, F(15)=>
      ImgReg1IN_31, F(14)=>ImgReg1IN_30, F(13)=>ImgReg1IN_29, F(12)=>
      ImgReg1IN_28, F(11)=>ImgReg1IN_27, F(10)=>ImgReg1IN_26, F(9)=>
      ImgReg1IN_25, F(8)=>ImgReg1IN_24, F(7)=>ImgReg1IN_23, F(6)=>
      ImgReg1IN_22, F(5)=>ImgReg1IN_21, F(4)=>ImgReg1IN_20, F(3)=>
      ImgReg1IN_19, F(2)=>ImgReg1IN_18, F(1)=>ImgReg1IN_17, F(0)=>
      ImgReg1IN_16);
   loop3_1_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_31_EXMPLR, D(14)=>OutputImg3_30_EXMPLR, D(13)=>
      OutputImg3_29_EXMPLR, D(12)=>OutputImg3_28_EXMPLR, D(11)=>
      OutputImg3_27_EXMPLR, D(10)=>OutputImg3_26_EXMPLR, D(9)=>
      OutputImg3_25_EXMPLR, D(8)=>OutputImg3_24_EXMPLR, D(7)=>
      OutputImg3_23_EXMPLR, D(6)=>OutputImg3_22_EXMPLR, D(5)=>
      OutputImg3_21_EXMPLR, D(4)=>OutputImg3_20_EXMPLR, D(3)=>
      OutputImg3_19_EXMPLR, D(2)=>OutputImg3_18_EXMPLR, D(1)=>
      OutputImg3_17_EXMPLR, D(0)=>OutputImg3_16_EXMPLR, EN=>nx23788, F(15)=>
      ImgReg2IN_31, F(14)=>ImgReg2IN_30, F(13)=>ImgReg2IN_29, F(12)=>
      ImgReg2IN_28, F(11)=>ImgReg2IN_27, F(10)=>ImgReg2IN_26, F(9)=>
      ImgReg2IN_25, F(8)=>ImgReg2IN_24, F(7)=>ImgReg2IN_23, F(6)=>
      ImgReg2IN_22, F(5)=>ImgReg2IN_21, F(4)=>ImgReg2IN_20, F(3)=>
      ImgReg2IN_19, F(2)=>ImgReg2IN_18, F(1)=>ImgReg2IN_17, F(0)=>
      ImgReg2IN_16);
   loop3_1_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_31_EXMPLR, D(14)=>OutputImg4_30_EXMPLR, D(13)=>
      OutputImg4_29_EXMPLR, D(12)=>OutputImg4_28_EXMPLR, D(11)=>
      OutputImg4_27_EXMPLR, D(10)=>OutputImg4_26_EXMPLR, D(9)=>
      OutputImg4_25_EXMPLR, D(8)=>OutputImg4_24_EXMPLR, D(7)=>
      OutputImg4_23_EXMPLR, D(6)=>OutputImg4_22_EXMPLR, D(5)=>
      OutputImg4_21_EXMPLR, D(4)=>OutputImg4_20_EXMPLR, D(3)=>
      OutputImg4_19_EXMPLR, D(2)=>OutputImg4_18_EXMPLR, D(1)=>
      OutputImg4_17_EXMPLR, D(0)=>OutputImg4_16_EXMPLR, EN=>nx23788, F(15)=>
      ImgReg3IN_31, F(14)=>ImgReg3IN_30, F(13)=>ImgReg3IN_29, F(12)=>
      ImgReg3IN_28, F(11)=>ImgReg3IN_27, F(10)=>ImgReg3IN_26, F(9)=>
      ImgReg3IN_25, F(8)=>ImgReg3IN_24, F(7)=>ImgReg3IN_23, F(6)=>
      ImgReg3IN_22, F(5)=>ImgReg3IN_21, F(4)=>ImgReg3IN_20, F(3)=>
      ImgReg3IN_19, F(2)=>ImgReg3IN_18, F(1)=>ImgReg3IN_17, F(0)=>
      ImgReg3IN_16);
   loop3_1_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_31_EXMPLR, D(14)=>OutputImg5_30_EXMPLR, D(13)=>
      OutputImg5_29_EXMPLR, D(12)=>OutputImg5_28_EXMPLR, D(11)=>
      OutputImg5_27_EXMPLR, D(10)=>OutputImg5_26_EXMPLR, D(9)=>
      OutputImg5_25_EXMPLR, D(8)=>OutputImg5_24_EXMPLR, D(7)=>
      OutputImg5_23_EXMPLR, D(6)=>OutputImg5_22_EXMPLR, D(5)=>
      OutputImg5_21_EXMPLR, D(4)=>OutputImg5_20_EXMPLR, D(3)=>
      OutputImg5_19_EXMPLR, D(2)=>OutputImg5_18_EXMPLR, D(1)=>
      OutputImg5_17_EXMPLR, D(0)=>OutputImg5_16_EXMPLR, EN=>nx23788, F(15)=>
      ImgReg4IN_31, F(14)=>ImgReg4IN_30, F(13)=>ImgReg4IN_29, F(12)=>
      ImgReg4IN_28, F(11)=>ImgReg4IN_27, F(10)=>ImgReg4IN_26, F(9)=>
      ImgReg4IN_25, F(8)=>ImgReg4IN_24, F(7)=>ImgReg4IN_23, F(6)=>
      ImgReg4IN_22, F(5)=>ImgReg4IN_21, F(4)=>ImgReg4IN_20, F(3)=>
      ImgReg4IN_19, F(2)=>ImgReg4IN_18, F(1)=>ImgReg4IN_17, F(0)=>
      ImgReg4IN_16);
   loop3_1_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_31, D(14)=>
      ImgReg0IN_30, D(13)=>ImgReg0IN_29, D(12)=>ImgReg0IN_28, D(11)=>
      ImgReg0IN_27, D(10)=>ImgReg0IN_26, D(9)=>ImgReg0IN_25, D(8)=>
      ImgReg0IN_24, D(7)=>ImgReg0IN_23, D(6)=>ImgReg0IN_22, D(5)=>
      ImgReg0IN_21, D(4)=>ImgReg0IN_20, D(3)=>ImgReg0IN_19, D(2)=>
      ImgReg0IN_18, D(1)=>ImgReg0IN_17, D(0)=>ImgReg0IN_16, CLK=>nx23834, 
      RST=>RST, EN=>nx23718, Q(15)=>OutputImg0_31_EXMPLR, Q(14)=>
      OutputImg0_30_EXMPLR, Q(13)=>OutputImg0_29_EXMPLR, Q(12)=>
      OutputImg0_28_EXMPLR, Q(11)=>OutputImg0_27_EXMPLR, Q(10)=>
      OutputImg0_26_EXMPLR, Q(9)=>OutputImg0_25_EXMPLR, Q(8)=>
      OutputImg0_24_EXMPLR, Q(7)=>OutputImg0_23_EXMPLR, Q(6)=>
      OutputImg0_22_EXMPLR, Q(5)=>OutputImg0_21_EXMPLR, Q(4)=>
      OutputImg0_20_EXMPLR, Q(3)=>OutputImg0_19_EXMPLR, Q(2)=>
      OutputImg0_18_EXMPLR, Q(1)=>OutputImg0_17_EXMPLR, Q(0)=>
      OutputImg0_16_EXMPLR);
   loop3_1_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_31, D(14)=>
      ImgReg1IN_30, D(13)=>ImgReg1IN_29, D(12)=>ImgReg1IN_28, D(11)=>
      ImgReg1IN_27, D(10)=>ImgReg1IN_26, D(9)=>ImgReg1IN_25, D(8)=>
      ImgReg1IN_24, D(7)=>ImgReg1IN_23, D(6)=>ImgReg1IN_22, D(5)=>
      ImgReg1IN_21, D(4)=>ImgReg1IN_20, D(3)=>ImgReg1IN_19, D(2)=>
      ImgReg1IN_18, D(1)=>ImgReg1IN_17, D(0)=>ImgReg1IN_16, CLK=>nx23836, 
      RST=>RST, EN=>nx23728, Q(15)=>OutputImg1_31_EXMPLR, Q(14)=>
      OutputImg1_30_EXMPLR, Q(13)=>OutputImg1_29_EXMPLR, Q(12)=>
      OutputImg1_28_EXMPLR, Q(11)=>OutputImg1_27_EXMPLR, Q(10)=>
      OutputImg1_26_EXMPLR, Q(9)=>OutputImg1_25_EXMPLR, Q(8)=>
      OutputImg1_24_EXMPLR, Q(7)=>OutputImg1_23_EXMPLR, Q(6)=>
      OutputImg1_22_EXMPLR, Q(5)=>OutputImg1_21_EXMPLR, Q(4)=>
      OutputImg1_20_EXMPLR, Q(3)=>OutputImg1_19_EXMPLR, Q(2)=>
      OutputImg1_18_EXMPLR, Q(1)=>OutputImg1_17_EXMPLR, Q(0)=>
      OutputImg1_16_EXMPLR);
   loop3_1_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_31, D(14)=>
      ImgReg2IN_30, D(13)=>ImgReg2IN_29, D(12)=>ImgReg2IN_28, D(11)=>
      ImgReg2IN_27, D(10)=>ImgReg2IN_26, D(9)=>ImgReg2IN_25, D(8)=>
      ImgReg2IN_24, D(7)=>ImgReg2IN_23, D(6)=>ImgReg2IN_22, D(5)=>
      ImgReg2IN_21, D(4)=>ImgReg2IN_20, D(3)=>ImgReg2IN_19, D(2)=>
      ImgReg2IN_18, D(1)=>ImgReg2IN_17, D(0)=>ImgReg2IN_16, CLK=>nx23836, 
      RST=>RST, EN=>nx23738, Q(15)=>OutputImg2_31_EXMPLR, Q(14)=>
      OutputImg2_30_EXMPLR, Q(13)=>OutputImg2_29_EXMPLR, Q(12)=>
      OutputImg2_28_EXMPLR, Q(11)=>OutputImg2_27_EXMPLR, Q(10)=>
      OutputImg2_26_EXMPLR, Q(9)=>OutputImg2_25_EXMPLR, Q(8)=>
      OutputImg2_24_EXMPLR, Q(7)=>OutputImg2_23_EXMPLR, Q(6)=>
      OutputImg2_22_EXMPLR, Q(5)=>OutputImg2_21_EXMPLR, Q(4)=>
      OutputImg2_20_EXMPLR, Q(3)=>OutputImg2_19_EXMPLR, Q(2)=>
      OutputImg2_18_EXMPLR, Q(1)=>OutputImg2_17_EXMPLR, Q(0)=>
      OutputImg2_16_EXMPLR);
   loop3_1_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_31, D(14)=>
      ImgReg3IN_30, D(13)=>ImgReg3IN_29, D(12)=>ImgReg3IN_28, D(11)=>
      ImgReg3IN_27, D(10)=>ImgReg3IN_26, D(9)=>ImgReg3IN_25, D(8)=>
      ImgReg3IN_24, D(7)=>ImgReg3IN_23, D(6)=>ImgReg3IN_22, D(5)=>
      ImgReg3IN_21, D(4)=>ImgReg3IN_20, D(3)=>ImgReg3IN_19, D(2)=>
      ImgReg3IN_18, D(1)=>ImgReg3IN_17, D(0)=>ImgReg3IN_16, CLK=>nx23838, 
      RST=>RST, EN=>nx23748, Q(15)=>OutputImg3_31_EXMPLR, Q(14)=>
      OutputImg3_30_EXMPLR, Q(13)=>OutputImg3_29_EXMPLR, Q(12)=>
      OutputImg3_28_EXMPLR, Q(11)=>OutputImg3_27_EXMPLR, Q(10)=>
      OutputImg3_26_EXMPLR, Q(9)=>OutputImg3_25_EXMPLR, Q(8)=>
      OutputImg3_24_EXMPLR, Q(7)=>OutputImg3_23_EXMPLR, Q(6)=>
      OutputImg3_22_EXMPLR, Q(5)=>OutputImg3_21_EXMPLR, Q(4)=>
      OutputImg3_20_EXMPLR, Q(3)=>OutputImg3_19_EXMPLR, Q(2)=>
      OutputImg3_18_EXMPLR, Q(1)=>OutputImg3_17_EXMPLR, Q(0)=>
      OutputImg3_16_EXMPLR);
   loop3_1_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_31, D(14)=>
      ImgReg4IN_30, D(13)=>ImgReg4IN_29, D(12)=>ImgReg4IN_28, D(11)=>
      ImgReg4IN_27, D(10)=>ImgReg4IN_26, D(9)=>ImgReg4IN_25, D(8)=>
      ImgReg4IN_24, D(7)=>ImgReg4IN_23, D(6)=>ImgReg4IN_22, D(5)=>
      ImgReg4IN_21, D(4)=>ImgReg4IN_20, D(3)=>ImgReg4IN_19, D(2)=>
      ImgReg4IN_18, D(1)=>ImgReg4IN_17, D(0)=>ImgReg4IN_16, CLK=>nx23838, 
      RST=>RST, EN=>nx23758, Q(15)=>OutputImg4_31_EXMPLR, Q(14)=>
      OutputImg4_30_EXMPLR, Q(13)=>OutputImg4_29_EXMPLR, Q(12)=>
      OutputImg4_28_EXMPLR, Q(11)=>OutputImg4_27_EXMPLR, Q(10)=>
      OutputImg4_26_EXMPLR, Q(9)=>OutputImg4_25_EXMPLR, Q(8)=>
      OutputImg4_24_EXMPLR, Q(7)=>OutputImg4_23_EXMPLR, Q(6)=>
      OutputImg4_22_EXMPLR, Q(5)=>OutputImg4_21_EXMPLR, Q(4)=>
      OutputImg4_20_EXMPLR, Q(3)=>OutputImg4_19_EXMPLR, Q(2)=>
      OutputImg4_18_EXMPLR, Q(1)=>OutputImg4_17_EXMPLR, Q(0)=>
      OutputImg4_16_EXMPLR);
   loop3_1_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_31, D(14)=>
      ImgReg5IN_30, D(13)=>ImgReg5IN_29, D(12)=>ImgReg5IN_28, D(11)=>
      ImgReg5IN_27, D(10)=>ImgReg5IN_26, D(9)=>ImgReg5IN_25, D(8)=>
      ImgReg5IN_24, D(7)=>ImgReg5IN_23, D(6)=>ImgReg5IN_22, D(5)=>
      ImgReg5IN_21, D(4)=>ImgReg5IN_20, D(3)=>ImgReg5IN_19, D(2)=>
      ImgReg5IN_18, D(1)=>ImgReg5IN_17, D(0)=>ImgReg5IN_16, CLK=>nx23840, 
      RST=>RST, EN=>nx23768, Q(15)=>OutputImg5_31_EXMPLR, Q(14)=>
      OutputImg5_30_EXMPLR, Q(13)=>OutputImg5_29_EXMPLR, Q(12)=>
      OutputImg5_28_EXMPLR, Q(11)=>OutputImg5_27_EXMPLR, Q(10)=>
      OutputImg5_26_EXMPLR, Q(9)=>OutputImg5_25_EXMPLR, Q(8)=>
      OutputImg5_24_EXMPLR, Q(7)=>OutputImg5_23_EXMPLR, Q(6)=>
      OutputImg5_22_EXMPLR, Q(5)=>OutputImg5_21_EXMPLR, Q(4)=>
      OutputImg5_20_EXMPLR, Q(3)=>OutputImg5_19_EXMPLR, Q(2)=>
      OutputImg5_18_EXMPLR, Q(1)=>OutputImg5_17_EXMPLR, Q(0)=>
      OutputImg5_16_EXMPLR);
   loop3_2_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_63_EXMPLR, D(14)=>OutputImg0_62_EXMPLR, D(13)=>
      OutputImg0_61_EXMPLR, D(12)=>OutputImg0_60_EXMPLR, D(11)=>
      OutputImg0_59_EXMPLR, D(10)=>OutputImg0_58_EXMPLR, D(9)=>
      OutputImg0_57_EXMPLR, D(8)=>OutputImg0_56_EXMPLR, D(7)=>
      OutputImg0_55_EXMPLR, D(6)=>OutputImg0_54_EXMPLR, D(5)=>
      OutputImg0_53_EXMPLR, D(4)=>OutputImg0_52_EXMPLR, D(3)=>
      OutputImg0_51_EXMPLR, D(2)=>OutputImg0_50_EXMPLR, D(1)=>
      OutputImg0_49_EXMPLR, D(0)=>OutputImg0_48_EXMPLR, EN=>nx23668, F(15)=>
      ImgReg0IN_47, F(14)=>ImgReg0IN_46, F(13)=>ImgReg0IN_45, F(12)=>
      ImgReg0IN_44, F(11)=>ImgReg0IN_43, F(10)=>ImgReg0IN_42, F(9)=>
      ImgReg0IN_41, F(8)=>ImgReg0IN_40, F(7)=>ImgReg0IN_39, F(6)=>
      ImgReg0IN_38, F(5)=>ImgReg0IN_37, F(4)=>ImgReg0IN_36, F(3)=>
      ImgReg0IN_35, F(2)=>ImgReg0IN_34, F(1)=>ImgReg0IN_33, F(0)=>
      ImgReg0IN_32);
   loop3_2_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_63_EXMPLR, D(14)=>OutputImg1_62_EXMPLR, D(13)=>
      OutputImg1_61_EXMPLR, D(12)=>OutputImg1_60_EXMPLR, D(11)=>
      OutputImg1_59_EXMPLR, D(10)=>OutputImg1_58_EXMPLR, D(9)=>
      OutputImg1_57_EXMPLR, D(8)=>OutputImg1_56_EXMPLR, D(7)=>
      OutputImg1_55_EXMPLR, D(6)=>OutputImg1_54_EXMPLR, D(5)=>
      OutputImg1_53_EXMPLR, D(4)=>OutputImg1_52_EXMPLR, D(3)=>
      OutputImg1_51_EXMPLR, D(2)=>OutputImg1_50_EXMPLR, D(1)=>
      OutputImg1_49_EXMPLR, D(0)=>OutputImg1_48_EXMPLR, EN=>nx23668, F(15)=>
      ImgReg1IN_47, F(14)=>ImgReg1IN_46, F(13)=>ImgReg1IN_45, F(12)=>
      ImgReg1IN_44, F(11)=>ImgReg1IN_43, F(10)=>ImgReg1IN_42, F(9)=>
      ImgReg1IN_41, F(8)=>ImgReg1IN_40, F(7)=>ImgReg1IN_39, F(6)=>
      ImgReg1IN_38, F(5)=>ImgReg1IN_37, F(4)=>ImgReg1IN_36, F(3)=>
      ImgReg1IN_35, F(2)=>ImgReg1IN_34, F(1)=>ImgReg1IN_33, F(0)=>
      ImgReg1IN_32);
   loop3_2_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_63_EXMPLR, D(14)=>OutputImg2_62_EXMPLR, D(13)=>
      OutputImg2_61_EXMPLR, D(12)=>OutputImg2_60_EXMPLR, D(11)=>
      OutputImg2_59_EXMPLR, D(10)=>OutputImg2_58_EXMPLR, D(9)=>
      OutputImg2_57_EXMPLR, D(8)=>OutputImg2_56_EXMPLR, D(7)=>
      OutputImg2_55_EXMPLR, D(6)=>OutputImg2_54_EXMPLR, D(5)=>
      OutputImg2_53_EXMPLR, D(4)=>OutputImg2_52_EXMPLR, D(3)=>
      OutputImg2_51_EXMPLR, D(2)=>OutputImg2_50_EXMPLR, D(1)=>
      OutputImg2_49_EXMPLR, D(0)=>OutputImg2_48_EXMPLR, EN=>nx23670, F(15)=>
      ImgReg2IN_47, F(14)=>ImgReg2IN_46, F(13)=>ImgReg2IN_45, F(12)=>
      ImgReg2IN_44, F(11)=>ImgReg2IN_43, F(10)=>ImgReg2IN_42, F(9)=>
      ImgReg2IN_41, F(8)=>ImgReg2IN_40, F(7)=>ImgReg2IN_39, F(6)=>
      ImgReg2IN_38, F(5)=>ImgReg2IN_37, F(4)=>ImgReg2IN_36, F(3)=>
      ImgReg2IN_35, F(2)=>ImgReg2IN_34, F(1)=>ImgReg2IN_33, F(0)=>
      ImgReg2IN_32);
   loop3_2_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_63_EXMPLR, D(14)=>OutputImg3_62_EXMPLR, D(13)=>
      OutputImg3_61_EXMPLR, D(12)=>OutputImg3_60_EXMPLR, D(11)=>
      OutputImg3_59_EXMPLR, D(10)=>OutputImg3_58_EXMPLR, D(9)=>
      OutputImg3_57_EXMPLR, D(8)=>OutputImg3_56_EXMPLR, D(7)=>
      OutputImg3_55_EXMPLR, D(6)=>OutputImg3_54_EXMPLR, D(5)=>
      OutputImg3_53_EXMPLR, D(4)=>OutputImg3_52_EXMPLR, D(3)=>
      OutputImg3_51_EXMPLR, D(2)=>OutputImg3_50_EXMPLR, D(1)=>
      OutputImg3_49_EXMPLR, D(0)=>OutputImg3_48_EXMPLR, EN=>nx23670, F(15)=>
      ImgReg3IN_47, F(14)=>ImgReg3IN_46, F(13)=>ImgReg3IN_45, F(12)=>
      ImgReg3IN_44, F(11)=>ImgReg3IN_43, F(10)=>ImgReg3IN_42, F(9)=>
      ImgReg3IN_41, F(8)=>ImgReg3IN_40, F(7)=>ImgReg3IN_39, F(6)=>
      ImgReg3IN_38, F(5)=>ImgReg3IN_37, F(4)=>ImgReg3IN_36, F(3)=>
      ImgReg3IN_35, F(2)=>ImgReg3IN_34, F(1)=>ImgReg3IN_33, F(0)=>
      ImgReg3IN_32);
   loop3_2_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_63_EXMPLR, D(14)=>OutputImg4_62_EXMPLR, D(13)=>
      OutputImg4_61_EXMPLR, D(12)=>OutputImg4_60_EXMPLR, D(11)=>
      OutputImg4_59_EXMPLR, D(10)=>OutputImg4_58_EXMPLR, D(9)=>
      OutputImg4_57_EXMPLR, D(8)=>OutputImg4_56_EXMPLR, D(7)=>
      OutputImg4_55_EXMPLR, D(6)=>OutputImg4_54_EXMPLR, D(5)=>
      OutputImg4_53_EXMPLR, D(4)=>OutputImg4_52_EXMPLR, D(3)=>
      OutputImg4_51_EXMPLR, D(2)=>OutputImg4_50_EXMPLR, D(1)=>
      OutputImg4_49_EXMPLR, D(0)=>OutputImg4_48_EXMPLR, EN=>nx23670, F(15)=>
      ImgReg4IN_47, F(14)=>ImgReg4IN_46, F(13)=>ImgReg4IN_45, F(12)=>
      ImgReg4IN_44, F(11)=>ImgReg4IN_43, F(10)=>ImgReg4IN_42, F(9)=>
      ImgReg4IN_41, F(8)=>ImgReg4IN_40, F(7)=>ImgReg4IN_39, F(6)=>
      ImgReg4IN_38, F(5)=>ImgReg4IN_37, F(4)=>ImgReg4IN_36, F(3)=>
      ImgReg4IN_35, F(2)=>ImgReg4IN_34, F(1)=>ImgReg4IN_33, F(0)=>
      ImgReg4IN_32);
   loop3_2_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_63_EXMPLR, D(14)=>OutputImg5_62_EXMPLR, D(13)=>
      OutputImg5_61_EXMPLR, D(12)=>OutputImg5_60_EXMPLR, D(11)=>
      OutputImg5_59_EXMPLR, D(10)=>OutputImg5_58_EXMPLR, D(9)=>
      OutputImg5_57_EXMPLR, D(8)=>OutputImg5_56_EXMPLR, D(7)=>
      OutputImg5_55_EXMPLR, D(6)=>OutputImg5_54_EXMPLR, D(5)=>
      OutputImg5_53_EXMPLR, D(4)=>OutputImg5_52_EXMPLR, D(3)=>
      OutputImg5_51_EXMPLR, D(2)=>OutputImg5_50_EXMPLR, D(1)=>
      OutputImg5_49_EXMPLR, D(0)=>OutputImg5_48_EXMPLR, EN=>nx23670, F(15)=>
      ImgReg5IN_47, F(14)=>ImgReg5IN_46, F(13)=>ImgReg5IN_45, F(12)=>
      ImgReg5IN_44, F(11)=>ImgReg5IN_43, F(10)=>ImgReg5IN_42, F(9)=>
      ImgReg5IN_41, F(8)=>ImgReg5IN_40, F(7)=>ImgReg5IN_39, F(6)=>
      ImgReg5IN_38, F(5)=>ImgReg5IN_37, F(4)=>ImgReg5IN_36, F(3)=>
      ImgReg5IN_35, F(2)=>ImgReg5IN_34, F(1)=>ImgReg5IN_33, F(0)=>
      ImgReg5IN_32);
   loop3_2_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(47), D(14)
      =>DATA(46), D(13)=>DATA(45), D(12)=>DATA(44), D(11)=>DATA(43), D(10)=>
      DATA(42), D(9)=>DATA(41), D(8)=>DATA(40), D(7)=>DATA(39), D(6)=>
      DATA(38), D(5)=>DATA(37), D(4)=>DATA(36), D(3)=>DATA(35), D(2)=>
      DATA(34), D(1)=>DATA(33), D(0)=>DATA(32), EN=>nx23654, F(15)=>
      ImgReg0IN_47, F(14)=>ImgReg0IN_46, F(13)=>ImgReg0IN_45, F(12)=>
      ImgReg0IN_44, F(11)=>ImgReg0IN_43, F(10)=>ImgReg0IN_42, F(9)=>
      ImgReg0IN_41, F(8)=>ImgReg0IN_40, F(7)=>ImgReg0IN_39, F(6)=>
      ImgReg0IN_38, F(5)=>ImgReg0IN_37, F(4)=>ImgReg0IN_36, F(3)=>
      ImgReg0IN_35, F(2)=>ImgReg0IN_34, F(1)=>ImgReg0IN_33, F(0)=>
      ImgReg0IN_32);
   loop3_2_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(47), D(14)
      =>DATA(46), D(13)=>DATA(45), D(12)=>DATA(44), D(11)=>DATA(43), D(10)=>
      DATA(42), D(9)=>DATA(41), D(8)=>DATA(40), D(7)=>DATA(39), D(6)=>
      DATA(38), D(5)=>DATA(37), D(4)=>DATA(36), D(3)=>DATA(35), D(2)=>
      DATA(34), D(1)=>DATA(33), D(0)=>DATA(32), EN=>nx23642, F(15)=>
      ImgReg1IN_47, F(14)=>ImgReg1IN_46, F(13)=>ImgReg1IN_45, F(12)=>
      ImgReg1IN_44, F(11)=>ImgReg1IN_43, F(10)=>ImgReg1IN_42, F(9)=>
      ImgReg1IN_41, F(8)=>ImgReg1IN_40, F(7)=>ImgReg1IN_39, F(6)=>
      ImgReg1IN_38, F(5)=>ImgReg1IN_37, F(4)=>ImgReg1IN_36, F(3)=>
      ImgReg1IN_35, F(2)=>ImgReg1IN_34, F(1)=>ImgReg1IN_33, F(0)=>
      ImgReg1IN_32);
   loop3_2_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(47), D(14)
      =>DATA(46), D(13)=>DATA(45), D(12)=>DATA(44), D(11)=>DATA(43), D(10)=>
      DATA(42), D(9)=>DATA(41), D(8)=>DATA(40), D(7)=>DATA(39), D(6)=>
      DATA(38), D(5)=>DATA(37), D(4)=>DATA(36), D(3)=>DATA(35), D(2)=>
      DATA(34), D(1)=>DATA(33), D(0)=>DATA(32), EN=>nx23630, F(15)=>
      ImgReg2IN_47, F(14)=>ImgReg2IN_46, F(13)=>ImgReg2IN_45, F(12)=>
      ImgReg2IN_44, F(11)=>ImgReg2IN_43, F(10)=>ImgReg2IN_42, F(9)=>
      ImgReg2IN_41, F(8)=>ImgReg2IN_40, F(7)=>ImgReg2IN_39, F(6)=>
      ImgReg2IN_38, F(5)=>ImgReg2IN_37, F(4)=>ImgReg2IN_36, F(3)=>
      ImgReg2IN_35, F(2)=>ImgReg2IN_34, F(1)=>ImgReg2IN_33, F(0)=>
      ImgReg2IN_32);
   loop3_2_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(47), D(14)
      =>DATA(46), D(13)=>DATA(45), D(12)=>DATA(44), D(11)=>DATA(43), D(10)=>
      DATA(42), D(9)=>DATA(41), D(8)=>DATA(40), D(7)=>DATA(39), D(6)=>
      DATA(38), D(5)=>DATA(37), D(4)=>DATA(36), D(3)=>DATA(35), D(2)=>
      DATA(34), D(1)=>DATA(33), D(0)=>DATA(32), EN=>nx23618, F(15)=>
      ImgReg3IN_47, F(14)=>ImgReg3IN_46, F(13)=>ImgReg3IN_45, F(12)=>
      ImgReg3IN_44, F(11)=>ImgReg3IN_43, F(10)=>ImgReg3IN_42, F(9)=>
      ImgReg3IN_41, F(8)=>ImgReg3IN_40, F(7)=>ImgReg3IN_39, F(6)=>
      ImgReg3IN_38, F(5)=>ImgReg3IN_37, F(4)=>ImgReg3IN_36, F(3)=>
      ImgReg3IN_35, F(2)=>ImgReg3IN_34, F(1)=>ImgReg3IN_33, F(0)=>
      ImgReg3IN_32);
   loop3_2_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(47), D(14)
      =>DATA(46), D(13)=>DATA(45), D(12)=>DATA(44), D(11)=>DATA(43), D(10)=>
      DATA(42), D(9)=>DATA(41), D(8)=>DATA(40), D(7)=>DATA(39), D(6)=>
      DATA(38), D(5)=>DATA(37), D(4)=>DATA(36), D(3)=>DATA(35), D(2)=>
      DATA(34), D(1)=>DATA(33), D(0)=>DATA(32), EN=>nx23606, F(15)=>
      ImgReg4IN_47, F(14)=>ImgReg4IN_46, F(13)=>ImgReg4IN_45, F(12)=>
      ImgReg4IN_44, F(11)=>ImgReg4IN_43, F(10)=>ImgReg4IN_42, F(9)=>
      ImgReg4IN_41, F(8)=>ImgReg4IN_40, F(7)=>ImgReg4IN_39, F(6)=>
      ImgReg4IN_38, F(5)=>ImgReg4IN_37, F(4)=>ImgReg4IN_36, F(3)=>
      ImgReg4IN_35, F(2)=>ImgReg4IN_34, F(1)=>ImgReg4IN_33, F(0)=>
      ImgReg4IN_32);
   loop3_2_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(47), D(14)
      =>DATA(46), D(13)=>DATA(45), D(12)=>DATA(44), D(11)=>DATA(43), D(10)=>
      DATA(42), D(9)=>DATA(41), D(8)=>DATA(40), D(7)=>DATA(39), D(6)=>
      DATA(38), D(5)=>DATA(37), D(4)=>DATA(36), D(3)=>DATA(35), D(2)=>
      DATA(34), D(1)=>DATA(33), D(0)=>DATA(32), EN=>nx23594, F(15)=>
      ImgReg5IN_47, F(14)=>ImgReg5IN_46, F(13)=>ImgReg5IN_45, F(12)=>
      ImgReg5IN_44, F(11)=>ImgReg5IN_43, F(10)=>ImgReg5IN_42, F(9)=>
      ImgReg5IN_41, F(8)=>ImgReg5IN_40, F(7)=>ImgReg5IN_39, F(6)=>
      ImgReg5IN_38, F(5)=>ImgReg5IN_37, F(4)=>ImgReg5IN_36, F(3)=>
      ImgReg5IN_35, F(2)=>ImgReg5IN_34, F(1)=>ImgReg5IN_33, F(0)=>
      ImgReg5IN_32);
   loop3_2_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_47_EXMPLR, D(14)=>OutputImg1_46_EXMPLR, D(13)=>
      OutputImg1_45_EXMPLR, D(12)=>OutputImg1_44_EXMPLR, D(11)=>
      OutputImg1_43_EXMPLR, D(10)=>OutputImg1_42_EXMPLR, D(9)=>
      OutputImg1_41_EXMPLR, D(8)=>OutputImg1_40_EXMPLR, D(7)=>
      OutputImg1_39_EXMPLR, D(6)=>OutputImg1_38_EXMPLR, D(5)=>
      OutputImg1_37_EXMPLR, D(4)=>OutputImg1_36_EXMPLR, D(3)=>
      OutputImg1_35_EXMPLR, D(2)=>OutputImg1_34_EXMPLR, D(1)=>
      OutputImg1_33_EXMPLR, D(0)=>OutputImg1_32_EXMPLR, EN=>nx23788, F(15)=>
      ImgReg0IN_47, F(14)=>ImgReg0IN_46, F(13)=>ImgReg0IN_45, F(12)=>
      ImgReg0IN_44, F(11)=>ImgReg0IN_43, F(10)=>ImgReg0IN_42, F(9)=>
      ImgReg0IN_41, F(8)=>ImgReg0IN_40, F(7)=>ImgReg0IN_39, F(6)=>
      ImgReg0IN_38, F(5)=>ImgReg0IN_37, F(4)=>ImgReg0IN_36, F(3)=>
      ImgReg0IN_35, F(2)=>ImgReg0IN_34, F(1)=>ImgReg0IN_33, F(0)=>
      ImgReg0IN_32);
   loop3_2_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_47_EXMPLR, D(14)=>OutputImg2_46_EXMPLR, D(13)=>
      OutputImg2_45_EXMPLR, D(12)=>OutputImg2_44_EXMPLR, D(11)=>
      OutputImg2_43_EXMPLR, D(10)=>OutputImg2_42_EXMPLR, D(9)=>
      OutputImg2_41_EXMPLR, D(8)=>OutputImg2_40_EXMPLR, D(7)=>
      OutputImg2_39_EXMPLR, D(6)=>OutputImg2_38_EXMPLR, D(5)=>
      OutputImg2_37_EXMPLR, D(4)=>OutputImg2_36_EXMPLR, D(3)=>
      OutputImg2_35_EXMPLR, D(2)=>OutputImg2_34_EXMPLR, D(1)=>
      OutputImg2_33_EXMPLR, D(0)=>OutputImg2_32_EXMPLR, EN=>nx23788, F(15)=>
      ImgReg1IN_47, F(14)=>ImgReg1IN_46, F(13)=>ImgReg1IN_45, F(12)=>
      ImgReg1IN_44, F(11)=>ImgReg1IN_43, F(10)=>ImgReg1IN_42, F(9)=>
      ImgReg1IN_41, F(8)=>ImgReg1IN_40, F(7)=>ImgReg1IN_39, F(6)=>
      ImgReg1IN_38, F(5)=>ImgReg1IN_37, F(4)=>ImgReg1IN_36, F(3)=>
      ImgReg1IN_35, F(2)=>ImgReg1IN_34, F(1)=>ImgReg1IN_33, F(0)=>
      ImgReg1IN_32);
   loop3_2_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_47_EXMPLR, D(14)=>OutputImg3_46_EXMPLR, D(13)=>
      OutputImg3_45_EXMPLR, D(12)=>OutputImg3_44_EXMPLR, D(11)=>
      OutputImg3_43_EXMPLR, D(10)=>OutputImg3_42_EXMPLR, D(9)=>
      OutputImg3_41_EXMPLR, D(8)=>OutputImg3_40_EXMPLR, D(7)=>
      OutputImg3_39_EXMPLR, D(6)=>OutputImg3_38_EXMPLR, D(5)=>
      OutputImg3_37_EXMPLR, D(4)=>OutputImg3_36_EXMPLR, D(3)=>
      OutputImg3_35_EXMPLR, D(2)=>OutputImg3_34_EXMPLR, D(1)=>
      OutputImg3_33_EXMPLR, D(0)=>OutputImg3_32_EXMPLR, EN=>nx23788, F(15)=>
      ImgReg2IN_47, F(14)=>ImgReg2IN_46, F(13)=>ImgReg2IN_45, F(12)=>
      ImgReg2IN_44, F(11)=>ImgReg2IN_43, F(10)=>ImgReg2IN_42, F(9)=>
      ImgReg2IN_41, F(8)=>ImgReg2IN_40, F(7)=>ImgReg2IN_39, F(6)=>
      ImgReg2IN_38, F(5)=>ImgReg2IN_37, F(4)=>ImgReg2IN_36, F(3)=>
      ImgReg2IN_35, F(2)=>ImgReg2IN_34, F(1)=>ImgReg2IN_33, F(0)=>
      ImgReg2IN_32);
   loop3_2_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_47_EXMPLR, D(14)=>OutputImg4_46_EXMPLR, D(13)=>
      OutputImg4_45_EXMPLR, D(12)=>OutputImg4_44_EXMPLR, D(11)=>
      OutputImg4_43_EXMPLR, D(10)=>OutputImg4_42_EXMPLR, D(9)=>
      OutputImg4_41_EXMPLR, D(8)=>OutputImg4_40_EXMPLR, D(7)=>
      OutputImg4_39_EXMPLR, D(6)=>OutputImg4_38_EXMPLR, D(5)=>
      OutputImg4_37_EXMPLR, D(4)=>OutputImg4_36_EXMPLR, D(3)=>
      OutputImg4_35_EXMPLR, D(2)=>OutputImg4_34_EXMPLR, D(1)=>
      OutputImg4_33_EXMPLR, D(0)=>OutputImg4_32_EXMPLR, EN=>nx23788, F(15)=>
      ImgReg3IN_47, F(14)=>ImgReg3IN_46, F(13)=>ImgReg3IN_45, F(12)=>
      ImgReg3IN_44, F(11)=>ImgReg3IN_43, F(10)=>ImgReg3IN_42, F(9)=>
      ImgReg3IN_41, F(8)=>ImgReg3IN_40, F(7)=>ImgReg3IN_39, F(6)=>
      ImgReg3IN_38, F(5)=>ImgReg3IN_37, F(4)=>ImgReg3IN_36, F(3)=>
      ImgReg3IN_35, F(2)=>ImgReg3IN_34, F(1)=>ImgReg3IN_33, F(0)=>
      ImgReg3IN_32);
   loop3_2_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_47_EXMPLR, D(14)=>OutputImg5_46_EXMPLR, D(13)=>
      OutputImg5_45_EXMPLR, D(12)=>OutputImg5_44_EXMPLR, D(11)=>
      OutputImg5_43_EXMPLR, D(10)=>OutputImg5_42_EXMPLR, D(9)=>
      OutputImg5_41_EXMPLR, D(8)=>OutputImg5_40_EXMPLR, D(7)=>
      OutputImg5_39_EXMPLR, D(6)=>OutputImg5_38_EXMPLR, D(5)=>
      OutputImg5_37_EXMPLR, D(4)=>OutputImg5_36_EXMPLR, D(3)=>
      OutputImg5_35_EXMPLR, D(2)=>OutputImg5_34_EXMPLR, D(1)=>
      OutputImg5_33_EXMPLR, D(0)=>OutputImg5_32_EXMPLR, EN=>nx23790, F(15)=>
      ImgReg4IN_47, F(14)=>ImgReg4IN_46, F(13)=>ImgReg4IN_45, F(12)=>
      ImgReg4IN_44, F(11)=>ImgReg4IN_43, F(10)=>ImgReg4IN_42, F(9)=>
      ImgReg4IN_41, F(8)=>ImgReg4IN_40, F(7)=>ImgReg4IN_39, F(6)=>
      ImgReg4IN_38, F(5)=>ImgReg4IN_37, F(4)=>ImgReg4IN_36, F(3)=>
      ImgReg4IN_35, F(2)=>ImgReg4IN_34, F(1)=>ImgReg4IN_33, F(0)=>
      ImgReg4IN_32);
   loop3_2_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_47, D(14)=>
      ImgReg0IN_46, D(13)=>ImgReg0IN_45, D(12)=>ImgReg0IN_44, D(11)=>
      ImgReg0IN_43, D(10)=>ImgReg0IN_42, D(9)=>ImgReg0IN_41, D(8)=>
      ImgReg0IN_40, D(7)=>ImgReg0IN_39, D(6)=>ImgReg0IN_38, D(5)=>
      ImgReg0IN_37, D(4)=>ImgReg0IN_36, D(3)=>ImgReg0IN_35, D(2)=>
      ImgReg0IN_34, D(1)=>ImgReg0IN_33, D(0)=>ImgReg0IN_32, CLK=>nx23840, 
      RST=>RST, EN=>nx23718, Q(15)=>OutputImg0_47_EXMPLR, Q(14)=>
      OutputImg0_46_EXMPLR, Q(13)=>OutputImg0_45_EXMPLR, Q(12)=>
      OutputImg0_44_EXMPLR, Q(11)=>OutputImg0_43_EXMPLR, Q(10)=>
      OutputImg0_42_EXMPLR, Q(9)=>OutputImg0_41_EXMPLR, Q(8)=>
      OutputImg0_40_EXMPLR, Q(7)=>OutputImg0_39_EXMPLR, Q(6)=>
      OutputImg0_38_EXMPLR, Q(5)=>OutputImg0_37_EXMPLR, Q(4)=>
      OutputImg0_36_EXMPLR, Q(3)=>OutputImg0_35_EXMPLR, Q(2)=>
      OutputImg0_34_EXMPLR, Q(1)=>OutputImg0_33_EXMPLR, Q(0)=>
      OutputImg0_32_EXMPLR);
   loop3_2_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_47, D(14)=>
      ImgReg1IN_46, D(13)=>ImgReg1IN_45, D(12)=>ImgReg1IN_44, D(11)=>
      ImgReg1IN_43, D(10)=>ImgReg1IN_42, D(9)=>ImgReg1IN_41, D(8)=>
      ImgReg1IN_40, D(7)=>ImgReg1IN_39, D(6)=>ImgReg1IN_38, D(5)=>
      ImgReg1IN_37, D(4)=>ImgReg1IN_36, D(3)=>ImgReg1IN_35, D(2)=>
      ImgReg1IN_34, D(1)=>ImgReg1IN_33, D(0)=>ImgReg1IN_32, CLK=>nx23842, 
      RST=>RST, EN=>nx23728, Q(15)=>OutputImg1_47_EXMPLR, Q(14)=>
      OutputImg1_46_EXMPLR, Q(13)=>OutputImg1_45_EXMPLR, Q(12)=>
      OutputImg1_44_EXMPLR, Q(11)=>OutputImg1_43_EXMPLR, Q(10)=>
      OutputImg1_42_EXMPLR, Q(9)=>OutputImg1_41_EXMPLR, Q(8)=>
      OutputImg1_40_EXMPLR, Q(7)=>OutputImg1_39_EXMPLR, Q(6)=>
      OutputImg1_38_EXMPLR, Q(5)=>OutputImg1_37_EXMPLR, Q(4)=>
      OutputImg1_36_EXMPLR, Q(3)=>OutputImg1_35_EXMPLR, Q(2)=>
      OutputImg1_34_EXMPLR, Q(1)=>OutputImg1_33_EXMPLR, Q(0)=>
      OutputImg1_32_EXMPLR);
   loop3_2_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_47, D(14)=>
      ImgReg2IN_46, D(13)=>ImgReg2IN_45, D(12)=>ImgReg2IN_44, D(11)=>
      ImgReg2IN_43, D(10)=>ImgReg2IN_42, D(9)=>ImgReg2IN_41, D(8)=>
      ImgReg2IN_40, D(7)=>ImgReg2IN_39, D(6)=>ImgReg2IN_38, D(5)=>
      ImgReg2IN_37, D(4)=>ImgReg2IN_36, D(3)=>ImgReg2IN_35, D(2)=>
      ImgReg2IN_34, D(1)=>ImgReg2IN_33, D(0)=>ImgReg2IN_32, CLK=>nx23842, 
      RST=>RST, EN=>nx23738, Q(15)=>OutputImg2_47_EXMPLR, Q(14)=>
      OutputImg2_46_EXMPLR, Q(13)=>OutputImg2_45_EXMPLR, Q(12)=>
      OutputImg2_44_EXMPLR, Q(11)=>OutputImg2_43_EXMPLR, Q(10)=>
      OutputImg2_42_EXMPLR, Q(9)=>OutputImg2_41_EXMPLR, Q(8)=>
      OutputImg2_40_EXMPLR, Q(7)=>OutputImg2_39_EXMPLR, Q(6)=>
      OutputImg2_38_EXMPLR, Q(5)=>OutputImg2_37_EXMPLR, Q(4)=>
      OutputImg2_36_EXMPLR, Q(3)=>OutputImg2_35_EXMPLR, Q(2)=>
      OutputImg2_34_EXMPLR, Q(1)=>OutputImg2_33_EXMPLR, Q(0)=>
      OutputImg2_32_EXMPLR);
   loop3_2_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_47, D(14)=>
      ImgReg3IN_46, D(13)=>ImgReg3IN_45, D(12)=>ImgReg3IN_44, D(11)=>
      ImgReg3IN_43, D(10)=>ImgReg3IN_42, D(9)=>ImgReg3IN_41, D(8)=>
      ImgReg3IN_40, D(7)=>ImgReg3IN_39, D(6)=>ImgReg3IN_38, D(5)=>
      ImgReg3IN_37, D(4)=>ImgReg3IN_36, D(3)=>ImgReg3IN_35, D(2)=>
      ImgReg3IN_34, D(1)=>ImgReg3IN_33, D(0)=>ImgReg3IN_32, CLK=>nx23844, 
      RST=>RST, EN=>nx23748, Q(15)=>OutputImg3_47_EXMPLR, Q(14)=>
      OutputImg3_46_EXMPLR, Q(13)=>OutputImg3_45_EXMPLR, Q(12)=>
      OutputImg3_44_EXMPLR, Q(11)=>OutputImg3_43_EXMPLR, Q(10)=>
      OutputImg3_42_EXMPLR, Q(9)=>OutputImg3_41_EXMPLR, Q(8)=>
      OutputImg3_40_EXMPLR, Q(7)=>OutputImg3_39_EXMPLR, Q(6)=>
      OutputImg3_38_EXMPLR, Q(5)=>OutputImg3_37_EXMPLR, Q(4)=>
      OutputImg3_36_EXMPLR, Q(3)=>OutputImg3_35_EXMPLR, Q(2)=>
      OutputImg3_34_EXMPLR, Q(1)=>OutputImg3_33_EXMPLR, Q(0)=>
      OutputImg3_32_EXMPLR);
   loop3_2_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_47, D(14)=>
      ImgReg4IN_46, D(13)=>ImgReg4IN_45, D(12)=>ImgReg4IN_44, D(11)=>
      ImgReg4IN_43, D(10)=>ImgReg4IN_42, D(9)=>ImgReg4IN_41, D(8)=>
      ImgReg4IN_40, D(7)=>ImgReg4IN_39, D(6)=>ImgReg4IN_38, D(5)=>
      ImgReg4IN_37, D(4)=>ImgReg4IN_36, D(3)=>ImgReg4IN_35, D(2)=>
      ImgReg4IN_34, D(1)=>ImgReg4IN_33, D(0)=>ImgReg4IN_32, CLK=>nx23844, 
      RST=>RST, EN=>nx23758, Q(15)=>OutputImg4_47_EXMPLR, Q(14)=>
      OutputImg4_46_EXMPLR, Q(13)=>OutputImg4_45_EXMPLR, Q(12)=>
      OutputImg4_44_EXMPLR, Q(11)=>OutputImg4_43_EXMPLR, Q(10)=>
      OutputImg4_42_EXMPLR, Q(9)=>OutputImg4_41_EXMPLR, Q(8)=>
      OutputImg4_40_EXMPLR, Q(7)=>OutputImg4_39_EXMPLR, Q(6)=>
      OutputImg4_38_EXMPLR, Q(5)=>OutputImg4_37_EXMPLR, Q(4)=>
      OutputImg4_36_EXMPLR, Q(3)=>OutputImg4_35_EXMPLR, Q(2)=>
      OutputImg4_34_EXMPLR, Q(1)=>OutputImg4_33_EXMPLR, Q(0)=>
      OutputImg4_32_EXMPLR);
   loop3_2_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_47, D(14)=>
      ImgReg5IN_46, D(13)=>ImgReg5IN_45, D(12)=>ImgReg5IN_44, D(11)=>
      ImgReg5IN_43, D(10)=>ImgReg5IN_42, D(9)=>ImgReg5IN_41, D(8)=>
      ImgReg5IN_40, D(7)=>ImgReg5IN_39, D(6)=>ImgReg5IN_38, D(5)=>
      ImgReg5IN_37, D(4)=>ImgReg5IN_36, D(3)=>ImgReg5IN_35, D(2)=>
      ImgReg5IN_34, D(1)=>ImgReg5IN_33, D(0)=>ImgReg5IN_32, CLK=>nx23846, 
      RST=>RST, EN=>nx23768, Q(15)=>OutputImg5_47_EXMPLR, Q(14)=>
      OutputImg5_46_EXMPLR, Q(13)=>OutputImg5_45_EXMPLR, Q(12)=>
      OutputImg5_44_EXMPLR, Q(11)=>OutputImg5_43_EXMPLR, Q(10)=>
      OutputImg5_42_EXMPLR, Q(9)=>OutputImg5_41_EXMPLR, Q(8)=>
      OutputImg5_40_EXMPLR, Q(7)=>OutputImg5_39_EXMPLR, Q(6)=>
      OutputImg5_38_EXMPLR, Q(5)=>OutputImg5_37_EXMPLR, Q(4)=>
      OutputImg5_36_EXMPLR, Q(3)=>OutputImg5_35_EXMPLR, Q(2)=>
      OutputImg5_34_EXMPLR, Q(1)=>OutputImg5_33_EXMPLR, Q(0)=>
      OutputImg5_32_EXMPLR);
   loop3_3_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_79_EXMPLR, D(14)=>OutputImg0_78_EXMPLR, D(13)=>
      OutputImg0_77_EXMPLR, D(12)=>OutputImg0_76_EXMPLR, D(11)=>
      OutputImg0_75_EXMPLR, D(10)=>OutputImg0_74_EXMPLR, D(9)=>
      OutputImg0_73_EXMPLR, D(8)=>OutputImg0_72_EXMPLR, D(7)=>
      OutputImg0_71_EXMPLR, D(6)=>OutputImg0_70_EXMPLR, D(5)=>
      OutputImg0_69_EXMPLR, D(4)=>OutputImg0_68_EXMPLR, D(3)=>
      OutputImg0_67_EXMPLR, D(2)=>OutputImg0_66_EXMPLR, D(1)=>
      OutputImg0_65_EXMPLR, D(0)=>OutputImg0_64_EXMPLR, EN=>nx23670, F(15)=>
      ImgReg0IN_63, F(14)=>ImgReg0IN_62, F(13)=>ImgReg0IN_61, F(12)=>
      ImgReg0IN_60, F(11)=>ImgReg0IN_59, F(10)=>ImgReg0IN_58, F(9)=>
      ImgReg0IN_57, F(8)=>ImgReg0IN_56, F(7)=>ImgReg0IN_55, F(6)=>
      ImgReg0IN_54, F(5)=>ImgReg0IN_53, F(4)=>ImgReg0IN_52, F(3)=>
      ImgReg0IN_51, F(2)=>ImgReg0IN_50, F(1)=>ImgReg0IN_49, F(0)=>
      ImgReg0IN_48);
   loop3_3_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_79_EXMPLR, D(14)=>OutputImg1_78_EXMPLR, D(13)=>
      OutputImg1_77_EXMPLR, D(12)=>OutputImg1_76_EXMPLR, D(11)=>
      OutputImg1_75_EXMPLR, D(10)=>OutputImg1_74_EXMPLR, D(9)=>
      OutputImg1_73_EXMPLR, D(8)=>OutputImg1_72_EXMPLR, D(7)=>
      OutputImg1_71_EXMPLR, D(6)=>OutputImg1_70_EXMPLR, D(5)=>
      OutputImg1_69_EXMPLR, D(4)=>OutputImg1_68_EXMPLR, D(3)=>
      OutputImg1_67_EXMPLR, D(2)=>OutputImg1_66_EXMPLR, D(1)=>
      OutputImg1_65_EXMPLR, D(0)=>OutputImg1_64_EXMPLR, EN=>nx23670, F(15)=>
      ImgReg1IN_63, F(14)=>ImgReg1IN_62, F(13)=>ImgReg1IN_61, F(12)=>
      ImgReg1IN_60, F(11)=>ImgReg1IN_59, F(10)=>ImgReg1IN_58, F(9)=>
      ImgReg1IN_57, F(8)=>ImgReg1IN_56, F(7)=>ImgReg1IN_55, F(6)=>
      ImgReg1IN_54, F(5)=>ImgReg1IN_53, F(4)=>ImgReg1IN_52, F(3)=>
      ImgReg1IN_51, F(2)=>ImgReg1IN_50, F(1)=>ImgReg1IN_49, F(0)=>
      ImgReg1IN_48);
   loop3_3_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_79_EXMPLR, D(14)=>OutputImg2_78_EXMPLR, D(13)=>
      OutputImg2_77_EXMPLR, D(12)=>OutputImg2_76_EXMPLR, D(11)=>
      OutputImg2_75_EXMPLR, D(10)=>OutputImg2_74_EXMPLR, D(9)=>
      OutputImg2_73_EXMPLR, D(8)=>OutputImg2_72_EXMPLR, D(7)=>
      OutputImg2_71_EXMPLR, D(6)=>OutputImg2_70_EXMPLR, D(5)=>
      OutputImg2_69_EXMPLR, D(4)=>OutputImg2_68_EXMPLR, D(3)=>
      OutputImg2_67_EXMPLR, D(2)=>OutputImg2_66_EXMPLR, D(1)=>
      OutputImg2_65_EXMPLR, D(0)=>OutputImg2_64_EXMPLR, EN=>nx23670, F(15)=>
      ImgReg2IN_63, F(14)=>ImgReg2IN_62, F(13)=>ImgReg2IN_61, F(12)=>
      ImgReg2IN_60, F(11)=>ImgReg2IN_59, F(10)=>ImgReg2IN_58, F(9)=>
      ImgReg2IN_57, F(8)=>ImgReg2IN_56, F(7)=>ImgReg2IN_55, F(6)=>
      ImgReg2IN_54, F(5)=>ImgReg2IN_53, F(4)=>ImgReg2IN_52, F(3)=>
      ImgReg2IN_51, F(2)=>ImgReg2IN_50, F(1)=>ImgReg2IN_49, F(0)=>
      ImgReg2IN_48);
   loop3_3_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_79_EXMPLR, D(14)=>OutputImg3_78_EXMPLR, D(13)=>
      OutputImg3_77_EXMPLR, D(12)=>OutputImg3_76_EXMPLR, D(11)=>
      OutputImg3_75_EXMPLR, D(10)=>OutputImg3_74_EXMPLR, D(9)=>
      OutputImg3_73_EXMPLR, D(8)=>OutputImg3_72_EXMPLR, D(7)=>
      OutputImg3_71_EXMPLR, D(6)=>OutputImg3_70_EXMPLR, D(5)=>
      OutputImg3_69_EXMPLR, D(4)=>OutputImg3_68_EXMPLR, D(3)=>
      OutputImg3_67_EXMPLR, D(2)=>OutputImg3_66_EXMPLR, D(1)=>
      OutputImg3_65_EXMPLR, D(0)=>OutputImg3_64_EXMPLR, EN=>nx23672, F(15)=>
      ImgReg3IN_63, F(14)=>ImgReg3IN_62, F(13)=>ImgReg3IN_61, F(12)=>
      ImgReg3IN_60, F(11)=>ImgReg3IN_59, F(10)=>ImgReg3IN_58, F(9)=>
      ImgReg3IN_57, F(8)=>ImgReg3IN_56, F(7)=>ImgReg3IN_55, F(6)=>
      ImgReg3IN_54, F(5)=>ImgReg3IN_53, F(4)=>ImgReg3IN_52, F(3)=>
      ImgReg3IN_51, F(2)=>ImgReg3IN_50, F(1)=>ImgReg3IN_49, F(0)=>
      ImgReg3IN_48);
   loop3_3_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_79_EXMPLR, D(14)=>OutputImg4_78_EXMPLR, D(13)=>
      OutputImg4_77_EXMPLR, D(12)=>OutputImg4_76_EXMPLR, D(11)=>
      OutputImg4_75_EXMPLR, D(10)=>OutputImg4_74_EXMPLR, D(9)=>
      OutputImg4_73_EXMPLR, D(8)=>OutputImg4_72_EXMPLR, D(7)=>
      OutputImg4_71_EXMPLR, D(6)=>OutputImg4_70_EXMPLR, D(5)=>
      OutputImg4_69_EXMPLR, D(4)=>OutputImg4_68_EXMPLR, D(3)=>
      OutputImg4_67_EXMPLR, D(2)=>OutputImg4_66_EXMPLR, D(1)=>
      OutputImg4_65_EXMPLR, D(0)=>OutputImg4_64_EXMPLR, EN=>nx23672, F(15)=>
      ImgReg4IN_63, F(14)=>ImgReg4IN_62, F(13)=>ImgReg4IN_61, F(12)=>
      ImgReg4IN_60, F(11)=>ImgReg4IN_59, F(10)=>ImgReg4IN_58, F(9)=>
      ImgReg4IN_57, F(8)=>ImgReg4IN_56, F(7)=>ImgReg4IN_55, F(6)=>
      ImgReg4IN_54, F(5)=>ImgReg4IN_53, F(4)=>ImgReg4IN_52, F(3)=>
      ImgReg4IN_51, F(2)=>ImgReg4IN_50, F(1)=>ImgReg4IN_49, F(0)=>
      ImgReg4IN_48);
   loop3_3_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_79_EXMPLR, D(14)=>OutputImg5_78_EXMPLR, D(13)=>
      OutputImg5_77_EXMPLR, D(12)=>OutputImg5_76_EXMPLR, D(11)=>
      OutputImg5_75_EXMPLR, D(10)=>OutputImg5_74_EXMPLR, D(9)=>
      OutputImg5_73_EXMPLR, D(8)=>OutputImg5_72_EXMPLR, D(7)=>
      OutputImg5_71_EXMPLR, D(6)=>OutputImg5_70_EXMPLR, D(5)=>
      OutputImg5_69_EXMPLR, D(4)=>OutputImg5_68_EXMPLR, D(3)=>
      OutputImg5_67_EXMPLR, D(2)=>OutputImg5_66_EXMPLR, D(1)=>
      OutputImg5_65_EXMPLR, D(0)=>OutputImg5_64_EXMPLR, EN=>nx23672, F(15)=>
      ImgReg5IN_63, F(14)=>ImgReg5IN_62, F(13)=>ImgReg5IN_61, F(12)=>
      ImgReg5IN_60, F(11)=>ImgReg5IN_59, F(10)=>ImgReg5IN_58, F(9)=>
      ImgReg5IN_57, F(8)=>ImgReg5IN_56, F(7)=>ImgReg5IN_55, F(6)=>
      ImgReg5IN_54, F(5)=>ImgReg5IN_53, F(4)=>ImgReg5IN_52, F(3)=>
      ImgReg5IN_51, F(2)=>ImgReg5IN_50, F(1)=>ImgReg5IN_49, F(0)=>
      ImgReg5IN_48);
   loop3_3_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(63), D(14)
      =>DATA(62), D(13)=>DATA(61), D(12)=>DATA(60), D(11)=>DATA(59), D(10)=>
      DATA(58), D(9)=>DATA(57), D(8)=>DATA(56), D(7)=>DATA(55), D(6)=>
      DATA(54), D(5)=>DATA(53), D(4)=>DATA(52), D(3)=>DATA(51), D(2)=>
      DATA(50), D(1)=>DATA(49), D(0)=>DATA(48), EN=>nx23654, F(15)=>
      ImgReg0IN_63, F(14)=>ImgReg0IN_62, F(13)=>ImgReg0IN_61, F(12)=>
      ImgReg0IN_60, F(11)=>ImgReg0IN_59, F(10)=>ImgReg0IN_58, F(9)=>
      ImgReg0IN_57, F(8)=>ImgReg0IN_56, F(7)=>ImgReg0IN_55, F(6)=>
      ImgReg0IN_54, F(5)=>ImgReg0IN_53, F(4)=>ImgReg0IN_52, F(3)=>
      ImgReg0IN_51, F(2)=>ImgReg0IN_50, F(1)=>ImgReg0IN_49, F(0)=>
      ImgReg0IN_48);
   loop3_3_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(63), D(14)
      =>DATA(62), D(13)=>DATA(61), D(12)=>DATA(60), D(11)=>DATA(59), D(10)=>
      DATA(58), D(9)=>DATA(57), D(8)=>DATA(56), D(7)=>DATA(55), D(6)=>
      DATA(54), D(5)=>DATA(53), D(4)=>DATA(52), D(3)=>DATA(51), D(2)=>
      DATA(50), D(1)=>DATA(49), D(0)=>DATA(48), EN=>nx23642, F(15)=>
      ImgReg1IN_63, F(14)=>ImgReg1IN_62, F(13)=>ImgReg1IN_61, F(12)=>
      ImgReg1IN_60, F(11)=>ImgReg1IN_59, F(10)=>ImgReg1IN_58, F(9)=>
      ImgReg1IN_57, F(8)=>ImgReg1IN_56, F(7)=>ImgReg1IN_55, F(6)=>
      ImgReg1IN_54, F(5)=>ImgReg1IN_53, F(4)=>ImgReg1IN_52, F(3)=>
      ImgReg1IN_51, F(2)=>ImgReg1IN_50, F(1)=>ImgReg1IN_49, F(0)=>
      ImgReg1IN_48);
   loop3_3_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(63), D(14)
      =>DATA(62), D(13)=>DATA(61), D(12)=>DATA(60), D(11)=>DATA(59), D(10)=>
      DATA(58), D(9)=>DATA(57), D(8)=>DATA(56), D(7)=>DATA(55), D(6)=>
      DATA(54), D(5)=>DATA(53), D(4)=>DATA(52), D(3)=>DATA(51), D(2)=>
      DATA(50), D(1)=>DATA(49), D(0)=>DATA(48), EN=>nx23630, F(15)=>
      ImgReg2IN_63, F(14)=>ImgReg2IN_62, F(13)=>ImgReg2IN_61, F(12)=>
      ImgReg2IN_60, F(11)=>ImgReg2IN_59, F(10)=>ImgReg2IN_58, F(9)=>
      ImgReg2IN_57, F(8)=>ImgReg2IN_56, F(7)=>ImgReg2IN_55, F(6)=>
      ImgReg2IN_54, F(5)=>ImgReg2IN_53, F(4)=>ImgReg2IN_52, F(3)=>
      ImgReg2IN_51, F(2)=>ImgReg2IN_50, F(1)=>ImgReg2IN_49, F(0)=>
      ImgReg2IN_48);
   loop3_3_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(63), D(14)
      =>DATA(62), D(13)=>DATA(61), D(12)=>DATA(60), D(11)=>DATA(59), D(10)=>
      DATA(58), D(9)=>DATA(57), D(8)=>DATA(56), D(7)=>DATA(55), D(6)=>
      DATA(54), D(5)=>DATA(53), D(4)=>DATA(52), D(3)=>DATA(51), D(2)=>
      DATA(50), D(1)=>DATA(49), D(0)=>DATA(48), EN=>nx23618, F(15)=>
      ImgReg3IN_63, F(14)=>ImgReg3IN_62, F(13)=>ImgReg3IN_61, F(12)=>
      ImgReg3IN_60, F(11)=>ImgReg3IN_59, F(10)=>ImgReg3IN_58, F(9)=>
      ImgReg3IN_57, F(8)=>ImgReg3IN_56, F(7)=>ImgReg3IN_55, F(6)=>
      ImgReg3IN_54, F(5)=>ImgReg3IN_53, F(4)=>ImgReg3IN_52, F(3)=>
      ImgReg3IN_51, F(2)=>ImgReg3IN_50, F(1)=>ImgReg3IN_49, F(0)=>
      ImgReg3IN_48);
   loop3_3_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(63), D(14)
      =>DATA(62), D(13)=>DATA(61), D(12)=>DATA(60), D(11)=>DATA(59), D(10)=>
      DATA(58), D(9)=>DATA(57), D(8)=>DATA(56), D(7)=>DATA(55), D(6)=>
      DATA(54), D(5)=>DATA(53), D(4)=>DATA(52), D(3)=>DATA(51), D(2)=>
      DATA(50), D(1)=>DATA(49), D(0)=>DATA(48), EN=>nx23606, F(15)=>
      ImgReg4IN_63, F(14)=>ImgReg4IN_62, F(13)=>ImgReg4IN_61, F(12)=>
      ImgReg4IN_60, F(11)=>ImgReg4IN_59, F(10)=>ImgReg4IN_58, F(9)=>
      ImgReg4IN_57, F(8)=>ImgReg4IN_56, F(7)=>ImgReg4IN_55, F(6)=>
      ImgReg4IN_54, F(5)=>ImgReg4IN_53, F(4)=>ImgReg4IN_52, F(3)=>
      ImgReg4IN_51, F(2)=>ImgReg4IN_50, F(1)=>ImgReg4IN_49, F(0)=>
      ImgReg4IN_48);
   loop3_3_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(63), D(14)
      =>DATA(62), D(13)=>DATA(61), D(12)=>DATA(60), D(11)=>DATA(59), D(10)=>
      DATA(58), D(9)=>DATA(57), D(8)=>DATA(56), D(7)=>DATA(55), D(6)=>
      DATA(54), D(5)=>DATA(53), D(4)=>DATA(52), D(3)=>DATA(51), D(2)=>
      DATA(50), D(1)=>DATA(49), D(0)=>DATA(48), EN=>nx23594, F(15)=>
      ImgReg5IN_63, F(14)=>ImgReg5IN_62, F(13)=>ImgReg5IN_61, F(12)=>
      ImgReg5IN_60, F(11)=>ImgReg5IN_59, F(10)=>ImgReg5IN_58, F(9)=>
      ImgReg5IN_57, F(8)=>ImgReg5IN_56, F(7)=>ImgReg5IN_55, F(6)=>
      ImgReg5IN_54, F(5)=>ImgReg5IN_53, F(4)=>ImgReg5IN_52, F(3)=>
      ImgReg5IN_51, F(2)=>ImgReg5IN_50, F(1)=>ImgReg5IN_49, F(0)=>
      ImgReg5IN_48);
   loop3_3_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_63_EXMPLR, D(14)=>OutputImg1_62_EXMPLR, D(13)=>
      OutputImg1_61_EXMPLR, D(12)=>OutputImg1_60_EXMPLR, D(11)=>
      OutputImg1_59_EXMPLR, D(10)=>OutputImg1_58_EXMPLR, D(9)=>
      OutputImg1_57_EXMPLR, D(8)=>OutputImg1_56_EXMPLR, D(7)=>
      OutputImg1_55_EXMPLR, D(6)=>OutputImg1_54_EXMPLR, D(5)=>
      OutputImg1_53_EXMPLR, D(4)=>OutputImg1_52_EXMPLR, D(3)=>
      OutputImg1_51_EXMPLR, D(2)=>OutputImg1_50_EXMPLR, D(1)=>
      OutputImg1_49_EXMPLR, D(0)=>OutputImg1_48_EXMPLR, EN=>nx23790, F(15)=>
      ImgReg0IN_63, F(14)=>ImgReg0IN_62, F(13)=>ImgReg0IN_61, F(12)=>
      ImgReg0IN_60, F(11)=>ImgReg0IN_59, F(10)=>ImgReg0IN_58, F(9)=>
      ImgReg0IN_57, F(8)=>ImgReg0IN_56, F(7)=>ImgReg0IN_55, F(6)=>
      ImgReg0IN_54, F(5)=>ImgReg0IN_53, F(4)=>ImgReg0IN_52, F(3)=>
      ImgReg0IN_51, F(2)=>ImgReg0IN_50, F(1)=>ImgReg0IN_49, F(0)=>
      ImgReg0IN_48);
   loop3_3_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_63_EXMPLR, D(14)=>OutputImg2_62_EXMPLR, D(13)=>
      OutputImg2_61_EXMPLR, D(12)=>OutputImg2_60_EXMPLR, D(11)=>
      OutputImg2_59_EXMPLR, D(10)=>OutputImg2_58_EXMPLR, D(9)=>
      OutputImg2_57_EXMPLR, D(8)=>OutputImg2_56_EXMPLR, D(7)=>
      OutputImg2_55_EXMPLR, D(6)=>OutputImg2_54_EXMPLR, D(5)=>
      OutputImg2_53_EXMPLR, D(4)=>OutputImg2_52_EXMPLR, D(3)=>
      OutputImg2_51_EXMPLR, D(2)=>OutputImg2_50_EXMPLR, D(1)=>
      OutputImg2_49_EXMPLR, D(0)=>OutputImg2_48_EXMPLR, EN=>nx23790, F(15)=>
      ImgReg1IN_63, F(14)=>ImgReg1IN_62, F(13)=>ImgReg1IN_61, F(12)=>
      ImgReg1IN_60, F(11)=>ImgReg1IN_59, F(10)=>ImgReg1IN_58, F(9)=>
      ImgReg1IN_57, F(8)=>ImgReg1IN_56, F(7)=>ImgReg1IN_55, F(6)=>
      ImgReg1IN_54, F(5)=>ImgReg1IN_53, F(4)=>ImgReg1IN_52, F(3)=>
      ImgReg1IN_51, F(2)=>ImgReg1IN_50, F(1)=>ImgReg1IN_49, F(0)=>
      ImgReg1IN_48);
   loop3_3_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_63_EXMPLR, D(14)=>OutputImg3_62_EXMPLR, D(13)=>
      OutputImg3_61_EXMPLR, D(12)=>OutputImg3_60_EXMPLR, D(11)=>
      OutputImg3_59_EXMPLR, D(10)=>OutputImg3_58_EXMPLR, D(9)=>
      OutputImg3_57_EXMPLR, D(8)=>OutputImg3_56_EXMPLR, D(7)=>
      OutputImg3_55_EXMPLR, D(6)=>OutputImg3_54_EXMPLR, D(5)=>
      OutputImg3_53_EXMPLR, D(4)=>OutputImg3_52_EXMPLR, D(3)=>
      OutputImg3_51_EXMPLR, D(2)=>OutputImg3_50_EXMPLR, D(1)=>
      OutputImg3_49_EXMPLR, D(0)=>OutputImg3_48_EXMPLR, EN=>nx23790, F(15)=>
      ImgReg2IN_63, F(14)=>ImgReg2IN_62, F(13)=>ImgReg2IN_61, F(12)=>
      ImgReg2IN_60, F(11)=>ImgReg2IN_59, F(10)=>ImgReg2IN_58, F(9)=>
      ImgReg2IN_57, F(8)=>ImgReg2IN_56, F(7)=>ImgReg2IN_55, F(6)=>
      ImgReg2IN_54, F(5)=>ImgReg2IN_53, F(4)=>ImgReg2IN_52, F(3)=>
      ImgReg2IN_51, F(2)=>ImgReg2IN_50, F(1)=>ImgReg2IN_49, F(0)=>
      ImgReg2IN_48);
   loop3_3_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_63_EXMPLR, D(14)=>OutputImg4_62_EXMPLR, D(13)=>
      OutputImg4_61_EXMPLR, D(12)=>OutputImg4_60_EXMPLR, D(11)=>
      OutputImg4_59_EXMPLR, D(10)=>OutputImg4_58_EXMPLR, D(9)=>
      OutputImg4_57_EXMPLR, D(8)=>OutputImg4_56_EXMPLR, D(7)=>
      OutputImg4_55_EXMPLR, D(6)=>OutputImg4_54_EXMPLR, D(5)=>
      OutputImg4_53_EXMPLR, D(4)=>OutputImg4_52_EXMPLR, D(3)=>
      OutputImg4_51_EXMPLR, D(2)=>OutputImg4_50_EXMPLR, D(1)=>
      OutputImg4_49_EXMPLR, D(0)=>OutputImg4_48_EXMPLR, EN=>nx23790, F(15)=>
      ImgReg3IN_63, F(14)=>ImgReg3IN_62, F(13)=>ImgReg3IN_61, F(12)=>
      ImgReg3IN_60, F(11)=>ImgReg3IN_59, F(10)=>ImgReg3IN_58, F(9)=>
      ImgReg3IN_57, F(8)=>ImgReg3IN_56, F(7)=>ImgReg3IN_55, F(6)=>
      ImgReg3IN_54, F(5)=>ImgReg3IN_53, F(4)=>ImgReg3IN_52, F(3)=>
      ImgReg3IN_51, F(2)=>ImgReg3IN_50, F(1)=>ImgReg3IN_49, F(0)=>
      ImgReg3IN_48);
   loop3_3_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_63_EXMPLR, D(14)=>OutputImg5_62_EXMPLR, D(13)=>
      OutputImg5_61_EXMPLR, D(12)=>OutputImg5_60_EXMPLR, D(11)=>
      OutputImg5_59_EXMPLR, D(10)=>OutputImg5_58_EXMPLR, D(9)=>
      OutputImg5_57_EXMPLR, D(8)=>OutputImg5_56_EXMPLR, D(7)=>
      OutputImg5_55_EXMPLR, D(6)=>OutputImg5_54_EXMPLR, D(5)=>
      OutputImg5_53_EXMPLR, D(4)=>OutputImg5_52_EXMPLR, D(3)=>
      OutputImg5_51_EXMPLR, D(2)=>OutputImg5_50_EXMPLR, D(1)=>
      OutputImg5_49_EXMPLR, D(0)=>OutputImg5_48_EXMPLR, EN=>nx23790, F(15)=>
      ImgReg4IN_63, F(14)=>ImgReg4IN_62, F(13)=>ImgReg4IN_61, F(12)=>
      ImgReg4IN_60, F(11)=>ImgReg4IN_59, F(10)=>ImgReg4IN_58, F(9)=>
      ImgReg4IN_57, F(8)=>ImgReg4IN_56, F(7)=>ImgReg4IN_55, F(6)=>
      ImgReg4IN_54, F(5)=>ImgReg4IN_53, F(4)=>ImgReg4IN_52, F(3)=>
      ImgReg4IN_51, F(2)=>ImgReg4IN_50, F(1)=>ImgReg4IN_49, F(0)=>
      ImgReg4IN_48);
   loop3_3_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_63, D(14)=>
      ImgReg0IN_62, D(13)=>ImgReg0IN_61, D(12)=>ImgReg0IN_60, D(11)=>
      ImgReg0IN_59, D(10)=>ImgReg0IN_58, D(9)=>ImgReg0IN_57, D(8)=>
      ImgReg0IN_56, D(7)=>ImgReg0IN_55, D(6)=>ImgReg0IN_54, D(5)=>
      ImgReg0IN_53, D(4)=>ImgReg0IN_52, D(3)=>ImgReg0IN_51, D(2)=>
      ImgReg0IN_50, D(1)=>ImgReg0IN_49, D(0)=>ImgReg0IN_48, CLK=>nx23846, 
      RST=>RST, EN=>nx23718, Q(15)=>OutputImg0_63_EXMPLR, Q(14)=>
      OutputImg0_62_EXMPLR, Q(13)=>OutputImg0_61_EXMPLR, Q(12)=>
      OutputImg0_60_EXMPLR, Q(11)=>OutputImg0_59_EXMPLR, Q(10)=>
      OutputImg0_58_EXMPLR, Q(9)=>OutputImg0_57_EXMPLR, Q(8)=>
      OutputImg0_56_EXMPLR, Q(7)=>OutputImg0_55_EXMPLR, Q(6)=>
      OutputImg0_54_EXMPLR, Q(5)=>OutputImg0_53_EXMPLR, Q(4)=>
      OutputImg0_52_EXMPLR, Q(3)=>OutputImg0_51_EXMPLR, Q(2)=>
      OutputImg0_50_EXMPLR, Q(1)=>OutputImg0_49_EXMPLR, Q(0)=>
      OutputImg0_48_EXMPLR);
   loop3_3_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_63, D(14)=>
      ImgReg1IN_62, D(13)=>ImgReg1IN_61, D(12)=>ImgReg1IN_60, D(11)=>
      ImgReg1IN_59, D(10)=>ImgReg1IN_58, D(9)=>ImgReg1IN_57, D(8)=>
      ImgReg1IN_56, D(7)=>ImgReg1IN_55, D(6)=>ImgReg1IN_54, D(5)=>
      ImgReg1IN_53, D(4)=>ImgReg1IN_52, D(3)=>ImgReg1IN_51, D(2)=>
      ImgReg1IN_50, D(1)=>ImgReg1IN_49, D(0)=>ImgReg1IN_48, CLK=>nx23848, 
      RST=>RST, EN=>nx23728, Q(15)=>OutputImg1_63_EXMPLR, Q(14)=>
      OutputImg1_62_EXMPLR, Q(13)=>OutputImg1_61_EXMPLR, Q(12)=>
      OutputImg1_60_EXMPLR, Q(11)=>OutputImg1_59_EXMPLR, Q(10)=>
      OutputImg1_58_EXMPLR, Q(9)=>OutputImg1_57_EXMPLR, Q(8)=>
      OutputImg1_56_EXMPLR, Q(7)=>OutputImg1_55_EXMPLR, Q(6)=>
      OutputImg1_54_EXMPLR, Q(5)=>OutputImg1_53_EXMPLR, Q(4)=>
      OutputImg1_52_EXMPLR, Q(3)=>OutputImg1_51_EXMPLR, Q(2)=>
      OutputImg1_50_EXMPLR, Q(1)=>OutputImg1_49_EXMPLR, Q(0)=>
      OutputImg1_48_EXMPLR);
   loop3_3_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_63, D(14)=>
      ImgReg2IN_62, D(13)=>ImgReg2IN_61, D(12)=>ImgReg2IN_60, D(11)=>
      ImgReg2IN_59, D(10)=>ImgReg2IN_58, D(9)=>ImgReg2IN_57, D(8)=>
      ImgReg2IN_56, D(7)=>ImgReg2IN_55, D(6)=>ImgReg2IN_54, D(5)=>
      ImgReg2IN_53, D(4)=>ImgReg2IN_52, D(3)=>ImgReg2IN_51, D(2)=>
      ImgReg2IN_50, D(1)=>ImgReg2IN_49, D(0)=>ImgReg2IN_48, CLK=>nx23848, 
      RST=>RST, EN=>nx23738, Q(15)=>OutputImg2_63_EXMPLR, Q(14)=>
      OutputImg2_62_EXMPLR, Q(13)=>OutputImg2_61_EXMPLR, Q(12)=>
      OutputImg2_60_EXMPLR, Q(11)=>OutputImg2_59_EXMPLR, Q(10)=>
      OutputImg2_58_EXMPLR, Q(9)=>OutputImg2_57_EXMPLR, Q(8)=>
      OutputImg2_56_EXMPLR, Q(7)=>OutputImg2_55_EXMPLR, Q(6)=>
      OutputImg2_54_EXMPLR, Q(5)=>OutputImg2_53_EXMPLR, Q(4)=>
      OutputImg2_52_EXMPLR, Q(3)=>OutputImg2_51_EXMPLR, Q(2)=>
      OutputImg2_50_EXMPLR, Q(1)=>OutputImg2_49_EXMPLR, Q(0)=>
      OutputImg2_48_EXMPLR);
   loop3_3_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_63, D(14)=>
      ImgReg3IN_62, D(13)=>ImgReg3IN_61, D(12)=>ImgReg3IN_60, D(11)=>
      ImgReg3IN_59, D(10)=>ImgReg3IN_58, D(9)=>ImgReg3IN_57, D(8)=>
      ImgReg3IN_56, D(7)=>ImgReg3IN_55, D(6)=>ImgReg3IN_54, D(5)=>
      ImgReg3IN_53, D(4)=>ImgReg3IN_52, D(3)=>ImgReg3IN_51, D(2)=>
      ImgReg3IN_50, D(1)=>ImgReg3IN_49, D(0)=>ImgReg3IN_48, CLK=>nx23850, 
      RST=>RST, EN=>nx23748, Q(15)=>OutputImg3_63_EXMPLR, Q(14)=>
      OutputImg3_62_EXMPLR, Q(13)=>OutputImg3_61_EXMPLR, Q(12)=>
      OutputImg3_60_EXMPLR, Q(11)=>OutputImg3_59_EXMPLR, Q(10)=>
      OutputImg3_58_EXMPLR, Q(9)=>OutputImg3_57_EXMPLR, Q(8)=>
      OutputImg3_56_EXMPLR, Q(7)=>OutputImg3_55_EXMPLR, Q(6)=>
      OutputImg3_54_EXMPLR, Q(5)=>OutputImg3_53_EXMPLR, Q(4)=>
      OutputImg3_52_EXMPLR, Q(3)=>OutputImg3_51_EXMPLR, Q(2)=>
      OutputImg3_50_EXMPLR, Q(1)=>OutputImg3_49_EXMPLR, Q(0)=>
      OutputImg3_48_EXMPLR);
   loop3_3_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_63, D(14)=>
      ImgReg4IN_62, D(13)=>ImgReg4IN_61, D(12)=>ImgReg4IN_60, D(11)=>
      ImgReg4IN_59, D(10)=>ImgReg4IN_58, D(9)=>ImgReg4IN_57, D(8)=>
      ImgReg4IN_56, D(7)=>ImgReg4IN_55, D(6)=>ImgReg4IN_54, D(5)=>
      ImgReg4IN_53, D(4)=>ImgReg4IN_52, D(3)=>ImgReg4IN_51, D(2)=>
      ImgReg4IN_50, D(1)=>ImgReg4IN_49, D(0)=>ImgReg4IN_48, CLK=>nx23850, 
      RST=>RST, EN=>nx23758, Q(15)=>OutputImg4_63_EXMPLR, Q(14)=>
      OutputImg4_62_EXMPLR, Q(13)=>OutputImg4_61_EXMPLR, Q(12)=>
      OutputImg4_60_EXMPLR, Q(11)=>OutputImg4_59_EXMPLR, Q(10)=>
      OutputImg4_58_EXMPLR, Q(9)=>OutputImg4_57_EXMPLR, Q(8)=>
      OutputImg4_56_EXMPLR, Q(7)=>OutputImg4_55_EXMPLR, Q(6)=>
      OutputImg4_54_EXMPLR, Q(5)=>OutputImg4_53_EXMPLR, Q(4)=>
      OutputImg4_52_EXMPLR, Q(3)=>OutputImg4_51_EXMPLR, Q(2)=>
      OutputImg4_50_EXMPLR, Q(1)=>OutputImg4_49_EXMPLR, Q(0)=>
      OutputImg4_48_EXMPLR);
   loop3_3_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_63, D(14)=>
      ImgReg5IN_62, D(13)=>ImgReg5IN_61, D(12)=>ImgReg5IN_60, D(11)=>
      ImgReg5IN_59, D(10)=>ImgReg5IN_58, D(9)=>ImgReg5IN_57, D(8)=>
      ImgReg5IN_56, D(7)=>ImgReg5IN_55, D(6)=>ImgReg5IN_54, D(5)=>
      ImgReg5IN_53, D(4)=>ImgReg5IN_52, D(3)=>ImgReg5IN_51, D(2)=>
      ImgReg5IN_50, D(1)=>ImgReg5IN_49, D(0)=>ImgReg5IN_48, CLK=>nx23852, 
      RST=>RST, EN=>nx23768, Q(15)=>OutputImg5_63_EXMPLR, Q(14)=>
      OutputImg5_62_EXMPLR, Q(13)=>OutputImg5_61_EXMPLR, Q(12)=>
      OutputImg5_60_EXMPLR, Q(11)=>OutputImg5_59_EXMPLR, Q(10)=>
      OutputImg5_58_EXMPLR, Q(9)=>OutputImg5_57_EXMPLR, Q(8)=>
      OutputImg5_56_EXMPLR, Q(7)=>OutputImg5_55_EXMPLR, Q(6)=>
      OutputImg5_54_EXMPLR, Q(5)=>OutputImg5_53_EXMPLR, Q(4)=>
      OutputImg5_52_EXMPLR, Q(3)=>OutputImg5_51_EXMPLR, Q(2)=>
      OutputImg5_50_EXMPLR, Q(1)=>OutputImg5_49_EXMPLR, Q(0)=>
      OutputImg5_48_EXMPLR);
   loop3_4_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_95_EXMPLR, D(14)=>OutputImg0_94_EXMPLR, D(13)=>
      OutputImg0_93_EXMPLR, D(12)=>OutputImg0_92_EXMPLR, D(11)=>
      OutputImg0_91_EXMPLR, D(10)=>OutputImg0_90_EXMPLR, D(9)=>
      OutputImg0_89_EXMPLR, D(8)=>OutputImg0_88_EXMPLR, D(7)=>
      OutputImg0_87_EXMPLR, D(6)=>OutputImg0_86_EXMPLR, D(5)=>
      OutputImg0_85_EXMPLR, D(4)=>OutputImg0_84_EXMPLR, D(3)=>
      OutputImg0_83_EXMPLR, D(2)=>OutputImg0_82_EXMPLR, D(1)=>
      OutputImg0_81_EXMPLR, D(0)=>OutputImg0_80_EXMPLR, EN=>nx23672, F(15)=>
      ImgReg0IN_79, F(14)=>ImgReg0IN_78, F(13)=>ImgReg0IN_77, F(12)=>
      ImgReg0IN_76, F(11)=>ImgReg0IN_75, F(10)=>ImgReg0IN_74, F(9)=>
      ImgReg0IN_73, F(8)=>ImgReg0IN_72, F(7)=>ImgReg0IN_71, F(6)=>
      ImgReg0IN_70, F(5)=>ImgReg0IN_69, F(4)=>ImgReg0IN_68, F(3)=>
      ImgReg0IN_67, F(2)=>ImgReg0IN_66, F(1)=>ImgReg0IN_65, F(0)=>
      ImgReg0IN_64);
   loop3_4_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_95_EXMPLR, D(14)=>OutputImg1_94_EXMPLR, D(13)=>
      OutputImg1_93_EXMPLR, D(12)=>OutputImg1_92_EXMPLR, D(11)=>
      OutputImg1_91_EXMPLR, D(10)=>OutputImg1_90_EXMPLR, D(9)=>
      OutputImg1_89_EXMPLR, D(8)=>OutputImg1_88_EXMPLR, D(7)=>
      OutputImg1_87_EXMPLR, D(6)=>OutputImg1_86_EXMPLR, D(5)=>
      OutputImg1_85_EXMPLR, D(4)=>OutputImg1_84_EXMPLR, D(3)=>
      OutputImg1_83_EXMPLR, D(2)=>OutputImg1_82_EXMPLR, D(1)=>
      OutputImg1_81_EXMPLR, D(0)=>OutputImg1_80_EXMPLR, EN=>nx23672, F(15)=>
      ImgReg1IN_79, F(14)=>ImgReg1IN_78, F(13)=>ImgReg1IN_77, F(12)=>
      ImgReg1IN_76, F(11)=>ImgReg1IN_75, F(10)=>ImgReg1IN_74, F(9)=>
      ImgReg1IN_73, F(8)=>ImgReg1IN_72, F(7)=>ImgReg1IN_71, F(6)=>
      ImgReg1IN_70, F(5)=>ImgReg1IN_69, F(4)=>ImgReg1IN_68, F(3)=>
      ImgReg1IN_67, F(2)=>ImgReg1IN_66, F(1)=>ImgReg1IN_65, F(0)=>
      ImgReg1IN_64);
   loop3_4_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_95_EXMPLR, D(14)=>OutputImg2_94_EXMPLR, D(13)=>
      OutputImg2_93_EXMPLR, D(12)=>OutputImg2_92_EXMPLR, D(11)=>
      OutputImg2_91_EXMPLR, D(10)=>OutputImg2_90_EXMPLR, D(9)=>
      OutputImg2_89_EXMPLR, D(8)=>OutputImg2_88_EXMPLR, D(7)=>
      OutputImg2_87_EXMPLR, D(6)=>OutputImg2_86_EXMPLR, D(5)=>
      OutputImg2_85_EXMPLR, D(4)=>OutputImg2_84_EXMPLR, D(3)=>
      OutputImg2_83_EXMPLR, D(2)=>OutputImg2_82_EXMPLR, D(1)=>
      OutputImg2_81_EXMPLR, D(0)=>OutputImg2_80_EXMPLR, EN=>nx23672, F(15)=>
      ImgReg2IN_79, F(14)=>ImgReg2IN_78, F(13)=>ImgReg2IN_77, F(12)=>
      ImgReg2IN_76, F(11)=>ImgReg2IN_75, F(10)=>ImgReg2IN_74, F(9)=>
      ImgReg2IN_73, F(8)=>ImgReg2IN_72, F(7)=>ImgReg2IN_71, F(6)=>
      ImgReg2IN_70, F(5)=>ImgReg2IN_69, F(4)=>ImgReg2IN_68, F(3)=>
      ImgReg2IN_67, F(2)=>ImgReg2IN_66, F(1)=>ImgReg2IN_65, F(0)=>
      ImgReg2IN_64);
   loop3_4_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_95_EXMPLR, D(14)=>OutputImg3_94_EXMPLR, D(13)=>
      OutputImg3_93_EXMPLR, D(12)=>OutputImg3_92_EXMPLR, D(11)=>
      OutputImg3_91_EXMPLR, D(10)=>OutputImg3_90_EXMPLR, D(9)=>
      OutputImg3_89_EXMPLR, D(8)=>OutputImg3_88_EXMPLR, D(7)=>
      OutputImg3_87_EXMPLR, D(6)=>OutputImg3_86_EXMPLR, D(5)=>
      OutputImg3_85_EXMPLR, D(4)=>OutputImg3_84_EXMPLR, D(3)=>
      OutputImg3_83_EXMPLR, D(2)=>OutputImg3_82_EXMPLR, D(1)=>
      OutputImg3_81_EXMPLR, D(0)=>OutputImg3_80_EXMPLR, EN=>nx23672, F(15)=>
      ImgReg3IN_79, F(14)=>ImgReg3IN_78, F(13)=>ImgReg3IN_77, F(12)=>
      ImgReg3IN_76, F(11)=>ImgReg3IN_75, F(10)=>ImgReg3IN_74, F(9)=>
      ImgReg3IN_73, F(8)=>ImgReg3IN_72, F(7)=>ImgReg3IN_71, F(6)=>
      ImgReg3IN_70, F(5)=>ImgReg3IN_69, F(4)=>ImgReg3IN_68, F(3)=>
      ImgReg3IN_67, F(2)=>ImgReg3IN_66, F(1)=>ImgReg3IN_65, F(0)=>
      ImgReg3IN_64);
   loop3_4_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_95_EXMPLR, D(14)=>OutputImg4_94_EXMPLR, D(13)=>
      OutputImg4_93_EXMPLR, D(12)=>OutputImg4_92_EXMPLR, D(11)=>
      OutputImg4_91_EXMPLR, D(10)=>OutputImg4_90_EXMPLR, D(9)=>
      OutputImg4_89_EXMPLR, D(8)=>OutputImg4_88_EXMPLR, D(7)=>
      OutputImg4_87_EXMPLR, D(6)=>OutputImg4_86_EXMPLR, D(5)=>
      OutputImg4_85_EXMPLR, D(4)=>OutputImg4_84_EXMPLR, D(3)=>
      OutputImg4_83_EXMPLR, D(2)=>OutputImg4_82_EXMPLR, D(1)=>
      OutputImg4_81_EXMPLR, D(0)=>OutputImg4_80_EXMPLR, EN=>nx23674, F(15)=>
      ImgReg4IN_79, F(14)=>ImgReg4IN_78, F(13)=>ImgReg4IN_77, F(12)=>
      ImgReg4IN_76, F(11)=>ImgReg4IN_75, F(10)=>ImgReg4IN_74, F(9)=>
      ImgReg4IN_73, F(8)=>ImgReg4IN_72, F(7)=>ImgReg4IN_71, F(6)=>
      ImgReg4IN_70, F(5)=>ImgReg4IN_69, F(4)=>ImgReg4IN_68, F(3)=>
      ImgReg4IN_67, F(2)=>ImgReg4IN_66, F(1)=>ImgReg4IN_65, F(0)=>
      ImgReg4IN_64);
   loop3_4_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_95_EXMPLR, D(14)=>OutputImg5_94_EXMPLR, D(13)=>
      OutputImg5_93_EXMPLR, D(12)=>OutputImg5_92_EXMPLR, D(11)=>
      OutputImg5_91_EXMPLR, D(10)=>OutputImg5_90_EXMPLR, D(9)=>
      OutputImg5_89_EXMPLR, D(8)=>OutputImg5_88_EXMPLR, D(7)=>
      OutputImg5_87_EXMPLR, D(6)=>OutputImg5_86_EXMPLR, D(5)=>
      OutputImg5_85_EXMPLR, D(4)=>OutputImg5_84_EXMPLR, D(3)=>
      OutputImg5_83_EXMPLR, D(2)=>OutputImg5_82_EXMPLR, D(1)=>
      OutputImg5_81_EXMPLR, D(0)=>OutputImg5_80_EXMPLR, EN=>nx23674, F(15)=>
      ImgReg5IN_79, F(14)=>ImgReg5IN_78, F(13)=>ImgReg5IN_77, F(12)=>
      ImgReg5IN_76, F(11)=>ImgReg5IN_75, F(10)=>ImgReg5IN_74, F(9)=>
      ImgReg5IN_73, F(8)=>ImgReg5IN_72, F(7)=>ImgReg5IN_71, F(6)=>
      ImgReg5IN_70, F(5)=>ImgReg5IN_69, F(4)=>ImgReg5IN_68, F(3)=>
      ImgReg5IN_67, F(2)=>ImgReg5IN_66, F(1)=>ImgReg5IN_65, F(0)=>
      ImgReg5IN_64);
   loop3_4_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(79), D(14)
      =>DATA(78), D(13)=>DATA(77), D(12)=>DATA(76), D(11)=>DATA(75), D(10)=>
      DATA(74), D(9)=>DATA(73), D(8)=>DATA(72), D(7)=>DATA(71), D(6)=>
      DATA(70), D(5)=>DATA(69), D(4)=>DATA(68), D(3)=>DATA(67), D(2)=>
      DATA(66), D(1)=>DATA(65), D(0)=>DATA(64), EN=>nx23654, F(15)=>
      ImgReg0IN_79, F(14)=>ImgReg0IN_78, F(13)=>ImgReg0IN_77, F(12)=>
      ImgReg0IN_76, F(11)=>ImgReg0IN_75, F(10)=>ImgReg0IN_74, F(9)=>
      ImgReg0IN_73, F(8)=>ImgReg0IN_72, F(7)=>ImgReg0IN_71, F(6)=>
      ImgReg0IN_70, F(5)=>ImgReg0IN_69, F(4)=>ImgReg0IN_68, F(3)=>
      ImgReg0IN_67, F(2)=>ImgReg0IN_66, F(1)=>ImgReg0IN_65, F(0)=>
      ImgReg0IN_64);
   loop3_4_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(79), D(14)
      =>DATA(78), D(13)=>DATA(77), D(12)=>DATA(76), D(11)=>DATA(75), D(10)=>
      DATA(74), D(9)=>DATA(73), D(8)=>DATA(72), D(7)=>DATA(71), D(6)=>
      DATA(70), D(5)=>DATA(69), D(4)=>DATA(68), D(3)=>DATA(67), D(2)=>
      DATA(66), D(1)=>DATA(65), D(0)=>DATA(64), EN=>nx23642, F(15)=>
      ImgReg1IN_79, F(14)=>ImgReg1IN_78, F(13)=>ImgReg1IN_77, F(12)=>
      ImgReg1IN_76, F(11)=>ImgReg1IN_75, F(10)=>ImgReg1IN_74, F(9)=>
      ImgReg1IN_73, F(8)=>ImgReg1IN_72, F(7)=>ImgReg1IN_71, F(6)=>
      ImgReg1IN_70, F(5)=>ImgReg1IN_69, F(4)=>ImgReg1IN_68, F(3)=>
      ImgReg1IN_67, F(2)=>ImgReg1IN_66, F(1)=>ImgReg1IN_65, F(0)=>
      ImgReg1IN_64);
   loop3_4_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(79), D(14)
      =>DATA(78), D(13)=>DATA(77), D(12)=>DATA(76), D(11)=>DATA(75), D(10)=>
      DATA(74), D(9)=>DATA(73), D(8)=>DATA(72), D(7)=>DATA(71), D(6)=>
      DATA(70), D(5)=>DATA(69), D(4)=>DATA(68), D(3)=>DATA(67), D(2)=>
      DATA(66), D(1)=>DATA(65), D(0)=>DATA(64), EN=>nx23630, F(15)=>
      ImgReg2IN_79, F(14)=>ImgReg2IN_78, F(13)=>ImgReg2IN_77, F(12)=>
      ImgReg2IN_76, F(11)=>ImgReg2IN_75, F(10)=>ImgReg2IN_74, F(9)=>
      ImgReg2IN_73, F(8)=>ImgReg2IN_72, F(7)=>ImgReg2IN_71, F(6)=>
      ImgReg2IN_70, F(5)=>ImgReg2IN_69, F(4)=>ImgReg2IN_68, F(3)=>
      ImgReg2IN_67, F(2)=>ImgReg2IN_66, F(1)=>ImgReg2IN_65, F(0)=>
      ImgReg2IN_64);
   loop3_4_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(79), D(14)
      =>DATA(78), D(13)=>DATA(77), D(12)=>DATA(76), D(11)=>DATA(75), D(10)=>
      DATA(74), D(9)=>DATA(73), D(8)=>DATA(72), D(7)=>DATA(71), D(6)=>
      DATA(70), D(5)=>DATA(69), D(4)=>DATA(68), D(3)=>DATA(67), D(2)=>
      DATA(66), D(1)=>DATA(65), D(0)=>DATA(64), EN=>nx23618, F(15)=>
      ImgReg3IN_79, F(14)=>ImgReg3IN_78, F(13)=>ImgReg3IN_77, F(12)=>
      ImgReg3IN_76, F(11)=>ImgReg3IN_75, F(10)=>ImgReg3IN_74, F(9)=>
      ImgReg3IN_73, F(8)=>ImgReg3IN_72, F(7)=>ImgReg3IN_71, F(6)=>
      ImgReg3IN_70, F(5)=>ImgReg3IN_69, F(4)=>ImgReg3IN_68, F(3)=>
      ImgReg3IN_67, F(2)=>ImgReg3IN_66, F(1)=>ImgReg3IN_65, F(0)=>
      ImgReg3IN_64);
   loop3_4_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(79), D(14)
      =>DATA(78), D(13)=>DATA(77), D(12)=>DATA(76), D(11)=>DATA(75), D(10)=>
      DATA(74), D(9)=>DATA(73), D(8)=>DATA(72), D(7)=>DATA(71), D(6)=>
      DATA(70), D(5)=>DATA(69), D(4)=>DATA(68), D(3)=>DATA(67), D(2)=>
      DATA(66), D(1)=>DATA(65), D(0)=>DATA(64), EN=>nx23606, F(15)=>
      ImgReg4IN_79, F(14)=>ImgReg4IN_78, F(13)=>ImgReg4IN_77, F(12)=>
      ImgReg4IN_76, F(11)=>ImgReg4IN_75, F(10)=>ImgReg4IN_74, F(9)=>
      ImgReg4IN_73, F(8)=>ImgReg4IN_72, F(7)=>ImgReg4IN_71, F(6)=>
      ImgReg4IN_70, F(5)=>ImgReg4IN_69, F(4)=>ImgReg4IN_68, F(3)=>
      ImgReg4IN_67, F(2)=>ImgReg4IN_66, F(1)=>ImgReg4IN_65, F(0)=>
      ImgReg4IN_64);
   loop3_4_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(79), D(14)
      =>DATA(78), D(13)=>DATA(77), D(12)=>DATA(76), D(11)=>DATA(75), D(10)=>
      DATA(74), D(9)=>DATA(73), D(8)=>DATA(72), D(7)=>DATA(71), D(6)=>
      DATA(70), D(5)=>DATA(69), D(4)=>DATA(68), D(3)=>DATA(67), D(2)=>
      DATA(66), D(1)=>DATA(65), D(0)=>DATA(64), EN=>nx23594, F(15)=>
      ImgReg5IN_79, F(14)=>ImgReg5IN_78, F(13)=>ImgReg5IN_77, F(12)=>
      ImgReg5IN_76, F(11)=>ImgReg5IN_75, F(10)=>ImgReg5IN_74, F(9)=>
      ImgReg5IN_73, F(8)=>ImgReg5IN_72, F(7)=>ImgReg5IN_71, F(6)=>
      ImgReg5IN_70, F(5)=>ImgReg5IN_69, F(4)=>ImgReg5IN_68, F(3)=>
      ImgReg5IN_67, F(2)=>ImgReg5IN_66, F(1)=>ImgReg5IN_65, F(0)=>
      ImgReg5IN_64);
   loop3_4_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_79_EXMPLR, D(14)=>OutputImg1_78_EXMPLR, D(13)=>
      OutputImg1_77_EXMPLR, D(12)=>OutputImg1_76_EXMPLR, D(11)=>
      OutputImg1_75_EXMPLR, D(10)=>OutputImg1_74_EXMPLR, D(9)=>
      OutputImg1_73_EXMPLR, D(8)=>OutputImg1_72_EXMPLR, D(7)=>
      OutputImg1_71_EXMPLR, D(6)=>OutputImg1_70_EXMPLR, D(5)=>
      OutputImg1_69_EXMPLR, D(4)=>OutputImg1_68_EXMPLR, D(3)=>
      OutputImg1_67_EXMPLR, D(2)=>OutputImg1_66_EXMPLR, D(1)=>
      OutputImg1_65_EXMPLR, D(0)=>OutputImg1_64_EXMPLR, EN=>nx23790, F(15)=>
      ImgReg0IN_79, F(14)=>ImgReg0IN_78, F(13)=>ImgReg0IN_77, F(12)=>
      ImgReg0IN_76, F(11)=>ImgReg0IN_75, F(10)=>ImgReg0IN_74, F(9)=>
      ImgReg0IN_73, F(8)=>ImgReg0IN_72, F(7)=>ImgReg0IN_71, F(6)=>
      ImgReg0IN_70, F(5)=>ImgReg0IN_69, F(4)=>ImgReg0IN_68, F(3)=>
      ImgReg0IN_67, F(2)=>ImgReg0IN_66, F(1)=>ImgReg0IN_65, F(0)=>
      ImgReg0IN_64);
   loop3_4_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_79_EXMPLR, D(14)=>OutputImg2_78_EXMPLR, D(13)=>
      OutputImg2_77_EXMPLR, D(12)=>OutputImg2_76_EXMPLR, D(11)=>
      OutputImg2_75_EXMPLR, D(10)=>OutputImg2_74_EXMPLR, D(9)=>
      OutputImg2_73_EXMPLR, D(8)=>OutputImg2_72_EXMPLR, D(7)=>
      OutputImg2_71_EXMPLR, D(6)=>OutputImg2_70_EXMPLR, D(5)=>
      OutputImg2_69_EXMPLR, D(4)=>OutputImg2_68_EXMPLR, D(3)=>
      OutputImg2_67_EXMPLR, D(2)=>OutputImg2_66_EXMPLR, D(1)=>
      OutputImg2_65_EXMPLR, D(0)=>OutputImg2_64_EXMPLR, EN=>nx23792, F(15)=>
      ImgReg1IN_79, F(14)=>ImgReg1IN_78, F(13)=>ImgReg1IN_77, F(12)=>
      ImgReg1IN_76, F(11)=>ImgReg1IN_75, F(10)=>ImgReg1IN_74, F(9)=>
      ImgReg1IN_73, F(8)=>ImgReg1IN_72, F(7)=>ImgReg1IN_71, F(6)=>
      ImgReg1IN_70, F(5)=>ImgReg1IN_69, F(4)=>ImgReg1IN_68, F(3)=>
      ImgReg1IN_67, F(2)=>ImgReg1IN_66, F(1)=>ImgReg1IN_65, F(0)=>
      ImgReg1IN_64);
   loop3_4_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_79_EXMPLR, D(14)=>OutputImg3_78_EXMPLR, D(13)=>
      OutputImg3_77_EXMPLR, D(12)=>OutputImg3_76_EXMPLR, D(11)=>
      OutputImg3_75_EXMPLR, D(10)=>OutputImg3_74_EXMPLR, D(9)=>
      OutputImg3_73_EXMPLR, D(8)=>OutputImg3_72_EXMPLR, D(7)=>
      OutputImg3_71_EXMPLR, D(6)=>OutputImg3_70_EXMPLR, D(5)=>
      OutputImg3_69_EXMPLR, D(4)=>OutputImg3_68_EXMPLR, D(3)=>
      OutputImg3_67_EXMPLR, D(2)=>OutputImg3_66_EXMPLR, D(1)=>
      OutputImg3_65_EXMPLR, D(0)=>OutputImg3_64_EXMPLR, EN=>nx23792, F(15)=>
      ImgReg2IN_79, F(14)=>ImgReg2IN_78, F(13)=>ImgReg2IN_77, F(12)=>
      ImgReg2IN_76, F(11)=>ImgReg2IN_75, F(10)=>ImgReg2IN_74, F(9)=>
      ImgReg2IN_73, F(8)=>ImgReg2IN_72, F(7)=>ImgReg2IN_71, F(6)=>
      ImgReg2IN_70, F(5)=>ImgReg2IN_69, F(4)=>ImgReg2IN_68, F(3)=>
      ImgReg2IN_67, F(2)=>ImgReg2IN_66, F(1)=>ImgReg2IN_65, F(0)=>
      ImgReg2IN_64);
   loop3_4_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_79_EXMPLR, D(14)=>OutputImg4_78_EXMPLR, D(13)=>
      OutputImg4_77_EXMPLR, D(12)=>OutputImg4_76_EXMPLR, D(11)=>
      OutputImg4_75_EXMPLR, D(10)=>OutputImg4_74_EXMPLR, D(9)=>
      OutputImg4_73_EXMPLR, D(8)=>OutputImg4_72_EXMPLR, D(7)=>
      OutputImg4_71_EXMPLR, D(6)=>OutputImg4_70_EXMPLR, D(5)=>
      OutputImg4_69_EXMPLR, D(4)=>OutputImg4_68_EXMPLR, D(3)=>
      OutputImg4_67_EXMPLR, D(2)=>OutputImg4_66_EXMPLR, D(1)=>
      OutputImg4_65_EXMPLR, D(0)=>OutputImg4_64_EXMPLR, EN=>nx23792, F(15)=>
      ImgReg3IN_79, F(14)=>ImgReg3IN_78, F(13)=>ImgReg3IN_77, F(12)=>
      ImgReg3IN_76, F(11)=>ImgReg3IN_75, F(10)=>ImgReg3IN_74, F(9)=>
      ImgReg3IN_73, F(8)=>ImgReg3IN_72, F(7)=>ImgReg3IN_71, F(6)=>
      ImgReg3IN_70, F(5)=>ImgReg3IN_69, F(4)=>ImgReg3IN_68, F(3)=>
      ImgReg3IN_67, F(2)=>ImgReg3IN_66, F(1)=>ImgReg3IN_65, F(0)=>
      ImgReg3IN_64);
   loop3_4_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_79_EXMPLR, D(14)=>OutputImg5_78_EXMPLR, D(13)=>
      OutputImg5_77_EXMPLR, D(12)=>OutputImg5_76_EXMPLR, D(11)=>
      OutputImg5_75_EXMPLR, D(10)=>OutputImg5_74_EXMPLR, D(9)=>
      OutputImg5_73_EXMPLR, D(8)=>OutputImg5_72_EXMPLR, D(7)=>
      OutputImg5_71_EXMPLR, D(6)=>OutputImg5_70_EXMPLR, D(5)=>
      OutputImg5_69_EXMPLR, D(4)=>OutputImg5_68_EXMPLR, D(3)=>
      OutputImg5_67_EXMPLR, D(2)=>OutputImg5_66_EXMPLR, D(1)=>
      OutputImg5_65_EXMPLR, D(0)=>OutputImg5_64_EXMPLR, EN=>nx23792, F(15)=>
      ImgReg4IN_79, F(14)=>ImgReg4IN_78, F(13)=>ImgReg4IN_77, F(12)=>
      ImgReg4IN_76, F(11)=>ImgReg4IN_75, F(10)=>ImgReg4IN_74, F(9)=>
      ImgReg4IN_73, F(8)=>ImgReg4IN_72, F(7)=>ImgReg4IN_71, F(6)=>
      ImgReg4IN_70, F(5)=>ImgReg4IN_69, F(4)=>ImgReg4IN_68, F(3)=>
      ImgReg4IN_67, F(2)=>ImgReg4IN_66, F(1)=>ImgReg4IN_65, F(0)=>
      ImgReg4IN_64);
   loop3_4_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_79, D(14)=>
      ImgReg0IN_78, D(13)=>ImgReg0IN_77, D(12)=>ImgReg0IN_76, D(11)=>
      ImgReg0IN_75, D(10)=>ImgReg0IN_74, D(9)=>ImgReg0IN_73, D(8)=>
      ImgReg0IN_72, D(7)=>ImgReg0IN_71, D(6)=>ImgReg0IN_70, D(5)=>
      ImgReg0IN_69, D(4)=>ImgReg0IN_68, D(3)=>ImgReg0IN_67, D(2)=>
      ImgReg0IN_66, D(1)=>ImgReg0IN_65, D(0)=>ImgReg0IN_64, CLK=>nx23852, 
      RST=>RST, EN=>nx23718, Q(15)=>OutputImg0_79_EXMPLR, Q(14)=>
      OutputImg0_78_EXMPLR, Q(13)=>OutputImg0_77_EXMPLR, Q(12)=>
      OutputImg0_76_EXMPLR, Q(11)=>OutputImg0_75_EXMPLR, Q(10)=>
      OutputImg0_74_EXMPLR, Q(9)=>OutputImg0_73_EXMPLR, Q(8)=>
      OutputImg0_72_EXMPLR, Q(7)=>OutputImg0_71_EXMPLR, Q(6)=>
      OutputImg0_70_EXMPLR, Q(5)=>OutputImg0_69_EXMPLR, Q(4)=>
      OutputImg0_68_EXMPLR, Q(3)=>OutputImg0_67_EXMPLR, Q(2)=>
      OutputImg0_66_EXMPLR, Q(1)=>OutputImg0_65_EXMPLR, Q(0)=>
      OutputImg0_64_EXMPLR);
   loop3_4_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_79, D(14)=>
      ImgReg1IN_78, D(13)=>ImgReg1IN_77, D(12)=>ImgReg1IN_76, D(11)=>
      ImgReg1IN_75, D(10)=>ImgReg1IN_74, D(9)=>ImgReg1IN_73, D(8)=>
      ImgReg1IN_72, D(7)=>ImgReg1IN_71, D(6)=>ImgReg1IN_70, D(5)=>
      ImgReg1IN_69, D(4)=>ImgReg1IN_68, D(3)=>ImgReg1IN_67, D(2)=>
      ImgReg1IN_66, D(1)=>ImgReg1IN_65, D(0)=>ImgReg1IN_64, CLK=>nx23854, 
      RST=>RST, EN=>nx23728, Q(15)=>OutputImg1_79_EXMPLR, Q(14)=>
      OutputImg1_78_EXMPLR, Q(13)=>OutputImg1_77_EXMPLR, Q(12)=>
      OutputImg1_76_EXMPLR, Q(11)=>OutputImg1_75_EXMPLR, Q(10)=>
      OutputImg1_74_EXMPLR, Q(9)=>OutputImg1_73_EXMPLR, Q(8)=>
      OutputImg1_72_EXMPLR, Q(7)=>OutputImg1_71_EXMPLR, Q(6)=>
      OutputImg1_70_EXMPLR, Q(5)=>OutputImg1_69_EXMPLR, Q(4)=>
      OutputImg1_68_EXMPLR, Q(3)=>OutputImg1_67_EXMPLR, Q(2)=>
      OutputImg1_66_EXMPLR, Q(1)=>OutputImg1_65_EXMPLR, Q(0)=>
      OutputImg1_64_EXMPLR);
   loop3_4_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_79, D(14)=>
      ImgReg2IN_78, D(13)=>ImgReg2IN_77, D(12)=>ImgReg2IN_76, D(11)=>
      ImgReg2IN_75, D(10)=>ImgReg2IN_74, D(9)=>ImgReg2IN_73, D(8)=>
      ImgReg2IN_72, D(7)=>ImgReg2IN_71, D(6)=>ImgReg2IN_70, D(5)=>
      ImgReg2IN_69, D(4)=>ImgReg2IN_68, D(3)=>ImgReg2IN_67, D(2)=>
      ImgReg2IN_66, D(1)=>ImgReg2IN_65, D(0)=>ImgReg2IN_64, CLK=>nx23854, 
      RST=>RST, EN=>nx23738, Q(15)=>OutputImg2_79_EXMPLR, Q(14)=>
      OutputImg2_78_EXMPLR, Q(13)=>OutputImg2_77_EXMPLR, Q(12)=>
      OutputImg2_76_EXMPLR, Q(11)=>OutputImg2_75_EXMPLR, Q(10)=>
      OutputImg2_74_EXMPLR, Q(9)=>OutputImg2_73_EXMPLR, Q(8)=>
      OutputImg2_72_EXMPLR, Q(7)=>OutputImg2_71_EXMPLR, Q(6)=>
      OutputImg2_70_EXMPLR, Q(5)=>OutputImg2_69_EXMPLR, Q(4)=>
      OutputImg2_68_EXMPLR, Q(3)=>OutputImg2_67_EXMPLR, Q(2)=>
      OutputImg2_66_EXMPLR, Q(1)=>OutputImg2_65_EXMPLR, Q(0)=>
      OutputImg2_64_EXMPLR);
   loop3_4_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_79, D(14)=>
      ImgReg3IN_78, D(13)=>ImgReg3IN_77, D(12)=>ImgReg3IN_76, D(11)=>
      ImgReg3IN_75, D(10)=>ImgReg3IN_74, D(9)=>ImgReg3IN_73, D(8)=>
      ImgReg3IN_72, D(7)=>ImgReg3IN_71, D(6)=>ImgReg3IN_70, D(5)=>
      ImgReg3IN_69, D(4)=>ImgReg3IN_68, D(3)=>ImgReg3IN_67, D(2)=>
      ImgReg3IN_66, D(1)=>ImgReg3IN_65, D(0)=>ImgReg3IN_64, CLK=>nx23856, 
      RST=>RST, EN=>nx23748, Q(15)=>OutputImg3_79_EXMPLR, Q(14)=>
      OutputImg3_78_EXMPLR, Q(13)=>OutputImg3_77_EXMPLR, Q(12)=>
      OutputImg3_76_EXMPLR, Q(11)=>OutputImg3_75_EXMPLR, Q(10)=>
      OutputImg3_74_EXMPLR, Q(9)=>OutputImg3_73_EXMPLR, Q(8)=>
      OutputImg3_72_EXMPLR, Q(7)=>OutputImg3_71_EXMPLR, Q(6)=>
      OutputImg3_70_EXMPLR, Q(5)=>OutputImg3_69_EXMPLR, Q(4)=>
      OutputImg3_68_EXMPLR, Q(3)=>OutputImg3_67_EXMPLR, Q(2)=>
      OutputImg3_66_EXMPLR, Q(1)=>OutputImg3_65_EXMPLR, Q(0)=>
      OutputImg3_64_EXMPLR);
   loop3_4_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_79, D(14)=>
      ImgReg4IN_78, D(13)=>ImgReg4IN_77, D(12)=>ImgReg4IN_76, D(11)=>
      ImgReg4IN_75, D(10)=>ImgReg4IN_74, D(9)=>ImgReg4IN_73, D(8)=>
      ImgReg4IN_72, D(7)=>ImgReg4IN_71, D(6)=>ImgReg4IN_70, D(5)=>
      ImgReg4IN_69, D(4)=>ImgReg4IN_68, D(3)=>ImgReg4IN_67, D(2)=>
      ImgReg4IN_66, D(1)=>ImgReg4IN_65, D(0)=>ImgReg4IN_64, CLK=>nx23856, 
      RST=>RST, EN=>nx23758, Q(15)=>OutputImg4_79_EXMPLR, Q(14)=>
      OutputImg4_78_EXMPLR, Q(13)=>OutputImg4_77_EXMPLR, Q(12)=>
      OutputImg4_76_EXMPLR, Q(11)=>OutputImg4_75_EXMPLR, Q(10)=>
      OutputImg4_74_EXMPLR, Q(9)=>OutputImg4_73_EXMPLR, Q(8)=>
      OutputImg4_72_EXMPLR, Q(7)=>OutputImg4_71_EXMPLR, Q(6)=>
      OutputImg4_70_EXMPLR, Q(5)=>OutputImg4_69_EXMPLR, Q(4)=>
      OutputImg4_68_EXMPLR, Q(3)=>OutputImg4_67_EXMPLR, Q(2)=>
      OutputImg4_66_EXMPLR, Q(1)=>OutputImg4_65_EXMPLR, Q(0)=>
      OutputImg4_64_EXMPLR);
   loop3_4_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_79, D(14)=>
      ImgReg5IN_78, D(13)=>ImgReg5IN_77, D(12)=>ImgReg5IN_76, D(11)=>
      ImgReg5IN_75, D(10)=>ImgReg5IN_74, D(9)=>ImgReg5IN_73, D(8)=>
      ImgReg5IN_72, D(7)=>ImgReg5IN_71, D(6)=>ImgReg5IN_70, D(5)=>
      ImgReg5IN_69, D(4)=>ImgReg5IN_68, D(3)=>ImgReg5IN_67, D(2)=>
      ImgReg5IN_66, D(1)=>ImgReg5IN_65, D(0)=>ImgReg5IN_64, CLK=>nx23858, 
      RST=>RST, EN=>nx23768, Q(15)=>OutputImg5_79_EXMPLR, Q(14)=>
      OutputImg5_78_EXMPLR, Q(13)=>OutputImg5_77_EXMPLR, Q(12)=>
      OutputImg5_76_EXMPLR, Q(11)=>OutputImg5_75_EXMPLR, Q(10)=>
      OutputImg5_74_EXMPLR, Q(9)=>OutputImg5_73_EXMPLR, Q(8)=>
      OutputImg5_72_EXMPLR, Q(7)=>OutputImg5_71_EXMPLR, Q(6)=>
      OutputImg5_70_EXMPLR, Q(5)=>OutputImg5_69_EXMPLR, Q(4)=>
      OutputImg5_68_EXMPLR, Q(3)=>OutputImg5_67_EXMPLR, Q(2)=>
      OutputImg5_66_EXMPLR, Q(1)=>OutputImg5_65_EXMPLR, Q(0)=>
      OutputImg5_64_EXMPLR);
   loop3_5_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_111_EXMPLR, D(14)=>OutputImg0_110_EXMPLR, D(13)=>
      OutputImg0_109_EXMPLR, D(12)=>OutputImg0_108_EXMPLR, D(11)=>
      OutputImg0_107_EXMPLR, D(10)=>OutputImg0_106_EXMPLR, D(9)=>
      OutputImg0_105_EXMPLR, D(8)=>OutputImg0_104_EXMPLR, D(7)=>
      OutputImg0_103_EXMPLR, D(6)=>OutputImg0_102_EXMPLR, D(5)=>
      OutputImg0_101_EXMPLR, D(4)=>OutputImg0_100_EXMPLR, D(3)=>
      OutputImg0_99_EXMPLR, D(2)=>OutputImg0_98_EXMPLR, D(1)=>
      OutputImg0_97_EXMPLR, D(0)=>OutputImg0_96_EXMPLR, EN=>nx23674, F(15)=>
      ImgReg0IN_95, F(14)=>ImgReg0IN_94, F(13)=>ImgReg0IN_93, F(12)=>
      ImgReg0IN_92, F(11)=>ImgReg0IN_91, F(10)=>ImgReg0IN_90, F(9)=>
      ImgReg0IN_89, F(8)=>ImgReg0IN_88, F(7)=>ImgReg0IN_87, F(6)=>
      ImgReg0IN_86, F(5)=>ImgReg0IN_85, F(4)=>ImgReg0IN_84, F(3)=>
      ImgReg0IN_83, F(2)=>ImgReg0IN_82, F(1)=>ImgReg0IN_81, F(0)=>
      ImgReg0IN_80);
   loop3_5_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_111_EXMPLR, D(14)=>OutputImg1_110_EXMPLR, D(13)=>
      OutputImg1_109_EXMPLR, D(12)=>OutputImg1_108_EXMPLR, D(11)=>
      OutputImg1_107_EXMPLR, D(10)=>OutputImg1_106_EXMPLR, D(9)=>
      OutputImg1_105_EXMPLR, D(8)=>OutputImg1_104_EXMPLR, D(7)=>
      OutputImg1_103_EXMPLR, D(6)=>OutputImg1_102_EXMPLR, D(5)=>
      OutputImg1_101_EXMPLR, D(4)=>OutputImg1_100_EXMPLR, D(3)=>
      OutputImg1_99_EXMPLR, D(2)=>OutputImg1_98_EXMPLR, D(1)=>
      OutputImg1_97_EXMPLR, D(0)=>OutputImg1_96_EXMPLR, EN=>nx23674, F(15)=>
      ImgReg1IN_95, F(14)=>ImgReg1IN_94, F(13)=>ImgReg1IN_93, F(12)=>
      ImgReg1IN_92, F(11)=>ImgReg1IN_91, F(10)=>ImgReg1IN_90, F(9)=>
      ImgReg1IN_89, F(8)=>ImgReg1IN_88, F(7)=>ImgReg1IN_87, F(6)=>
      ImgReg1IN_86, F(5)=>ImgReg1IN_85, F(4)=>ImgReg1IN_84, F(3)=>
      ImgReg1IN_83, F(2)=>ImgReg1IN_82, F(1)=>ImgReg1IN_81, F(0)=>
      ImgReg1IN_80);
   loop3_5_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_111_EXMPLR, D(14)=>OutputImg2_110_EXMPLR, D(13)=>
      OutputImg2_109_EXMPLR, D(12)=>OutputImg2_108_EXMPLR, D(11)=>
      OutputImg2_107_EXMPLR, D(10)=>OutputImg2_106_EXMPLR, D(9)=>
      OutputImg2_105_EXMPLR, D(8)=>OutputImg2_104_EXMPLR, D(7)=>
      OutputImg2_103_EXMPLR, D(6)=>OutputImg2_102_EXMPLR, D(5)=>
      OutputImg2_101_EXMPLR, D(4)=>OutputImg2_100_EXMPLR, D(3)=>
      OutputImg2_99_EXMPLR, D(2)=>OutputImg2_98_EXMPLR, D(1)=>
      OutputImg2_97_EXMPLR, D(0)=>OutputImg2_96_EXMPLR, EN=>nx23674, F(15)=>
      ImgReg2IN_95, F(14)=>ImgReg2IN_94, F(13)=>ImgReg2IN_93, F(12)=>
      ImgReg2IN_92, F(11)=>ImgReg2IN_91, F(10)=>ImgReg2IN_90, F(9)=>
      ImgReg2IN_89, F(8)=>ImgReg2IN_88, F(7)=>ImgReg2IN_87, F(6)=>
      ImgReg2IN_86, F(5)=>ImgReg2IN_85, F(4)=>ImgReg2IN_84, F(3)=>
      ImgReg2IN_83, F(2)=>ImgReg2IN_82, F(1)=>ImgReg2IN_81, F(0)=>
      ImgReg2IN_80);
   loop3_5_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_111_EXMPLR, D(14)=>OutputImg3_110_EXMPLR, D(13)=>
      OutputImg3_109_EXMPLR, D(12)=>OutputImg3_108_EXMPLR, D(11)=>
      OutputImg3_107_EXMPLR, D(10)=>OutputImg3_106_EXMPLR, D(9)=>
      OutputImg3_105_EXMPLR, D(8)=>OutputImg3_104_EXMPLR, D(7)=>
      OutputImg3_103_EXMPLR, D(6)=>OutputImg3_102_EXMPLR, D(5)=>
      OutputImg3_101_EXMPLR, D(4)=>OutputImg3_100_EXMPLR, D(3)=>
      OutputImg3_99_EXMPLR, D(2)=>OutputImg3_98_EXMPLR, D(1)=>
      OutputImg3_97_EXMPLR, D(0)=>OutputImg3_96_EXMPLR, EN=>nx23674, F(15)=>
      ImgReg3IN_95, F(14)=>ImgReg3IN_94, F(13)=>ImgReg3IN_93, F(12)=>
      ImgReg3IN_92, F(11)=>ImgReg3IN_91, F(10)=>ImgReg3IN_90, F(9)=>
      ImgReg3IN_89, F(8)=>ImgReg3IN_88, F(7)=>ImgReg3IN_87, F(6)=>
      ImgReg3IN_86, F(5)=>ImgReg3IN_85, F(4)=>ImgReg3IN_84, F(3)=>
      ImgReg3IN_83, F(2)=>ImgReg3IN_82, F(1)=>ImgReg3IN_81, F(0)=>
      ImgReg3IN_80);
   loop3_5_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_111_EXMPLR, D(14)=>OutputImg4_110_EXMPLR, D(13)=>
      OutputImg4_109_EXMPLR, D(12)=>OutputImg4_108_EXMPLR, D(11)=>
      OutputImg4_107_EXMPLR, D(10)=>OutputImg4_106_EXMPLR, D(9)=>
      OutputImg4_105_EXMPLR, D(8)=>OutputImg4_104_EXMPLR, D(7)=>
      OutputImg4_103_EXMPLR, D(6)=>OutputImg4_102_EXMPLR, D(5)=>
      OutputImg4_101_EXMPLR, D(4)=>OutputImg4_100_EXMPLR, D(3)=>
      OutputImg4_99_EXMPLR, D(2)=>OutputImg4_98_EXMPLR, D(1)=>
      OutputImg4_97_EXMPLR, D(0)=>OutputImg4_96_EXMPLR, EN=>nx23674, F(15)=>
      ImgReg4IN_95, F(14)=>ImgReg4IN_94, F(13)=>ImgReg4IN_93, F(12)=>
      ImgReg4IN_92, F(11)=>ImgReg4IN_91, F(10)=>ImgReg4IN_90, F(9)=>
      ImgReg4IN_89, F(8)=>ImgReg4IN_88, F(7)=>ImgReg4IN_87, F(6)=>
      ImgReg4IN_86, F(5)=>ImgReg4IN_85, F(4)=>ImgReg4IN_84, F(3)=>
      ImgReg4IN_83, F(2)=>ImgReg4IN_82, F(1)=>ImgReg4IN_81, F(0)=>
      ImgReg4IN_80);
   loop3_5_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_111_EXMPLR, D(14)=>OutputImg5_110_EXMPLR, D(13)=>
      OutputImg5_109_EXMPLR, D(12)=>OutputImg5_108_EXMPLR, D(11)=>
      OutputImg5_107_EXMPLR, D(10)=>OutputImg5_106_EXMPLR, D(9)=>
      OutputImg5_105_EXMPLR, D(8)=>OutputImg5_104_EXMPLR, D(7)=>
      OutputImg5_103_EXMPLR, D(6)=>OutputImg5_102_EXMPLR, D(5)=>
      OutputImg5_101_EXMPLR, D(4)=>OutputImg5_100_EXMPLR, D(3)=>
      OutputImg5_99_EXMPLR, D(2)=>OutputImg5_98_EXMPLR, D(1)=>
      OutputImg5_97_EXMPLR, D(0)=>OutputImg5_96_EXMPLR, EN=>nx23676, F(15)=>
      ImgReg5IN_95, F(14)=>ImgReg5IN_94, F(13)=>ImgReg5IN_93, F(12)=>
      ImgReg5IN_92, F(11)=>ImgReg5IN_91, F(10)=>ImgReg5IN_90, F(9)=>
      ImgReg5IN_89, F(8)=>ImgReg5IN_88, F(7)=>ImgReg5IN_87, F(6)=>
      ImgReg5IN_86, F(5)=>ImgReg5IN_85, F(4)=>ImgReg5IN_84, F(3)=>
      ImgReg5IN_83, F(2)=>ImgReg5IN_82, F(1)=>ImgReg5IN_81, F(0)=>
      ImgReg5IN_80);
   loop3_5_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(95), D(14)
      =>DATA(94), D(13)=>DATA(93), D(12)=>DATA(92), D(11)=>DATA(91), D(10)=>
      DATA(90), D(9)=>DATA(89), D(8)=>DATA(88), D(7)=>DATA(87), D(6)=>
      DATA(86), D(5)=>DATA(85), D(4)=>DATA(84), D(3)=>DATA(83), D(2)=>
      DATA(82), D(1)=>DATA(81), D(0)=>DATA(80), EN=>nx23654, F(15)=>
      ImgReg0IN_95, F(14)=>ImgReg0IN_94, F(13)=>ImgReg0IN_93, F(12)=>
      ImgReg0IN_92, F(11)=>ImgReg0IN_91, F(10)=>ImgReg0IN_90, F(9)=>
      ImgReg0IN_89, F(8)=>ImgReg0IN_88, F(7)=>ImgReg0IN_87, F(6)=>
      ImgReg0IN_86, F(5)=>ImgReg0IN_85, F(4)=>ImgReg0IN_84, F(3)=>
      ImgReg0IN_83, F(2)=>ImgReg0IN_82, F(1)=>ImgReg0IN_81, F(0)=>
      ImgReg0IN_80);
   loop3_5_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(95), D(14)
      =>DATA(94), D(13)=>DATA(93), D(12)=>DATA(92), D(11)=>DATA(91), D(10)=>
      DATA(90), D(9)=>DATA(89), D(8)=>DATA(88), D(7)=>DATA(87), D(6)=>
      DATA(86), D(5)=>DATA(85), D(4)=>DATA(84), D(3)=>DATA(83), D(2)=>
      DATA(82), D(1)=>DATA(81), D(0)=>DATA(80), EN=>nx23642, F(15)=>
      ImgReg1IN_95, F(14)=>ImgReg1IN_94, F(13)=>ImgReg1IN_93, F(12)=>
      ImgReg1IN_92, F(11)=>ImgReg1IN_91, F(10)=>ImgReg1IN_90, F(9)=>
      ImgReg1IN_89, F(8)=>ImgReg1IN_88, F(7)=>ImgReg1IN_87, F(6)=>
      ImgReg1IN_86, F(5)=>ImgReg1IN_85, F(4)=>ImgReg1IN_84, F(3)=>
      ImgReg1IN_83, F(2)=>ImgReg1IN_82, F(1)=>ImgReg1IN_81, F(0)=>
      ImgReg1IN_80);
   loop3_5_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(95), D(14)
      =>DATA(94), D(13)=>DATA(93), D(12)=>DATA(92), D(11)=>DATA(91), D(10)=>
      DATA(90), D(9)=>DATA(89), D(8)=>DATA(88), D(7)=>DATA(87), D(6)=>
      DATA(86), D(5)=>DATA(85), D(4)=>DATA(84), D(3)=>DATA(83), D(2)=>
      DATA(82), D(1)=>DATA(81), D(0)=>DATA(80), EN=>nx23630, F(15)=>
      ImgReg2IN_95, F(14)=>ImgReg2IN_94, F(13)=>ImgReg2IN_93, F(12)=>
      ImgReg2IN_92, F(11)=>ImgReg2IN_91, F(10)=>ImgReg2IN_90, F(9)=>
      ImgReg2IN_89, F(8)=>ImgReg2IN_88, F(7)=>ImgReg2IN_87, F(6)=>
      ImgReg2IN_86, F(5)=>ImgReg2IN_85, F(4)=>ImgReg2IN_84, F(3)=>
      ImgReg2IN_83, F(2)=>ImgReg2IN_82, F(1)=>ImgReg2IN_81, F(0)=>
      ImgReg2IN_80);
   loop3_5_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(95), D(14)
      =>DATA(94), D(13)=>DATA(93), D(12)=>DATA(92), D(11)=>DATA(91), D(10)=>
      DATA(90), D(9)=>DATA(89), D(8)=>DATA(88), D(7)=>DATA(87), D(6)=>
      DATA(86), D(5)=>DATA(85), D(4)=>DATA(84), D(3)=>DATA(83), D(2)=>
      DATA(82), D(1)=>DATA(81), D(0)=>DATA(80), EN=>nx23618, F(15)=>
      ImgReg3IN_95, F(14)=>ImgReg3IN_94, F(13)=>ImgReg3IN_93, F(12)=>
      ImgReg3IN_92, F(11)=>ImgReg3IN_91, F(10)=>ImgReg3IN_90, F(9)=>
      ImgReg3IN_89, F(8)=>ImgReg3IN_88, F(7)=>ImgReg3IN_87, F(6)=>
      ImgReg3IN_86, F(5)=>ImgReg3IN_85, F(4)=>ImgReg3IN_84, F(3)=>
      ImgReg3IN_83, F(2)=>ImgReg3IN_82, F(1)=>ImgReg3IN_81, F(0)=>
      ImgReg3IN_80);
   loop3_5_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(95), D(14)
      =>DATA(94), D(13)=>DATA(93), D(12)=>DATA(92), D(11)=>DATA(91), D(10)=>
      DATA(90), D(9)=>DATA(89), D(8)=>DATA(88), D(7)=>DATA(87), D(6)=>
      DATA(86), D(5)=>DATA(85), D(4)=>DATA(84), D(3)=>DATA(83), D(2)=>
      DATA(82), D(1)=>DATA(81), D(0)=>DATA(80), EN=>nx23606, F(15)=>
      ImgReg4IN_95, F(14)=>ImgReg4IN_94, F(13)=>ImgReg4IN_93, F(12)=>
      ImgReg4IN_92, F(11)=>ImgReg4IN_91, F(10)=>ImgReg4IN_90, F(9)=>
      ImgReg4IN_89, F(8)=>ImgReg4IN_88, F(7)=>ImgReg4IN_87, F(6)=>
      ImgReg4IN_86, F(5)=>ImgReg4IN_85, F(4)=>ImgReg4IN_84, F(3)=>
      ImgReg4IN_83, F(2)=>ImgReg4IN_82, F(1)=>ImgReg4IN_81, F(0)=>
      ImgReg4IN_80);
   loop3_5_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(95), D(14)
      =>DATA(94), D(13)=>DATA(93), D(12)=>DATA(92), D(11)=>DATA(91), D(10)=>
      DATA(90), D(9)=>DATA(89), D(8)=>DATA(88), D(7)=>DATA(87), D(6)=>
      DATA(86), D(5)=>DATA(85), D(4)=>DATA(84), D(3)=>DATA(83), D(2)=>
      DATA(82), D(1)=>DATA(81), D(0)=>DATA(80), EN=>nx23594, F(15)=>
      ImgReg5IN_95, F(14)=>ImgReg5IN_94, F(13)=>ImgReg5IN_93, F(12)=>
      ImgReg5IN_92, F(11)=>ImgReg5IN_91, F(10)=>ImgReg5IN_90, F(9)=>
      ImgReg5IN_89, F(8)=>ImgReg5IN_88, F(7)=>ImgReg5IN_87, F(6)=>
      ImgReg5IN_86, F(5)=>ImgReg5IN_85, F(4)=>ImgReg5IN_84, F(3)=>
      ImgReg5IN_83, F(2)=>ImgReg5IN_82, F(1)=>ImgReg5IN_81, F(0)=>
      ImgReg5IN_80);
   loop3_5_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_95_EXMPLR, D(14)=>OutputImg1_94_EXMPLR, D(13)=>
      OutputImg1_93_EXMPLR, D(12)=>OutputImg1_92_EXMPLR, D(11)=>
      OutputImg1_91_EXMPLR, D(10)=>OutputImg1_90_EXMPLR, D(9)=>
      OutputImg1_89_EXMPLR, D(8)=>OutputImg1_88_EXMPLR, D(7)=>
      OutputImg1_87_EXMPLR, D(6)=>OutputImg1_86_EXMPLR, D(5)=>
      OutputImg1_85_EXMPLR, D(4)=>OutputImg1_84_EXMPLR, D(3)=>
      OutputImg1_83_EXMPLR, D(2)=>OutputImg1_82_EXMPLR, D(1)=>
      OutputImg1_81_EXMPLR, D(0)=>OutputImg1_80_EXMPLR, EN=>nx23792, F(15)=>
      ImgReg0IN_95, F(14)=>ImgReg0IN_94, F(13)=>ImgReg0IN_93, F(12)=>
      ImgReg0IN_92, F(11)=>ImgReg0IN_91, F(10)=>ImgReg0IN_90, F(9)=>
      ImgReg0IN_89, F(8)=>ImgReg0IN_88, F(7)=>ImgReg0IN_87, F(6)=>
      ImgReg0IN_86, F(5)=>ImgReg0IN_85, F(4)=>ImgReg0IN_84, F(3)=>
      ImgReg0IN_83, F(2)=>ImgReg0IN_82, F(1)=>ImgReg0IN_81, F(0)=>
      ImgReg0IN_80);
   loop3_5_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_95_EXMPLR, D(14)=>OutputImg2_94_EXMPLR, D(13)=>
      OutputImg2_93_EXMPLR, D(12)=>OutputImg2_92_EXMPLR, D(11)=>
      OutputImg2_91_EXMPLR, D(10)=>OutputImg2_90_EXMPLR, D(9)=>
      OutputImg2_89_EXMPLR, D(8)=>OutputImg2_88_EXMPLR, D(7)=>
      OutputImg2_87_EXMPLR, D(6)=>OutputImg2_86_EXMPLR, D(5)=>
      OutputImg2_85_EXMPLR, D(4)=>OutputImg2_84_EXMPLR, D(3)=>
      OutputImg2_83_EXMPLR, D(2)=>OutputImg2_82_EXMPLR, D(1)=>
      OutputImg2_81_EXMPLR, D(0)=>OutputImg2_80_EXMPLR, EN=>nx23792, F(15)=>
      ImgReg1IN_95, F(14)=>ImgReg1IN_94, F(13)=>ImgReg1IN_93, F(12)=>
      ImgReg1IN_92, F(11)=>ImgReg1IN_91, F(10)=>ImgReg1IN_90, F(9)=>
      ImgReg1IN_89, F(8)=>ImgReg1IN_88, F(7)=>ImgReg1IN_87, F(6)=>
      ImgReg1IN_86, F(5)=>ImgReg1IN_85, F(4)=>ImgReg1IN_84, F(3)=>
      ImgReg1IN_83, F(2)=>ImgReg1IN_82, F(1)=>ImgReg1IN_81, F(0)=>
      ImgReg1IN_80);
   loop3_5_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_95_EXMPLR, D(14)=>OutputImg3_94_EXMPLR, D(13)=>
      OutputImg3_93_EXMPLR, D(12)=>OutputImg3_92_EXMPLR, D(11)=>
      OutputImg3_91_EXMPLR, D(10)=>OutputImg3_90_EXMPLR, D(9)=>
      OutputImg3_89_EXMPLR, D(8)=>OutputImg3_88_EXMPLR, D(7)=>
      OutputImg3_87_EXMPLR, D(6)=>OutputImg3_86_EXMPLR, D(5)=>
      OutputImg3_85_EXMPLR, D(4)=>OutputImg3_84_EXMPLR, D(3)=>
      OutputImg3_83_EXMPLR, D(2)=>OutputImg3_82_EXMPLR, D(1)=>
      OutputImg3_81_EXMPLR, D(0)=>OutputImg3_80_EXMPLR, EN=>nx23792, F(15)=>
      ImgReg2IN_95, F(14)=>ImgReg2IN_94, F(13)=>ImgReg2IN_93, F(12)=>
      ImgReg2IN_92, F(11)=>ImgReg2IN_91, F(10)=>ImgReg2IN_90, F(9)=>
      ImgReg2IN_89, F(8)=>ImgReg2IN_88, F(7)=>ImgReg2IN_87, F(6)=>
      ImgReg2IN_86, F(5)=>ImgReg2IN_85, F(4)=>ImgReg2IN_84, F(3)=>
      ImgReg2IN_83, F(2)=>ImgReg2IN_82, F(1)=>ImgReg2IN_81, F(0)=>
      ImgReg2IN_80);
   loop3_5_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_95_EXMPLR, D(14)=>OutputImg4_94_EXMPLR, D(13)=>
      OutputImg4_93_EXMPLR, D(12)=>OutputImg4_92_EXMPLR, D(11)=>
      OutputImg4_91_EXMPLR, D(10)=>OutputImg4_90_EXMPLR, D(9)=>
      OutputImg4_89_EXMPLR, D(8)=>OutputImg4_88_EXMPLR, D(7)=>
      OutputImg4_87_EXMPLR, D(6)=>OutputImg4_86_EXMPLR, D(5)=>
      OutputImg4_85_EXMPLR, D(4)=>OutputImg4_84_EXMPLR, D(3)=>
      OutputImg4_83_EXMPLR, D(2)=>OutputImg4_82_EXMPLR, D(1)=>
      OutputImg4_81_EXMPLR, D(0)=>OutputImg4_80_EXMPLR, EN=>nx23794, F(15)=>
      ImgReg3IN_95, F(14)=>ImgReg3IN_94, F(13)=>ImgReg3IN_93, F(12)=>
      ImgReg3IN_92, F(11)=>ImgReg3IN_91, F(10)=>ImgReg3IN_90, F(9)=>
      ImgReg3IN_89, F(8)=>ImgReg3IN_88, F(7)=>ImgReg3IN_87, F(6)=>
      ImgReg3IN_86, F(5)=>ImgReg3IN_85, F(4)=>ImgReg3IN_84, F(3)=>
      ImgReg3IN_83, F(2)=>ImgReg3IN_82, F(1)=>ImgReg3IN_81, F(0)=>
      ImgReg3IN_80);
   loop3_5_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_95_EXMPLR, D(14)=>OutputImg5_94_EXMPLR, D(13)=>
      OutputImg5_93_EXMPLR, D(12)=>OutputImg5_92_EXMPLR, D(11)=>
      OutputImg5_91_EXMPLR, D(10)=>OutputImg5_90_EXMPLR, D(9)=>
      OutputImg5_89_EXMPLR, D(8)=>OutputImg5_88_EXMPLR, D(7)=>
      OutputImg5_87_EXMPLR, D(6)=>OutputImg5_86_EXMPLR, D(5)=>
      OutputImg5_85_EXMPLR, D(4)=>OutputImg5_84_EXMPLR, D(3)=>
      OutputImg5_83_EXMPLR, D(2)=>OutputImg5_82_EXMPLR, D(1)=>
      OutputImg5_81_EXMPLR, D(0)=>OutputImg5_80_EXMPLR, EN=>nx23794, F(15)=>
      ImgReg4IN_95, F(14)=>ImgReg4IN_94, F(13)=>ImgReg4IN_93, F(12)=>
      ImgReg4IN_92, F(11)=>ImgReg4IN_91, F(10)=>ImgReg4IN_90, F(9)=>
      ImgReg4IN_89, F(8)=>ImgReg4IN_88, F(7)=>ImgReg4IN_87, F(6)=>
      ImgReg4IN_86, F(5)=>ImgReg4IN_85, F(4)=>ImgReg4IN_84, F(3)=>
      ImgReg4IN_83, F(2)=>ImgReg4IN_82, F(1)=>ImgReg4IN_81, F(0)=>
      ImgReg4IN_80);
   loop3_5_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_95, D(14)=>
      ImgReg0IN_94, D(13)=>ImgReg0IN_93, D(12)=>ImgReg0IN_92, D(11)=>
      ImgReg0IN_91, D(10)=>ImgReg0IN_90, D(9)=>ImgReg0IN_89, D(8)=>
      ImgReg0IN_88, D(7)=>ImgReg0IN_87, D(6)=>ImgReg0IN_86, D(5)=>
      ImgReg0IN_85, D(4)=>ImgReg0IN_84, D(3)=>ImgReg0IN_83, D(2)=>
      ImgReg0IN_82, D(1)=>ImgReg0IN_81, D(0)=>ImgReg0IN_80, CLK=>nx23858, 
      RST=>RST, EN=>nx23718, Q(15)=>OutputImg0_95_EXMPLR, Q(14)=>
      OutputImg0_94_EXMPLR, Q(13)=>OutputImg0_93_EXMPLR, Q(12)=>
      OutputImg0_92_EXMPLR, Q(11)=>OutputImg0_91_EXMPLR, Q(10)=>
      OutputImg0_90_EXMPLR, Q(9)=>OutputImg0_89_EXMPLR, Q(8)=>
      OutputImg0_88_EXMPLR, Q(7)=>OutputImg0_87_EXMPLR, Q(6)=>
      OutputImg0_86_EXMPLR, Q(5)=>OutputImg0_85_EXMPLR, Q(4)=>
      OutputImg0_84_EXMPLR, Q(3)=>OutputImg0_83_EXMPLR, Q(2)=>
      OutputImg0_82_EXMPLR, Q(1)=>OutputImg0_81_EXMPLR, Q(0)=>
      OutputImg0_80_EXMPLR);
   loop3_5_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_95, D(14)=>
      ImgReg1IN_94, D(13)=>ImgReg1IN_93, D(12)=>ImgReg1IN_92, D(11)=>
      ImgReg1IN_91, D(10)=>ImgReg1IN_90, D(9)=>ImgReg1IN_89, D(8)=>
      ImgReg1IN_88, D(7)=>ImgReg1IN_87, D(6)=>ImgReg1IN_86, D(5)=>
      ImgReg1IN_85, D(4)=>ImgReg1IN_84, D(3)=>ImgReg1IN_83, D(2)=>
      ImgReg1IN_82, D(1)=>ImgReg1IN_81, D(0)=>ImgReg1IN_80, CLK=>nx23860, 
      RST=>RST, EN=>nx23728, Q(15)=>OutputImg1_95_EXMPLR, Q(14)=>
      OutputImg1_94_EXMPLR, Q(13)=>OutputImg1_93_EXMPLR, Q(12)=>
      OutputImg1_92_EXMPLR, Q(11)=>OutputImg1_91_EXMPLR, Q(10)=>
      OutputImg1_90_EXMPLR, Q(9)=>OutputImg1_89_EXMPLR, Q(8)=>
      OutputImg1_88_EXMPLR, Q(7)=>OutputImg1_87_EXMPLR, Q(6)=>
      OutputImg1_86_EXMPLR, Q(5)=>OutputImg1_85_EXMPLR, Q(4)=>
      OutputImg1_84_EXMPLR, Q(3)=>OutputImg1_83_EXMPLR, Q(2)=>
      OutputImg1_82_EXMPLR, Q(1)=>OutputImg1_81_EXMPLR, Q(0)=>
      OutputImg1_80_EXMPLR);
   loop3_5_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_95, D(14)=>
      ImgReg2IN_94, D(13)=>ImgReg2IN_93, D(12)=>ImgReg2IN_92, D(11)=>
      ImgReg2IN_91, D(10)=>ImgReg2IN_90, D(9)=>ImgReg2IN_89, D(8)=>
      ImgReg2IN_88, D(7)=>ImgReg2IN_87, D(6)=>ImgReg2IN_86, D(5)=>
      ImgReg2IN_85, D(4)=>ImgReg2IN_84, D(3)=>ImgReg2IN_83, D(2)=>
      ImgReg2IN_82, D(1)=>ImgReg2IN_81, D(0)=>ImgReg2IN_80, CLK=>nx23860, 
      RST=>RST, EN=>nx23738, Q(15)=>OutputImg2_95_EXMPLR, Q(14)=>
      OutputImg2_94_EXMPLR, Q(13)=>OutputImg2_93_EXMPLR, Q(12)=>
      OutputImg2_92_EXMPLR, Q(11)=>OutputImg2_91_EXMPLR, Q(10)=>
      OutputImg2_90_EXMPLR, Q(9)=>OutputImg2_89_EXMPLR, Q(8)=>
      OutputImg2_88_EXMPLR, Q(7)=>OutputImg2_87_EXMPLR, Q(6)=>
      OutputImg2_86_EXMPLR, Q(5)=>OutputImg2_85_EXMPLR, Q(4)=>
      OutputImg2_84_EXMPLR, Q(3)=>OutputImg2_83_EXMPLR, Q(2)=>
      OutputImg2_82_EXMPLR, Q(1)=>OutputImg2_81_EXMPLR, Q(0)=>
      OutputImg2_80_EXMPLR);
   loop3_5_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_95, D(14)=>
      ImgReg3IN_94, D(13)=>ImgReg3IN_93, D(12)=>ImgReg3IN_92, D(11)=>
      ImgReg3IN_91, D(10)=>ImgReg3IN_90, D(9)=>ImgReg3IN_89, D(8)=>
      ImgReg3IN_88, D(7)=>ImgReg3IN_87, D(6)=>ImgReg3IN_86, D(5)=>
      ImgReg3IN_85, D(4)=>ImgReg3IN_84, D(3)=>ImgReg3IN_83, D(2)=>
      ImgReg3IN_82, D(1)=>ImgReg3IN_81, D(0)=>ImgReg3IN_80, CLK=>nx23862, 
      RST=>RST, EN=>nx23748, Q(15)=>OutputImg3_95_EXMPLR, Q(14)=>
      OutputImg3_94_EXMPLR, Q(13)=>OutputImg3_93_EXMPLR, Q(12)=>
      OutputImg3_92_EXMPLR, Q(11)=>OutputImg3_91_EXMPLR, Q(10)=>
      OutputImg3_90_EXMPLR, Q(9)=>OutputImg3_89_EXMPLR, Q(8)=>
      OutputImg3_88_EXMPLR, Q(7)=>OutputImg3_87_EXMPLR, Q(6)=>
      OutputImg3_86_EXMPLR, Q(5)=>OutputImg3_85_EXMPLR, Q(4)=>
      OutputImg3_84_EXMPLR, Q(3)=>OutputImg3_83_EXMPLR, Q(2)=>
      OutputImg3_82_EXMPLR, Q(1)=>OutputImg3_81_EXMPLR, Q(0)=>
      OutputImg3_80_EXMPLR);
   loop3_5_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_95, D(14)=>
      ImgReg4IN_94, D(13)=>ImgReg4IN_93, D(12)=>ImgReg4IN_92, D(11)=>
      ImgReg4IN_91, D(10)=>ImgReg4IN_90, D(9)=>ImgReg4IN_89, D(8)=>
      ImgReg4IN_88, D(7)=>ImgReg4IN_87, D(6)=>ImgReg4IN_86, D(5)=>
      ImgReg4IN_85, D(4)=>ImgReg4IN_84, D(3)=>ImgReg4IN_83, D(2)=>
      ImgReg4IN_82, D(1)=>ImgReg4IN_81, D(0)=>ImgReg4IN_80, CLK=>nx23862, 
      RST=>RST, EN=>nx23758, Q(15)=>OutputImg4_95_EXMPLR, Q(14)=>
      OutputImg4_94_EXMPLR, Q(13)=>OutputImg4_93_EXMPLR, Q(12)=>
      OutputImg4_92_EXMPLR, Q(11)=>OutputImg4_91_EXMPLR, Q(10)=>
      OutputImg4_90_EXMPLR, Q(9)=>OutputImg4_89_EXMPLR, Q(8)=>
      OutputImg4_88_EXMPLR, Q(7)=>OutputImg4_87_EXMPLR, Q(6)=>
      OutputImg4_86_EXMPLR, Q(5)=>OutputImg4_85_EXMPLR, Q(4)=>
      OutputImg4_84_EXMPLR, Q(3)=>OutputImg4_83_EXMPLR, Q(2)=>
      OutputImg4_82_EXMPLR, Q(1)=>OutputImg4_81_EXMPLR, Q(0)=>
      OutputImg4_80_EXMPLR);
   loop3_5_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_95, D(14)=>
      ImgReg5IN_94, D(13)=>ImgReg5IN_93, D(12)=>ImgReg5IN_92, D(11)=>
      ImgReg5IN_91, D(10)=>ImgReg5IN_90, D(9)=>ImgReg5IN_89, D(8)=>
      ImgReg5IN_88, D(7)=>ImgReg5IN_87, D(6)=>ImgReg5IN_86, D(5)=>
      ImgReg5IN_85, D(4)=>ImgReg5IN_84, D(3)=>ImgReg5IN_83, D(2)=>
      ImgReg5IN_82, D(1)=>ImgReg5IN_81, D(0)=>ImgReg5IN_80, CLK=>nx23864, 
      RST=>RST, EN=>nx23768, Q(15)=>OutputImg5_95_EXMPLR, Q(14)=>
      OutputImg5_94_EXMPLR, Q(13)=>OutputImg5_93_EXMPLR, Q(12)=>
      OutputImg5_92_EXMPLR, Q(11)=>OutputImg5_91_EXMPLR, Q(10)=>
      OutputImg5_90_EXMPLR, Q(9)=>OutputImg5_89_EXMPLR, Q(8)=>
      OutputImg5_88_EXMPLR, Q(7)=>OutputImg5_87_EXMPLR, Q(6)=>
      OutputImg5_86_EXMPLR, Q(5)=>OutputImg5_85_EXMPLR, Q(4)=>
      OutputImg5_84_EXMPLR, Q(3)=>OutputImg5_83_EXMPLR, Q(2)=>
      OutputImg5_82_EXMPLR, Q(1)=>OutputImg5_81_EXMPLR, Q(0)=>
      OutputImg5_80_EXMPLR);
   loop3_6_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_127_EXMPLR, D(14)=>OutputImg0_126_EXMPLR, D(13)=>
      OutputImg0_125_EXMPLR, D(12)=>OutputImg0_124_EXMPLR, D(11)=>
      OutputImg0_123_EXMPLR, D(10)=>OutputImg0_122_EXMPLR, D(9)=>
      OutputImg0_121_EXMPLR, D(8)=>OutputImg0_120_EXMPLR, D(7)=>
      OutputImg0_119_EXMPLR, D(6)=>OutputImg0_118_EXMPLR, D(5)=>
      OutputImg0_117_EXMPLR, D(4)=>OutputImg0_116_EXMPLR, D(3)=>
      OutputImg0_115_EXMPLR, D(2)=>OutputImg0_114_EXMPLR, D(1)=>
      OutputImg0_113_EXMPLR, D(0)=>OutputImg0_112_EXMPLR, EN=>nx23676, F(15)
      =>ImgReg0IN_111, F(14)=>ImgReg0IN_110, F(13)=>ImgReg0IN_109, F(12)=>
      ImgReg0IN_108, F(11)=>ImgReg0IN_107, F(10)=>ImgReg0IN_106, F(9)=>
      ImgReg0IN_105, F(8)=>ImgReg0IN_104, F(7)=>ImgReg0IN_103, F(6)=>
      ImgReg0IN_102, F(5)=>ImgReg0IN_101, F(4)=>ImgReg0IN_100, F(3)=>
      ImgReg0IN_99, F(2)=>ImgReg0IN_98, F(1)=>ImgReg0IN_97, F(0)=>
      ImgReg0IN_96);
   loop3_6_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_127_EXMPLR, D(14)=>OutputImg1_126_EXMPLR, D(13)=>
      OutputImg1_125_EXMPLR, D(12)=>OutputImg1_124_EXMPLR, D(11)=>
      OutputImg1_123_EXMPLR, D(10)=>OutputImg1_122_EXMPLR, D(9)=>
      OutputImg1_121_EXMPLR, D(8)=>OutputImg1_120_EXMPLR, D(7)=>
      OutputImg1_119_EXMPLR, D(6)=>OutputImg1_118_EXMPLR, D(5)=>
      OutputImg1_117_EXMPLR, D(4)=>OutputImg1_116_EXMPLR, D(3)=>
      OutputImg1_115_EXMPLR, D(2)=>OutputImg1_114_EXMPLR, D(1)=>
      OutputImg1_113_EXMPLR, D(0)=>OutputImg1_112_EXMPLR, EN=>nx23676, F(15)
      =>ImgReg1IN_111, F(14)=>ImgReg1IN_110, F(13)=>ImgReg1IN_109, F(12)=>
      ImgReg1IN_108, F(11)=>ImgReg1IN_107, F(10)=>ImgReg1IN_106, F(9)=>
      ImgReg1IN_105, F(8)=>ImgReg1IN_104, F(7)=>ImgReg1IN_103, F(6)=>
      ImgReg1IN_102, F(5)=>ImgReg1IN_101, F(4)=>ImgReg1IN_100, F(3)=>
      ImgReg1IN_99, F(2)=>ImgReg1IN_98, F(1)=>ImgReg1IN_97, F(0)=>
      ImgReg1IN_96);
   loop3_6_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_127_EXMPLR, D(14)=>OutputImg2_126_EXMPLR, D(13)=>
      OutputImg2_125_EXMPLR, D(12)=>OutputImg2_124_EXMPLR, D(11)=>
      OutputImg2_123_EXMPLR, D(10)=>OutputImg2_122_EXMPLR, D(9)=>
      OutputImg2_121_EXMPLR, D(8)=>OutputImg2_120_EXMPLR, D(7)=>
      OutputImg2_119_EXMPLR, D(6)=>OutputImg2_118_EXMPLR, D(5)=>
      OutputImg2_117_EXMPLR, D(4)=>OutputImg2_116_EXMPLR, D(3)=>
      OutputImg2_115_EXMPLR, D(2)=>OutputImg2_114_EXMPLR, D(1)=>
      OutputImg2_113_EXMPLR, D(0)=>OutputImg2_112_EXMPLR, EN=>nx23676, F(15)
      =>ImgReg2IN_111, F(14)=>ImgReg2IN_110, F(13)=>ImgReg2IN_109, F(12)=>
      ImgReg2IN_108, F(11)=>ImgReg2IN_107, F(10)=>ImgReg2IN_106, F(9)=>
      ImgReg2IN_105, F(8)=>ImgReg2IN_104, F(7)=>ImgReg2IN_103, F(6)=>
      ImgReg2IN_102, F(5)=>ImgReg2IN_101, F(4)=>ImgReg2IN_100, F(3)=>
      ImgReg2IN_99, F(2)=>ImgReg2IN_98, F(1)=>ImgReg2IN_97, F(0)=>
      ImgReg2IN_96);
   loop3_6_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_127_EXMPLR, D(14)=>OutputImg3_126_EXMPLR, D(13)=>
      OutputImg3_125_EXMPLR, D(12)=>OutputImg3_124_EXMPLR, D(11)=>
      OutputImg3_123_EXMPLR, D(10)=>OutputImg3_122_EXMPLR, D(9)=>
      OutputImg3_121_EXMPLR, D(8)=>OutputImg3_120_EXMPLR, D(7)=>
      OutputImg3_119_EXMPLR, D(6)=>OutputImg3_118_EXMPLR, D(5)=>
      OutputImg3_117_EXMPLR, D(4)=>OutputImg3_116_EXMPLR, D(3)=>
      OutputImg3_115_EXMPLR, D(2)=>OutputImg3_114_EXMPLR, D(1)=>
      OutputImg3_113_EXMPLR, D(0)=>OutputImg3_112_EXMPLR, EN=>nx23676, F(15)
      =>ImgReg3IN_111, F(14)=>ImgReg3IN_110, F(13)=>ImgReg3IN_109, F(12)=>
      ImgReg3IN_108, F(11)=>ImgReg3IN_107, F(10)=>ImgReg3IN_106, F(9)=>
      ImgReg3IN_105, F(8)=>ImgReg3IN_104, F(7)=>ImgReg3IN_103, F(6)=>
      ImgReg3IN_102, F(5)=>ImgReg3IN_101, F(4)=>ImgReg3IN_100, F(3)=>
      ImgReg3IN_99, F(2)=>ImgReg3IN_98, F(1)=>ImgReg3IN_97, F(0)=>
      ImgReg3IN_96);
   loop3_6_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_127_EXMPLR, D(14)=>OutputImg4_126_EXMPLR, D(13)=>
      OutputImg4_125_EXMPLR, D(12)=>OutputImg4_124_EXMPLR, D(11)=>
      OutputImg4_123_EXMPLR, D(10)=>OutputImg4_122_EXMPLR, D(9)=>
      OutputImg4_121_EXMPLR, D(8)=>OutputImg4_120_EXMPLR, D(7)=>
      OutputImg4_119_EXMPLR, D(6)=>OutputImg4_118_EXMPLR, D(5)=>
      OutputImg4_117_EXMPLR, D(4)=>OutputImg4_116_EXMPLR, D(3)=>
      OutputImg4_115_EXMPLR, D(2)=>OutputImg4_114_EXMPLR, D(1)=>
      OutputImg4_113_EXMPLR, D(0)=>OutputImg4_112_EXMPLR, EN=>nx23676, F(15)
      =>ImgReg4IN_111, F(14)=>ImgReg4IN_110, F(13)=>ImgReg4IN_109, F(12)=>
      ImgReg4IN_108, F(11)=>ImgReg4IN_107, F(10)=>ImgReg4IN_106, F(9)=>
      ImgReg4IN_105, F(8)=>ImgReg4IN_104, F(7)=>ImgReg4IN_103, F(6)=>
      ImgReg4IN_102, F(5)=>ImgReg4IN_101, F(4)=>ImgReg4IN_100, F(3)=>
      ImgReg4IN_99, F(2)=>ImgReg4IN_98, F(1)=>ImgReg4IN_97, F(0)=>
      ImgReg4IN_96);
   loop3_6_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_127_EXMPLR, D(14)=>OutputImg5_126_EXMPLR, D(13)=>
      OutputImg5_125_EXMPLR, D(12)=>OutputImg5_124_EXMPLR, D(11)=>
      OutputImg5_123_EXMPLR, D(10)=>OutputImg5_122_EXMPLR, D(9)=>
      OutputImg5_121_EXMPLR, D(8)=>OutputImg5_120_EXMPLR, D(7)=>
      OutputImg5_119_EXMPLR, D(6)=>OutputImg5_118_EXMPLR, D(5)=>
      OutputImg5_117_EXMPLR, D(4)=>OutputImg5_116_EXMPLR, D(3)=>
      OutputImg5_115_EXMPLR, D(2)=>OutputImg5_114_EXMPLR, D(1)=>
      OutputImg5_113_EXMPLR, D(0)=>OutputImg5_112_EXMPLR, EN=>nx23676, F(15)
      =>ImgReg5IN_111, F(14)=>ImgReg5IN_110, F(13)=>ImgReg5IN_109, F(12)=>
      ImgReg5IN_108, F(11)=>ImgReg5IN_107, F(10)=>ImgReg5IN_106, F(9)=>
      ImgReg5IN_105, F(8)=>ImgReg5IN_104, F(7)=>ImgReg5IN_103, F(6)=>
      ImgReg5IN_102, F(5)=>ImgReg5IN_101, F(4)=>ImgReg5IN_100, F(3)=>
      ImgReg5IN_99, F(2)=>ImgReg5IN_98, F(1)=>ImgReg5IN_97, F(0)=>
      ImgReg5IN_96);
   loop3_6_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(111), D(14)
      =>DATA(110), D(13)=>DATA(109), D(12)=>DATA(108), D(11)=>DATA(107), 
      D(10)=>DATA(106), D(9)=>DATA(105), D(8)=>DATA(104), D(7)=>DATA(103), 
      D(6)=>DATA(102), D(5)=>DATA(101), D(4)=>DATA(100), D(3)=>DATA(99), 
      D(2)=>DATA(98), D(1)=>DATA(97), D(0)=>DATA(96), EN=>nx23654, F(15)=>
      ImgReg0IN_111, F(14)=>ImgReg0IN_110, F(13)=>ImgReg0IN_109, F(12)=>
      ImgReg0IN_108, F(11)=>ImgReg0IN_107, F(10)=>ImgReg0IN_106, F(9)=>
      ImgReg0IN_105, F(8)=>ImgReg0IN_104, F(7)=>ImgReg0IN_103, F(6)=>
      ImgReg0IN_102, F(5)=>ImgReg0IN_101, F(4)=>ImgReg0IN_100, F(3)=>
      ImgReg0IN_99, F(2)=>ImgReg0IN_98, F(1)=>ImgReg0IN_97, F(0)=>
      ImgReg0IN_96);
   loop3_6_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(111), D(14)
      =>DATA(110), D(13)=>DATA(109), D(12)=>DATA(108), D(11)=>DATA(107), 
      D(10)=>DATA(106), D(9)=>DATA(105), D(8)=>DATA(104), D(7)=>DATA(103), 
      D(6)=>DATA(102), D(5)=>DATA(101), D(4)=>DATA(100), D(3)=>DATA(99), 
      D(2)=>DATA(98), D(1)=>DATA(97), D(0)=>DATA(96), EN=>nx23642, F(15)=>
      ImgReg1IN_111, F(14)=>ImgReg1IN_110, F(13)=>ImgReg1IN_109, F(12)=>
      ImgReg1IN_108, F(11)=>ImgReg1IN_107, F(10)=>ImgReg1IN_106, F(9)=>
      ImgReg1IN_105, F(8)=>ImgReg1IN_104, F(7)=>ImgReg1IN_103, F(6)=>
      ImgReg1IN_102, F(5)=>ImgReg1IN_101, F(4)=>ImgReg1IN_100, F(3)=>
      ImgReg1IN_99, F(2)=>ImgReg1IN_98, F(1)=>ImgReg1IN_97, F(0)=>
      ImgReg1IN_96);
   loop3_6_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(111), D(14)
      =>DATA(110), D(13)=>DATA(109), D(12)=>DATA(108), D(11)=>DATA(107), 
      D(10)=>DATA(106), D(9)=>DATA(105), D(8)=>DATA(104), D(7)=>DATA(103), 
      D(6)=>DATA(102), D(5)=>DATA(101), D(4)=>DATA(100), D(3)=>DATA(99), 
      D(2)=>DATA(98), D(1)=>DATA(97), D(0)=>DATA(96), EN=>nx23630, F(15)=>
      ImgReg2IN_111, F(14)=>ImgReg2IN_110, F(13)=>ImgReg2IN_109, F(12)=>
      ImgReg2IN_108, F(11)=>ImgReg2IN_107, F(10)=>ImgReg2IN_106, F(9)=>
      ImgReg2IN_105, F(8)=>ImgReg2IN_104, F(7)=>ImgReg2IN_103, F(6)=>
      ImgReg2IN_102, F(5)=>ImgReg2IN_101, F(4)=>ImgReg2IN_100, F(3)=>
      ImgReg2IN_99, F(2)=>ImgReg2IN_98, F(1)=>ImgReg2IN_97, F(0)=>
      ImgReg2IN_96);
   loop3_6_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(111), D(14)
      =>DATA(110), D(13)=>DATA(109), D(12)=>DATA(108), D(11)=>DATA(107), 
      D(10)=>DATA(106), D(9)=>DATA(105), D(8)=>DATA(104), D(7)=>DATA(103), 
      D(6)=>DATA(102), D(5)=>DATA(101), D(4)=>DATA(100), D(3)=>DATA(99), 
      D(2)=>DATA(98), D(1)=>DATA(97), D(0)=>DATA(96), EN=>nx23618, F(15)=>
      ImgReg3IN_111, F(14)=>ImgReg3IN_110, F(13)=>ImgReg3IN_109, F(12)=>
      ImgReg3IN_108, F(11)=>ImgReg3IN_107, F(10)=>ImgReg3IN_106, F(9)=>
      ImgReg3IN_105, F(8)=>ImgReg3IN_104, F(7)=>ImgReg3IN_103, F(6)=>
      ImgReg3IN_102, F(5)=>ImgReg3IN_101, F(4)=>ImgReg3IN_100, F(3)=>
      ImgReg3IN_99, F(2)=>ImgReg3IN_98, F(1)=>ImgReg3IN_97, F(0)=>
      ImgReg3IN_96);
   loop3_6_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(111), D(14)
      =>DATA(110), D(13)=>DATA(109), D(12)=>DATA(108), D(11)=>DATA(107), 
      D(10)=>DATA(106), D(9)=>DATA(105), D(8)=>DATA(104), D(7)=>DATA(103), 
      D(6)=>DATA(102), D(5)=>DATA(101), D(4)=>DATA(100), D(3)=>DATA(99), 
      D(2)=>DATA(98), D(1)=>DATA(97), D(0)=>DATA(96), EN=>nx23606, F(15)=>
      ImgReg4IN_111, F(14)=>ImgReg4IN_110, F(13)=>ImgReg4IN_109, F(12)=>
      ImgReg4IN_108, F(11)=>ImgReg4IN_107, F(10)=>ImgReg4IN_106, F(9)=>
      ImgReg4IN_105, F(8)=>ImgReg4IN_104, F(7)=>ImgReg4IN_103, F(6)=>
      ImgReg4IN_102, F(5)=>ImgReg4IN_101, F(4)=>ImgReg4IN_100, F(3)=>
      ImgReg4IN_99, F(2)=>ImgReg4IN_98, F(1)=>ImgReg4IN_97, F(0)=>
      ImgReg4IN_96);
   loop3_6_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(111), D(14)
      =>DATA(110), D(13)=>DATA(109), D(12)=>DATA(108), D(11)=>DATA(107), 
      D(10)=>DATA(106), D(9)=>DATA(105), D(8)=>DATA(104), D(7)=>DATA(103), 
      D(6)=>DATA(102), D(5)=>DATA(101), D(4)=>DATA(100), D(3)=>DATA(99), 
      D(2)=>DATA(98), D(1)=>DATA(97), D(0)=>DATA(96), EN=>nx23594, F(15)=>
      ImgReg5IN_111, F(14)=>ImgReg5IN_110, F(13)=>ImgReg5IN_109, F(12)=>
      ImgReg5IN_108, F(11)=>ImgReg5IN_107, F(10)=>ImgReg5IN_106, F(9)=>
      ImgReg5IN_105, F(8)=>ImgReg5IN_104, F(7)=>ImgReg5IN_103, F(6)=>
      ImgReg5IN_102, F(5)=>ImgReg5IN_101, F(4)=>ImgReg5IN_100, F(3)=>
      ImgReg5IN_99, F(2)=>ImgReg5IN_98, F(1)=>ImgReg5IN_97, F(0)=>
      ImgReg5IN_96);
   loop3_6_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_111_EXMPLR, D(14)=>OutputImg1_110_EXMPLR, D(13)=>
      OutputImg1_109_EXMPLR, D(12)=>OutputImg1_108_EXMPLR, D(11)=>
      OutputImg1_107_EXMPLR, D(10)=>OutputImg1_106_EXMPLR, D(9)=>
      OutputImg1_105_EXMPLR, D(8)=>OutputImg1_104_EXMPLR, D(7)=>
      OutputImg1_103_EXMPLR, D(6)=>OutputImg1_102_EXMPLR, D(5)=>
      OutputImg1_101_EXMPLR, D(4)=>OutputImg1_100_EXMPLR, D(3)=>
      OutputImg1_99_EXMPLR, D(2)=>OutputImg1_98_EXMPLR, D(1)=>
      OutputImg1_97_EXMPLR, D(0)=>OutputImg1_96_EXMPLR, EN=>nx23794, F(15)=>
      ImgReg0IN_111, F(14)=>ImgReg0IN_110, F(13)=>ImgReg0IN_109, F(12)=>
      ImgReg0IN_108, F(11)=>ImgReg0IN_107, F(10)=>ImgReg0IN_106, F(9)=>
      ImgReg0IN_105, F(8)=>ImgReg0IN_104, F(7)=>ImgReg0IN_103, F(6)=>
      ImgReg0IN_102, F(5)=>ImgReg0IN_101, F(4)=>ImgReg0IN_100, F(3)=>
      ImgReg0IN_99, F(2)=>ImgReg0IN_98, F(1)=>ImgReg0IN_97, F(0)=>
      ImgReg0IN_96);
   loop3_6_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_111_EXMPLR, D(14)=>OutputImg2_110_EXMPLR, D(13)=>
      OutputImg2_109_EXMPLR, D(12)=>OutputImg2_108_EXMPLR, D(11)=>
      OutputImg2_107_EXMPLR, D(10)=>OutputImg2_106_EXMPLR, D(9)=>
      OutputImg2_105_EXMPLR, D(8)=>OutputImg2_104_EXMPLR, D(7)=>
      OutputImg2_103_EXMPLR, D(6)=>OutputImg2_102_EXMPLR, D(5)=>
      OutputImg2_101_EXMPLR, D(4)=>OutputImg2_100_EXMPLR, D(3)=>
      OutputImg2_99_EXMPLR, D(2)=>OutputImg2_98_EXMPLR, D(1)=>
      OutputImg2_97_EXMPLR, D(0)=>OutputImg2_96_EXMPLR, EN=>nx23794, F(15)=>
      ImgReg1IN_111, F(14)=>ImgReg1IN_110, F(13)=>ImgReg1IN_109, F(12)=>
      ImgReg1IN_108, F(11)=>ImgReg1IN_107, F(10)=>ImgReg1IN_106, F(9)=>
      ImgReg1IN_105, F(8)=>ImgReg1IN_104, F(7)=>ImgReg1IN_103, F(6)=>
      ImgReg1IN_102, F(5)=>ImgReg1IN_101, F(4)=>ImgReg1IN_100, F(3)=>
      ImgReg1IN_99, F(2)=>ImgReg1IN_98, F(1)=>ImgReg1IN_97, F(0)=>
      ImgReg1IN_96);
   loop3_6_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_111_EXMPLR, D(14)=>OutputImg3_110_EXMPLR, D(13)=>
      OutputImg3_109_EXMPLR, D(12)=>OutputImg3_108_EXMPLR, D(11)=>
      OutputImg3_107_EXMPLR, D(10)=>OutputImg3_106_EXMPLR, D(9)=>
      OutputImg3_105_EXMPLR, D(8)=>OutputImg3_104_EXMPLR, D(7)=>
      OutputImg3_103_EXMPLR, D(6)=>OutputImg3_102_EXMPLR, D(5)=>
      OutputImg3_101_EXMPLR, D(4)=>OutputImg3_100_EXMPLR, D(3)=>
      OutputImg3_99_EXMPLR, D(2)=>OutputImg3_98_EXMPLR, D(1)=>
      OutputImg3_97_EXMPLR, D(0)=>OutputImg3_96_EXMPLR, EN=>nx23794, F(15)=>
      ImgReg2IN_111, F(14)=>ImgReg2IN_110, F(13)=>ImgReg2IN_109, F(12)=>
      ImgReg2IN_108, F(11)=>ImgReg2IN_107, F(10)=>ImgReg2IN_106, F(9)=>
      ImgReg2IN_105, F(8)=>ImgReg2IN_104, F(7)=>ImgReg2IN_103, F(6)=>
      ImgReg2IN_102, F(5)=>ImgReg2IN_101, F(4)=>ImgReg2IN_100, F(3)=>
      ImgReg2IN_99, F(2)=>ImgReg2IN_98, F(1)=>ImgReg2IN_97, F(0)=>
      ImgReg2IN_96);
   loop3_6_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_111_EXMPLR, D(14)=>OutputImg4_110_EXMPLR, D(13)=>
      OutputImg4_109_EXMPLR, D(12)=>OutputImg4_108_EXMPLR, D(11)=>
      OutputImg4_107_EXMPLR, D(10)=>OutputImg4_106_EXMPLR, D(9)=>
      OutputImg4_105_EXMPLR, D(8)=>OutputImg4_104_EXMPLR, D(7)=>
      OutputImg4_103_EXMPLR, D(6)=>OutputImg4_102_EXMPLR, D(5)=>
      OutputImg4_101_EXMPLR, D(4)=>OutputImg4_100_EXMPLR, D(3)=>
      OutputImg4_99_EXMPLR, D(2)=>OutputImg4_98_EXMPLR, D(1)=>
      OutputImg4_97_EXMPLR, D(0)=>OutputImg4_96_EXMPLR, EN=>nx23794, F(15)=>
      ImgReg3IN_111, F(14)=>ImgReg3IN_110, F(13)=>ImgReg3IN_109, F(12)=>
      ImgReg3IN_108, F(11)=>ImgReg3IN_107, F(10)=>ImgReg3IN_106, F(9)=>
      ImgReg3IN_105, F(8)=>ImgReg3IN_104, F(7)=>ImgReg3IN_103, F(6)=>
      ImgReg3IN_102, F(5)=>ImgReg3IN_101, F(4)=>ImgReg3IN_100, F(3)=>
      ImgReg3IN_99, F(2)=>ImgReg3IN_98, F(1)=>ImgReg3IN_97, F(0)=>
      ImgReg3IN_96);
   loop3_6_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_111_EXMPLR, D(14)=>OutputImg5_110_EXMPLR, D(13)=>
      OutputImg5_109_EXMPLR, D(12)=>OutputImg5_108_EXMPLR, D(11)=>
      OutputImg5_107_EXMPLR, D(10)=>OutputImg5_106_EXMPLR, D(9)=>
      OutputImg5_105_EXMPLR, D(8)=>OutputImg5_104_EXMPLR, D(7)=>
      OutputImg5_103_EXMPLR, D(6)=>OutputImg5_102_EXMPLR, D(5)=>
      OutputImg5_101_EXMPLR, D(4)=>OutputImg5_100_EXMPLR, D(3)=>
      OutputImg5_99_EXMPLR, D(2)=>OutputImg5_98_EXMPLR, D(1)=>
      OutputImg5_97_EXMPLR, D(0)=>OutputImg5_96_EXMPLR, EN=>nx23794, F(15)=>
      ImgReg4IN_111, F(14)=>ImgReg4IN_110, F(13)=>ImgReg4IN_109, F(12)=>
      ImgReg4IN_108, F(11)=>ImgReg4IN_107, F(10)=>ImgReg4IN_106, F(9)=>
      ImgReg4IN_105, F(8)=>ImgReg4IN_104, F(7)=>ImgReg4IN_103, F(6)=>
      ImgReg4IN_102, F(5)=>ImgReg4IN_101, F(4)=>ImgReg4IN_100, F(3)=>
      ImgReg4IN_99, F(2)=>ImgReg4IN_98, F(1)=>ImgReg4IN_97, F(0)=>
      ImgReg4IN_96);
   loop3_6_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_111, D(14)=>
      ImgReg0IN_110, D(13)=>ImgReg0IN_109, D(12)=>ImgReg0IN_108, D(11)=>
      ImgReg0IN_107, D(10)=>ImgReg0IN_106, D(9)=>ImgReg0IN_105, D(8)=>
      ImgReg0IN_104, D(7)=>ImgReg0IN_103, D(6)=>ImgReg0IN_102, D(5)=>
      ImgReg0IN_101, D(4)=>ImgReg0IN_100, D(3)=>ImgReg0IN_99, D(2)=>
      ImgReg0IN_98, D(1)=>ImgReg0IN_97, D(0)=>ImgReg0IN_96, CLK=>nx23864, 
      RST=>RST, EN=>nx23718, Q(15)=>OutputImg0_111_EXMPLR, Q(14)=>
      OutputImg0_110_EXMPLR, Q(13)=>OutputImg0_109_EXMPLR, Q(12)=>
      OutputImg0_108_EXMPLR, Q(11)=>OutputImg0_107_EXMPLR, Q(10)=>
      OutputImg0_106_EXMPLR, Q(9)=>OutputImg0_105_EXMPLR, Q(8)=>
      OutputImg0_104_EXMPLR, Q(7)=>OutputImg0_103_EXMPLR, Q(6)=>
      OutputImg0_102_EXMPLR, Q(5)=>OutputImg0_101_EXMPLR, Q(4)=>
      OutputImg0_100_EXMPLR, Q(3)=>OutputImg0_99_EXMPLR, Q(2)=>
      OutputImg0_98_EXMPLR, Q(1)=>OutputImg0_97_EXMPLR, Q(0)=>
      OutputImg0_96_EXMPLR);
   loop3_6_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_111, D(14)=>
      ImgReg1IN_110, D(13)=>ImgReg1IN_109, D(12)=>ImgReg1IN_108, D(11)=>
      ImgReg1IN_107, D(10)=>ImgReg1IN_106, D(9)=>ImgReg1IN_105, D(8)=>
      ImgReg1IN_104, D(7)=>ImgReg1IN_103, D(6)=>ImgReg1IN_102, D(5)=>
      ImgReg1IN_101, D(4)=>ImgReg1IN_100, D(3)=>ImgReg1IN_99, D(2)=>
      ImgReg1IN_98, D(1)=>ImgReg1IN_97, D(0)=>ImgReg1IN_96, CLK=>nx23866, 
      RST=>RST, EN=>nx23728, Q(15)=>OutputImg1_111_EXMPLR, Q(14)=>
      OutputImg1_110_EXMPLR, Q(13)=>OutputImg1_109_EXMPLR, Q(12)=>
      OutputImg1_108_EXMPLR, Q(11)=>OutputImg1_107_EXMPLR, Q(10)=>
      OutputImg1_106_EXMPLR, Q(9)=>OutputImg1_105_EXMPLR, Q(8)=>
      OutputImg1_104_EXMPLR, Q(7)=>OutputImg1_103_EXMPLR, Q(6)=>
      OutputImg1_102_EXMPLR, Q(5)=>OutputImg1_101_EXMPLR, Q(4)=>
      OutputImg1_100_EXMPLR, Q(3)=>OutputImg1_99_EXMPLR, Q(2)=>
      OutputImg1_98_EXMPLR, Q(1)=>OutputImg1_97_EXMPLR, Q(0)=>
      OutputImg1_96_EXMPLR);
   loop3_6_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_111, D(14)=>
      ImgReg2IN_110, D(13)=>ImgReg2IN_109, D(12)=>ImgReg2IN_108, D(11)=>
      ImgReg2IN_107, D(10)=>ImgReg2IN_106, D(9)=>ImgReg2IN_105, D(8)=>
      ImgReg2IN_104, D(7)=>ImgReg2IN_103, D(6)=>ImgReg2IN_102, D(5)=>
      ImgReg2IN_101, D(4)=>ImgReg2IN_100, D(3)=>ImgReg2IN_99, D(2)=>
      ImgReg2IN_98, D(1)=>ImgReg2IN_97, D(0)=>ImgReg2IN_96, CLK=>nx23866, 
      RST=>RST, EN=>nx23738, Q(15)=>OutputImg2_111_EXMPLR, Q(14)=>
      OutputImg2_110_EXMPLR, Q(13)=>OutputImg2_109_EXMPLR, Q(12)=>
      OutputImg2_108_EXMPLR, Q(11)=>OutputImg2_107_EXMPLR, Q(10)=>
      OutputImg2_106_EXMPLR, Q(9)=>OutputImg2_105_EXMPLR, Q(8)=>
      OutputImg2_104_EXMPLR, Q(7)=>OutputImg2_103_EXMPLR, Q(6)=>
      OutputImg2_102_EXMPLR, Q(5)=>OutputImg2_101_EXMPLR, Q(4)=>
      OutputImg2_100_EXMPLR, Q(3)=>OutputImg2_99_EXMPLR, Q(2)=>
      OutputImg2_98_EXMPLR, Q(1)=>OutputImg2_97_EXMPLR, Q(0)=>
      OutputImg2_96_EXMPLR);
   loop3_6_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_111, D(14)=>
      ImgReg3IN_110, D(13)=>ImgReg3IN_109, D(12)=>ImgReg3IN_108, D(11)=>
      ImgReg3IN_107, D(10)=>ImgReg3IN_106, D(9)=>ImgReg3IN_105, D(8)=>
      ImgReg3IN_104, D(7)=>ImgReg3IN_103, D(6)=>ImgReg3IN_102, D(5)=>
      ImgReg3IN_101, D(4)=>ImgReg3IN_100, D(3)=>ImgReg3IN_99, D(2)=>
      ImgReg3IN_98, D(1)=>ImgReg3IN_97, D(0)=>ImgReg3IN_96, CLK=>nx23868, 
      RST=>RST, EN=>nx23748, Q(15)=>OutputImg3_111_EXMPLR, Q(14)=>
      OutputImg3_110_EXMPLR, Q(13)=>OutputImg3_109_EXMPLR, Q(12)=>
      OutputImg3_108_EXMPLR, Q(11)=>OutputImg3_107_EXMPLR, Q(10)=>
      OutputImg3_106_EXMPLR, Q(9)=>OutputImg3_105_EXMPLR, Q(8)=>
      OutputImg3_104_EXMPLR, Q(7)=>OutputImg3_103_EXMPLR, Q(6)=>
      OutputImg3_102_EXMPLR, Q(5)=>OutputImg3_101_EXMPLR, Q(4)=>
      OutputImg3_100_EXMPLR, Q(3)=>OutputImg3_99_EXMPLR, Q(2)=>
      OutputImg3_98_EXMPLR, Q(1)=>OutputImg3_97_EXMPLR, Q(0)=>
      OutputImg3_96_EXMPLR);
   loop3_6_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_111, D(14)=>
      ImgReg4IN_110, D(13)=>ImgReg4IN_109, D(12)=>ImgReg4IN_108, D(11)=>
      ImgReg4IN_107, D(10)=>ImgReg4IN_106, D(9)=>ImgReg4IN_105, D(8)=>
      ImgReg4IN_104, D(7)=>ImgReg4IN_103, D(6)=>ImgReg4IN_102, D(5)=>
      ImgReg4IN_101, D(4)=>ImgReg4IN_100, D(3)=>ImgReg4IN_99, D(2)=>
      ImgReg4IN_98, D(1)=>ImgReg4IN_97, D(0)=>ImgReg4IN_96, CLK=>nx23868, 
      RST=>RST, EN=>nx23758, Q(15)=>OutputImg4_111_EXMPLR, Q(14)=>
      OutputImg4_110_EXMPLR, Q(13)=>OutputImg4_109_EXMPLR, Q(12)=>
      OutputImg4_108_EXMPLR, Q(11)=>OutputImg4_107_EXMPLR, Q(10)=>
      OutputImg4_106_EXMPLR, Q(9)=>OutputImg4_105_EXMPLR, Q(8)=>
      OutputImg4_104_EXMPLR, Q(7)=>OutputImg4_103_EXMPLR, Q(6)=>
      OutputImg4_102_EXMPLR, Q(5)=>OutputImg4_101_EXMPLR, Q(4)=>
      OutputImg4_100_EXMPLR, Q(3)=>OutputImg4_99_EXMPLR, Q(2)=>
      OutputImg4_98_EXMPLR, Q(1)=>OutputImg4_97_EXMPLR, Q(0)=>
      OutputImg4_96_EXMPLR);
   loop3_6_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_111, D(14)=>
      ImgReg5IN_110, D(13)=>ImgReg5IN_109, D(12)=>ImgReg5IN_108, D(11)=>
      ImgReg5IN_107, D(10)=>ImgReg5IN_106, D(9)=>ImgReg5IN_105, D(8)=>
      ImgReg5IN_104, D(7)=>ImgReg5IN_103, D(6)=>ImgReg5IN_102, D(5)=>
      ImgReg5IN_101, D(4)=>ImgReg5IN_100, D(3)=>ImgReg5IN_99, D(2)=>
      ImgReg5IN_98, D(1)=>ImgReg5IN_97, D(0)=>ImgReg5IN_96, CLK=>nx23870, 
      RST=>RST, EN=>nx23768, Q(15)=>OutputImg5_111_EXMPLR, Q(14)=>
      OutputImg5_110_EXMPLR, Q(13)=>OutputImg5_109_EXMPLR, Q(12)=>
      OutputImg5_108_EXMPLR, Q(11)=>OutputImg5_107_EXMPLR, Q(10)=>
      OutputImg5_106_EXMPLR, Q(9)=>OutputImg5_105_EXMPLR, Q(8)=>
      OutputImg5_104_EXMPLR, Q(7)=>OutputImg5_103_EXMPLR, Q(6)=>
      OutputImg5_102_EXMPLR, Q(5)=>OutputImg5_101_EXMPLR, Q(4)=>
      OutputImg5_100_EXMPLR, Q(3)=>OutputImg5_99_EXMPLR, Q(2)=>
      OutputImg5_98_EXMPLR, Q(1)=>OutputImg5_97_EXMPLR, Q(0)=>
      OutputImg5_96_EXMPLR);
   loop3_7_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_143_EXMPLR, D(14)=>OutputImg0_142_EXMPLR, D(13)=>
      OutputImg0_141_EXMPLR, D(12)=>OutputImg0_140_EXMPLR, D(11)=>
      OutputImg0_139_EXMPLR, D(10)=>OutputImg0_138_EXMPLR, D(9)=>
      OutputImg0_137_EXMPLR, D(8)=>OutputImg0_136_EXMPLR, D(7)=>
      OutputImg0_135_EXMPLR, D(6)=>OutputImg0_134_EXMPLR, D(5)=>
      OutputImg0_133_EXMPLR, D(4)=>OutputImg0_132_EXMPLR, D(3)=>
      OutputImg0_131_EXMPLR, D(2)=>OutputImg0_130_EXMPLR, D(1)=>
      OutputImg0_129_EXMPLR, D(0)=>OutputImg0_128_EXMPLR, EN=>nx23678, F(15)
      =>ImgReg0IN_127, F(14)=>ImgReg0IN_126, F(13)=>ImgReg0IN_125, F(12)=>
      ImgReg0IN_124, F(11)=>ImgReg0IN_123, F(10)=>ImgReg0IN_122, F(9)=>
      ImgReg0IN_121, F(8)=>ImgReg0IN_120, F(7)=>ImgReg0IN_119, F(6)=>
      ImgReg0IN_118, F(5)=>ImgReg0IN_117, F(4)=>ImgReg0IN_116, F(3)=>
      ImgReg0IN_115, F(2)=>ImgReg0IN_114, F(1)=>ImgReg0IN_113, F(0)=>
      ImgReg0IN_112);
   loop3_7_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_143_EXMPLR, D(14)=>OutputImg1_142_EXMPLR, D(13)=>
      OutputImg1_141_EXMPLR, D(12)=>OutputImg1_140_EXMPLR, D(11)=>
      OutputImg1_139_EXMPLR, D(10)=>OutputImg1_138_EXMPLR, D(9)=>
      OutputImg1_137_EXMPLR, D(8)=>OutputImg1_136_EXMPLR, D(7)=>
      OutputImg1_135_EXMPLR, D(6)=>OutputImg1_134_EXMPLR, D(5)=>
      OutputImg1_133_EXMPLR, D(4)=>OutputImg1_132_EXMPLR, D(3)=>
      OutputImg1_131_EXMPLR, D(2)=>OutputImg1_130_EXMPLR, D(1)=>
      OutputImg1_129_EXMPLR, D(0)=>OutputImg1_128_EXMPLR, EN=>nx23678, F(15)
      =>ImgReg1IN_127, F(14)=>ImgReg1IN_126, F(13)=>ImgReg1IN_125, F(12)=>
      ImgReg1IN_124, F(11)=>ImgReg1IN_123, F(10)=>ImgReg1IN_122, F(9)=>
      ImgReg1IN_121, F(8)=>ImgReg1IN_120, F(7)=>ImgReg1IN_119, F(6)=>
      ImgReg1IN_118, F(5)=>ImgReg1IN_117, F(4)=>ImgReg1IN_116, F(3)=>
      ImgReg1IN_115, F(2)=>ImgReg1IN_114, F(1)=>ImgReg1IN_113, F(0)=>
      ImgReg1IN_112);
   loop3_7_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_143_EXMPLR, D(14)=>OutputImg2_142_EXMPLR, D(13)=>
      OutputImg2_141_EXMPLR, D(12)=>OutputImg2_140_EXMPLR, D(11)=>
      OutputImg2_139_EXMPLR, D(10)=>OutputImg2_138_EXMPLR, D(9)=>
      OutputImg2_137_EXMPLR, D(8)=>OutputImg2_136_EXMPLR, D(7)=>
      OutputImg2_135_EXMPLR, D(6)=>OutputImg2_134_EXMPLR, D(5)=>
      OutputImg2_133_EXMPLR, D(4)=>OutputImg2_132_EXMPLR, D(3)=>
      OutputImg2_131_EXMPLR, D(2)=>OutputImg2_130_EXMPLR, D(1)=>
      OutputImg2_129_EXMPLR, D(0)=>OutputImg2_128_EXMPLR, EN=>nx23678, F(15)
      =>ImgReg2IN_127, F(14)=>ImgReg2IN_126, F(13)=>ImgReg2IN_125, F(12)=>
      ImgReg2IN_124, F(11)=>ImgReg2IN_123, F(10)=>ImgReg2IN_122, F(9)=>
      ImgReg2IN_121, F(8)=>ImgReg2IN_120, F(7)=>ImgReg2IN_119, F(6)=>
      ImgReg2IN_118, F(5)=>ImgReg2IN_117, F(4)=>ImgReg2IN_116, F(3)=>
      ImgReg2IN_115, F(2)=>ImgReg2IN_114, F(1)=>ImgReg2IN_113, F(0)=>
      ImgReg2IN_112);
   loop3_7_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_143_EXMPLR, D(14)=>OutputImg3_142_EXMPLR, D(13)=>
      OutputImg3_141_EXMPLR, D(12)=>OutputImg3_140_EXMPLR, D(11)=>
      OutputImg3_139_EXMPLR, D(10)=>OutputImg3_138_EXMPLR, D(9)=>
      OutputImg3_137_EXMPLR, D(8)=>OutputImg3_136_EXMPLR, D(7)=>
      OutputImg3_135_EXMPLR, D(6)=>OutputImg3_134_EXMPLR, D(5)=>
      OutputImg3_133_EXMPLR, D(4)=>OutputImg3_132_EXMPLR, D(3)=>
      OutputImg3_131_EXMPLR, D(2)=>OutputImg3_130_EXMPLR, D(1)=>
      OutputImg3_129_EXMPLR, D(0)=>OutputImg3_128_EXMPLR, EN=>nx23678, F(15)
      =>ImgReg3IN_127, F(14)=>ImgReg3IN_126, F(13)=>ImgReg3IN_125, F(12)=>
      ImgReg3IN_124, F(11)=>ImgReg3IN_123, F(10)=>ImgReg3IN_122, F(9)=>
      ImgReg3IN_121, F(8)=>ImgReg3IN_120, F(7)=>ImgReg3IN_119, F(6)=>
      ImgReg3IN_118, F(5)=>ImgReg3IN_117, F(4)=>ImgReg3IN_116, F(3)=>
      ImgReg3IN_115, F(2)=>ImgReg3IN_114, F(1)=>ImgReg3IN_113, F(0)=>
      ImgReg3IN_112);
   loop3_7_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_143_EXMPLR, D(14)=>OutputImg4_142_EXMPLR, D(13)=>
      OutputImg4_141_EXMPLR, D(12)=>OutputImg4_140_EXMPLR, D(11)=>
      OutputImg4_139_EXMPLR, D(10)=>OutputImg4_138_EXMPLR, D(9)=>
      OutputImg4_137_EXMPLR, D(8)=>OutputImg4_136_EXMPLR, D(7)=>
      OutputImg4_135_EXMPLR, D(6)=>OutputImg4_134_EXMPLR, D(5)=>
      OutputImg4_133_EXMPLR, D(4)=>OutputImg4_132_EXMPLR, D(3)=>
      OutputImg4_131_EXMPLR, D(2)=>OutputImg4_130_EXMPLR, D(1)=>
      OutputImg4_129_EXMPLR, D(0)=>OutputImg4_128_EXMPLR, EN=>nx23678, F(15)
      =>ImgReg4IN_127, F(14)=>ImgReg4IN_126, F(13)=>ImgReg4IN_125, F(12)=>
      ImgReg4IN_124, F(11)=>ImgReg4IN_123, F(10)=>ImgReg4IN_122, F(9)=>
      ImgReg4IN_121, F(8)=>ImgReg4IN_120, F(7)=>ImgReg4IN_119, F(6)=>
      ImgReg4IN_118, F(5)=>ImgReg4IN_117, F(4)=>ImgReg4IN_116, F(3)=>
      ImgReg4IN_115, F(2)=>ImgReg4IN_114, F(1)=>ImgReg4IN_113, F(0)=>
      ImgReg4IN_112);
   loop3_7_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_143_EXMPLR, D(14)=>OutputImg5_142_EXMPLR, D(13)=>
      OutputImg5_141_EXMPLR, D(12)=>OutputImg5_140_EXMPLR, D(11)=>
      OutputImg5_139_EXMPLR, D(10)=>OutputImg5_138_EXMPLR, D(9)=>
      OutputImg5_137_EXMPLR, D(8)=>OutputImg5_136_EXMPLR, D(7)=>
      OutputImg5_135_EXMPLR, D(6)=>OutputImg5_134_EXMPLR, D(5)=>
      OutputImg5_133_EXMPLR, D(4)=>OutputImg5_132_EXMPLR, D(3)=>
      OutputImg5_131_EXMPLR, D(2)=>OutputImg5_130_EXMPLR, D(1)=>
      OutputImg5_129_EXMPLR, D(0)=>OutputImg5_128_EXMPLR, EN=>nx23678, F(15)
      =>ImgReg5IN_127, F(14)=>ImgReg5IN_126, F(13)=>ImgReg5IN_125, F(12)=>
      ImgReg5IN_124, F(11)=>ImgReg5IN_123, F(10)=>ImgReg5IN_122, F(9)=>
      ImgReg5IN_121, F(8)=>ImgReg5IN_120, F(7)=>ImgReg5IN_119, F(6)=>
      ImgReg5IN_118, F(5)=>ImgReg5IN_117, F(4)=>ImgReg5IN_116, F(3)=>
      ImgReg5IN_115, F(2)=>ImgReg5IN_114, F(1)=>ImgReg5IN_113, F(0)=>
      ImgReg5IN_112);
   loop3_7_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(127), D(14)
      =>DATA(126), D(13)=>DATA(125), D(12)=>DATA(124), D(11)=>DATA(123), 
      D(10)=>DATA(122), D(9)=>DATA(121), D(8)=>DATA(120), D(7)=>DATA(119), 
      D(6)=>DATA(118), D(5)=>DATA(117), D(4)=>DATA(116), D(3)=>DATA(115), 
      D(2)=>DATA(114), D(1)=>DATA(113), D(0)=>DATA(112), EN=>nx23656, F(15)
      =>ImgReg0IN_127, F(14)=>ImgReg0IN_126, F(13)=>ImgReg0IN_125, F(12)=>
      ImgReg0IN_124, F(11)=>ImgReg0IN_123, F(10)=>ImgReg0IN_122, F(9)=>
      ImgReg0IN_121, F(8)=>ImgReg0IN_120, F(7)=>ImgReg0IN_119, F(6)=>
      ImgReg0IN_118, F(5)=>ImgReg0IN_117, F(4)=>ImgReg0IN_116, F(3)=>
      ImgReg0IN_115, F(2)=>ImgReg0IN_114, F(1)=>ImgReg0IN_113, F(0)=>
      ImgReg0IN_112);
   loop3_7_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(127), D(14)
      =>DATA(126), D(13)=>DATA(125), D(12)=>DATA(124), D(11)=>DATA(123), 
      D(10)=>DATA(122), D(9)=>DATA(121), D(8)=>DATA(120), D(7)=>DATA(119), 
      D(6)=>DATA(118), D(5)=>DATA(117), D(4)=>DATA(116), D(3)=>DATA(115), 
      D(2)=>DATA(114), D(1)=>DATA(113), D(0)=>DATA(112), EN=>nx23644, F(15)
      =>ImgReg1IN_127, F(14)=>ImgReg1IN_126, F(13)=>ImgReg1IN_125, F(12)=>
      ImgReg1IN_124, F(11)=>ImgReg1IN_123, F(10)=>ImgReg1IN_122, F(9)=>
      ImgReg1IN_121, F(8)=>ImgReg1IN_120, F(7)=>ImgReg1IN_119, F(6)=>
      ImgReg1IN_118, F(5)=>ImgReg1IN_117, F(4)=>ImgReg1IN_116, F(3)=>
      ImgReg1IN_115, F(2)=>ImgReg1IN_114, F(1)=>ImgReg1IN_113, F(0)=>
      ImgReg1IN_112);
   loop3_7_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(127), D(14)
      =>DATA(126), D(13)=>DATA(125), D(12)=>DATA(124), D(11)=>DATA(123), 
      D(10)=>DATA(122), D(9)=>DATA(121), D(8)=>DATA(120), D(7)=>DATA(119), 
      D(6)=>DATA(118), D(5)=>DATA(117), D(4)=>DATA(116), D(3)=>DATA(115), 
      D(2)=>DATA(114), D(1)=>DATA(113), D(0)=>DATA(112), EN=>nx23632, F(15)
      =>ImgReg2IN_127, F(14)=>ImgReg2IN_126, F(13)=>ImgReg2IN_125, F(12)=>
      ImgReg2IN_124, F(11)=>ImgReg2IN_123, F(10)=>ImgReg2IN_122, F(9)=>
      ImgReg2IN_121, F(8)=>ImgReg2IN_120, F(7)=>ImgReg2IN_119, F(6)=>
      ImgReg2IN_118, F(5)=>ImgReg2IN_117, F(4)=>ImgReg2IN_116, F(3)=>
      ImgReg2IN_115, F(2)=>ImgReg2IN_114, F(1)=>ImgReg2IN_113, F(0)=>
      ImgReg2IN_112);
   loop3_7_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(127), D(14)
      =>DATA(126), D(13)=>DATA(125), D(12)=>DATA(124), D(11)=>DATA(123), 
      D(10)=>DATA(122), D(9)=>DATA(121), D(8)=>DATA(120), D(7)=>DATA(119), 
      D(6)=>DATA(118), D(5)=>DATA(117), D(4)=>DATA(116), D(3)=>DATA(115), 
      D(2)=>DATA(114), D(1)=>DATA(113), D(0)=>DATA(112), EN=>nx23620, F(15)
      =>ImgReg3IN_127, F(14)=>ImgReg3IN_126, F(13)=>ImgReg3IN_125, F(12)=>
      ImgReg3IN_124, F(11)=>ImgReg3IN_123, F(10)=>ImgReg3IN_122, F(9)=>
      ImgReg3IN_121, F(8)=>ImgReg3IN_120, F(7)=>ImgReg3IN_119, F(6)=>
      ImgReg3IN_118, F(5)=>ImgReg3IN_117, F(4)=>ImgReg3IN_116, F(3)=>
      ImgReg3IN_115, F(2)=>ImgReg3IN_114, F(1)=>ImgReg3IN_113, F(0)=>
      ImgReg3IN_112);
   loop3_7_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(127), D(14)
      =>DATA(126), D(13)=>DATA(125), D(12)=>DATA(124), D(11)=>DATA(123), 
      D(10)=>DATA(122), D(9)=>DATA(121), D(8)=>DATA(120), D(7)=>DATA(119), 
      D(6)=>DATA(118), D(5)=>DATA(117), D(4)=>DATA(116), D(3)=>DATA(115), 
      D(2)=>DATA(114), D(1)=>DATA(113), D(0)=>DATA(112), EN=>nx23608, F(15)
      =>ImgReg4IN_127, F(14)=>ImgReg4IN_126, F(13)=>ImgReg4IN_125, F(12)=>
      ImgReg4IN_124, F(11)=>ImgReg4IN_123, F(10)=>ImgReg4IN_122, F(9)=>
      ImgReg4IN_121, F(8)=>ImgReg4IN_120, F(7)=>ImgReg4IN_119, F(6)=>
      ImgReg4IN_118, F(5)=>ImgReg4IN_117, F(4)=>ImgReg4IN_116, F(3)=>
      ImgReg4IN_115, F(2)=>ImgReg4IN_114, F(1)=>ImgReg4IN_113, F(0)=>
      ImgReg4IN_112);
   loop3_7_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(127), D(14)
      =>DATA(126), D(13)=>DATA(125), D(12)=>DATA(124), D(11)=>DATA(123), 
      D(10)=>DATA(122), D(9)=>DATA(121), D(8)=>DATA(120), D(7)=>DATA(119), 
      D(6)=>DATA(118), D(5)=>DATA(117), D(4)=>DATA(116), D(3)=>DATA(115), 
      D(2)=>DATA(114), D(1)=>DATA(113), D(0)=>DATA(112), EN=>nx23596, F(15)
      =>ImgReg5IN_127, F(14)=>ImgReg5IN_126, F(13)=>ImgReg5IN_125, F(12)=>
      ImgReg5IN_124, F(11)=>ImgReg5IN_123, F(10)=>ImgReg5IN_122, F(9)=>
      ImgReg5IN_121, F(8)=>ImgReg5IN_120, F(7)=>ImgReg5IN_119, F(6)=>
      ImgReg5IN_118, F(5)=>ImgReg5IN_117, F(4)=>ImgReg5IN_116, F(3)=>
      ImgReg5IN_115, F(2)=>ImgReg5IN_114, F(1)=>ImgReg5IN_113, F(0)=>
      ImgReg5IN_112);
   loop3_7_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_127_EXMPLR, D(14)=>OutputImg1_126_EXMPLR, D(13)=>
      OutputImg1_125_EXMPLR, D(12)=>OutputImg1_124_EXMPLR, D(11)=>
      OutputImg1_123_EXMPLR, D(10)=>OutputImg1_122_EXMPLR, D(9)=>
      OutputImg1_121_EXMPLR, D(8)=>OutputImg1_120_EXMPLR, D(7)=>
      OutputImg1_119_EXMPLR, D(6)=>OutputImg1_118_EXMPLR, D(5)=>
      OutputImg1_117_EXMPLR, D(4)=>OutputImg1_116_EXMPLR, D(3)=>
      OutputImg1_115_EXMPLR, D(2)=>OutputImg1_114_EXMPLR, D(1)=>
      OutputImg1_113_EXMPLR, D(0)=>OutputImg1_112_EXMPLR, EN=>nx23796, F(15)
      =>ImgReg0IN_127, F(14)=>ImgReg0IN_126, F(13)=>ImgReg0IN_125, F(12)=>
      ImgReg0IN_124, F(11)=>ImgReg0IN_123, F(10)=>ImgReg0IN_122, F(9)=>
      ImgReg0IN_121, F(8)=>ImgReg0IN_120, F(7)=>ImgReg0IN_119, F(6)=>
      ImgReg0IN_118, F(5)=>ImgReg0IN_117, F(4)=>ImgReg0IN_116, F(3)=>
      ImgReg0IN_115, F(2)=>ImgReg0IN_114, F(1)=>ImgReg0IN_113, F(0)=>
      ImgReg0IN_112);
   loop3_7_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_127_EXMPLR, D(14)=>OutputImg2_126_EXMPLR, D(13)=>
      OutputImg2_125_EXMPLR, D(12)=>OutputImg2_124_EXMPLR, D(11)=>
      OutputImg2_123_EXMPLR, D(10)=>OutputImg2_122_EXMPLR, D(9)=>
      OutputImg2_121_EXMPLR, D(8)=>OutputImg2_120_EXMPLR, D(7)=>
      OutputImg2_119_EXMPLR, D(6)=>OutputImg2_118_EXMPLR, D(5)=>
      OutputImg2_117_EXMPLR, D(4)=>OutputImg2_116_EXMPLR, D(3)=>
      OutputImg2_115_EXMPLR, D(2)=>OutputImg2_114_EXMPLR, D(1)=>
      OutputImg2_113_EXMPLR, D(0)=>OutputImg2_112_EXMPLR, EN=>nx23796, F(15)
      =>ImgReg1IN_127, F(14)=>ImgReg1IN_126, F(13)=>ImgReg1IN_125, F(12)=>
      ImgReg1IN_124, F(11)=>ImgReg1IN_123, F(10)=>ImgReg1IN_122, F(9)=>
      ImgReg1IN_121, F(8)=>ImgReg1IN_120, F(7)=>ImgReg1IN_119, F(6)=>
      ImgReg1IN_118, F(5)=>ImgReg1IN_117, F(4)=>ImgReg1IN_116, F(3)=>
      ImgReg1IN_115, F(2)=>ImgReg1IN_114, F(1)=>ImgReg1IN_113, F(0)=>
      ImgReg1IN_112);
   loop3_7_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_127_EXMPLR, D(14)=>OutputImg3_126_EXMPLR, D(13)=>
      OutputImg3_125_EXMPLR, D(12)=>OutputImg3_124_EXMPLR, D(11)=>
      OutputImg3_123_EXMPLR, D(10)=>OutputImg3_122_EXMPLR, D(9)=>
      OutputImg3_121_EXMPLR, D(8)=>OutputImg3_120_EXMPLR, D(7)=>
      OutputImg3_119_EXMPLR, D(6)=>OutputImg3_118_EXMPLR, D(5)=>
      OutputImg3_117_EXMPLR, D(4)=>OutputImg3_116_EXMPLR, D(3)=>
      OutputImg3_115_EXMPLR, D(2)=>OutputImg3_114_EXMPLR, D(1)=>
      OutputImg3_113_EXMPLR, D(0)=>OutputImg3_112_EXMPLR, EN=>nx23796, F(15)
      =>ImgReg2IN_127, F(14)=>ImgReg2IN_126, F(13)=>ImgReg2IN_125, F(12)=>
      ImgReg2IN_124, F(11)=>ImgReg2IN_123, F(10)=>ImgReg2IN_122, F(9)=>
      ImgReg2IN_121, F(8)=>ImgReg2IN_120, F(7)=>ImgReg2IN_119, F(6)=>
      ImgReg2IN_118, F(5)=>ImgReg2IN_117, F(4)=>ImgReg2IN_116, F(3)=>
      ImgReg2IN_115, F(2)=>ImgReg2IN_114, F(1)=>ImgReg2IN_113, F(0)=>
      ImgReg2IN_112);
   loop3_7_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_127_EXMPLR, D(14)=>OutputImg4_126_EXMPLR, D(13)=>
      OutputImg4_125_EXMPLR, D(12)=>OutputImg4_124_EXMPLR, D(11)=>
      OutputImg4_123_EXMPLR, D(10)=>OutputImg4_122_EXMPLR, D(9)=>
      OutputImg4_121_EXMPLR, D(8)=>OutputImg4_120_EXMPLR, D(7)=>
      OutputImg4_119_EXMPLR, D(6)=>OutputImg4_118_EXMPLR, D(5)=>
      OutputImg4_117_EXMPLR, D(4)=>OutputImg4_116_EXMPLR, D(3)=>
      OutputImg4_115_EXMPLR, D(2)=>OutputImg4_114_EXMPLR, D(1)=>
      OutputImg4_113_EXMPLR, D(0)=>OutputImg4_112_EXMPLR, EN=>nx23796, F(15)
      =>ImgReg3IN_127, F(14)=>ImgReg3IN_126, F(13)=>ImgReg3IN_125, F(12)=>
      ImgReg3IN_124, F(11)=>ImgReg3IN_123, F(10)=>ImgReg3IN_122, F(9)=>
      ImgReg3IN_121, F(8)=>ImgReg3IN_120, F(7)=>ImgReg3IN_119, F(6)=>
      ImgReg3IN_118, F(5)=>ImgReg3IN_117, F(4)=>ImgReg3IN_116, F(3)=>
      ImgReg3IN_115, F(2)=>ImgReg3IN_114, F(1)=>ImgReg3IN_113, F(0)=>
      ImgReg3IN_112);
   loop3_7_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_127_EXMPLR, D(14)=>OutputImg5_126_EXMPLR, D(13)=>
      OutputImg5_125_EXMPLR, D(12)=>OutputImg5_124_EXMPLR, D(11)=>
      OutputImg5_123_EXMPLR, D(10)=>OutputImg5_122_EXMPLR, D(9)=>
      OutputImg5_121_EXMPLR, D(8)=>OutputImg5_120_EXMPLR, D(7)=>
      OutputImg5_119_EXMPLR, D(6)=>OutputImg5_118_EXMPLR, D(5)=>
      OutputImg5_117_EXMPLR, D(4)=>OutputImg5_116_EXMPLR, D(3)=>
      OutputImg5_115_EXMPLR, D(2)=>OutputImg5_114_EXMPLR, D(1)=>
      OutputImg5_113_EXMPLR, D(0)=>OutputImg5_112_EXMPLR, EN=>nx23796, F(15)
      =>ImgReg4IN_127, F(14)=>ImgReg4IN_126, F(13)=>ImgReg4IN_125, F(12)=>
      ImgReg4IN_124, F(11)=>ImgReg4IN_123, F(10)=>ImgReg4IN_122, F(9)=>
      ImgReg4IN_121, F(8)=>ImgReg4IN_120, F(7)=>ImgReg4IN_119, F(6)=>
      ImgReg4IN_118, F(5)=>ImgReg4IN_117, F(4)=>ImgReg4IN_116, F(3)=>
      ImgReg4IN_115, F(2)=>ImgReg4IN_114, F(1)=>ImgReg4IN_113, F(0)=>
      ImgReg4IN_112);
   loop3_7_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_127, D(14)=>
      ImgReg0IN_126, D(13)=>ImgReg0IN_125, D(12)=>ImgReg0IN_124, D(11)=>
      ImgReg0IN_123, D(10)=>ImgReg0IN_122, D(9)=>ImgReg0IN_121, D(8)=>
      ImgReg0IN_120, D(7)=>ImgReg0IN_119, D(6)=>ImgReg0IN_118, D(5)=>
      ImgReg0IN_117, D(4)=>ImgReg0IN_116, D(3)=>ImgReg0IN_115, D(2)=>
      ImgReg0IN_114, D(1)=>ImgReg0IN_113, D(0)=>ImgReg0IN_112, CLK=>nx23870, 
      RST=>RST, EN=>nx23720, Q(15)=>OutputImg0_127_EXMPLR, Q(14)=>
      OutputImg0_126_EXMPLR, Q(13)=>OutputImg0_125_EXMPLR, Q(12)=>
      OutputImg0_124_EXMPLR, Q(11)=>OutputImg0_123_EXMPLR, Q(10)=>
      OutputImg0_122_EXMPLR, Q(9)=>OutputImg0_121_EXMPLR, Q(8)=>
      OutputImg0_120_EXMPLR, Q(7)=>OutputImg0_119_EXMPLR, Q(6)=>
      OutputImg0_118_EXMPLR, Q(5)=>OutputImg0_117_EXMPLR, Q(4)=>
      OutputImg0_116_EXMPLR, Q(3)=>OutputImg0_115_EXMPLR, Q(2)=>
      OutputImg0_114_EXMPLR, Q(1)=>OutputImg0_113_EXMPLR, Q(0)=>
      OutputImg0_112_EXMPLR);
   loop3_7_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_127, D(14)=>
      ImgReg1IN_126, D(13)=>ImgReg1IN_125, D(12)=>ImgReg1IN_124, D(11)=>
      ImgReg1IN_123, D(10)=>ImgReg1IN_122, D(9)=>ImgReg1IN_121, D(8)=>
      ImgReg1IN_120, D(7)=>ImgReg1IN_119, D(6)=>ImgReg1IN_118, D(5)=>
      ImgReg1IN_117, D(4)=>ImgReg1IN_116, D(3)=>ImgReg1IN_115, D(2)=>
      ImgReg1IN_114, D(1)=>ImgReg1IN_113, D(0)=>ImgReg1IN_112, CLK=>nx23872, 
      RST=>RST, EN=>nx23730, Q(15)=>OutputImg1_127_EXMPLR, Q(14)=>
      OutputImg1_126_EXMPLR, Q(13)=>OutputImg1_125_EXMPLR, Q(12)=>
      OutputImg1_124_EXMPLR, Q(11)=>OutputImg1_123_EXMPLR, Q(10)=>
      OutputImg1_122_EXMPLR, Q(9)=>OutputImg1_121_EXMPLR, Q(8)=>
      OutputImg1_120_EXMPLR, Q(7)=>OutputImg1_119_EXMPLR, Q(6)=>
      OutputImg1_118_EXMPLR, Q(5)=>OutputImg1_117_EXMPLR, Q(4)=>
      OutputImg1_116_EXMPLR, Q(3)=>OutputImg1_115_EXMPLR, Q(2)=>
      OutputImg1_114_EXMPLR, Q(1)=>OutputImg1_113_EXMPLR, Q(0)=>
      OutputImg1_112_EXMPLR);
   loop3_7_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_127, D(14)=>
      ImgReg2IN_126, D(13)=>ImgReg2IN_125, D(12)=>ImgReg2IN_124, D(11)=>
      ImgReg2IN_123, D(10)=>ImgReg2IN_122, D(9)=>ImgReg2IN_121, D(8)=>
      ImgReg2IN_120, D(7)=>ImgReg2IN_119, D(6)=>ImgReg2IN_118, D(5)=>
      ImgReg2IN_117, D(4)=>ImgReg2IN_116, D(3)=>ImgReg2IN_115, D(2)=>
      ImgReg2IN_114, D(1)=>ImgReg2IN_113, D(0)=>ImgReg2IN_112, CLK=>nx23872, 
      RST=>RST, EN=>nx23740, Q(15)=>OutputImg2_127_EXMPLR, Q(14)=>
      OutputImg2_126_EXMPLR, Q(13)=>OutputImg2_125_EXMPLR, Q(12)=>
      OutputImg2_124_EXMPLR, Q(11)=>OutputImg2_123_EXMPLR, Q(10)=>
      OutputImg2_122_EXMPLR, Q(9)=>OutputImg2_121_EXMPLR, Q(8)=>
      OutputImg2_120_EXMPLR, Q(7)=>OutputImg2_119_EXMPLR, Q(6)=>
      OutputImg2_118_EXMPLR, Q(5)=>OutputImg2_117_EXMPLR, Q(4)=>
      OutputImg2_116_EXMPLR, Q(3)=>OutputImg2_115_EXMPLR, Q(2)=>
      OutputImg2_114_EXMPLR, Q(1)=>OutputImg2_113_EXMPLR, Q(0)=>
      OutputImg2_112_EXMPLR);
   loop3_7_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_127, D(14)=>
      ImgReg3IN_126, D(13)=>ImgReg3IN_125, D(12)=>ImgReg3IN_124, D(11)=>
      ImgReg3IN_123, D(10)=>ImgReg3IN_122, D(9)=>ImgReg3IN_121, D(8)=>
      ImgReg3IN_120, D(7)=>ImgReg3IN_119, D(6)=>ImgReg3IN_118, D(5)=>
      ImgReg3IN_117, D(4)=>ImgReg3IN_116, D(3)=>ImgReg3IN_115, D(2)=>
      ImgReg3IN_114, D(1)=>ImgReg3IN_113, D(0)=>ImgReg3IN_112, CLK=>nx23874, 
      RST=>RST, EN=>nx23750, Q(15)=>OutputImg3_127_EXMPLR, Q(14)=>
      OutputImg3_126_EXMPLR, Q(13)=>OutputImg3_125_EXMPLR, Q(12)=>
      OutputImg3_124_EXMPLR, Q(11)=>OutputImg3_123_EXMPLR, Q(10)=>
      OutputImg3_122_EXMPLR, Q(9)=>OutputImg3_121_EXMPLR, Q(8)=>
      OutputImg3_120_EXMPLR, Q(7)=>OutputImg3_119_EXMPLR, Q(6)=>
      OutputImg3_118_EXMPLR, Q(5)=>OutputImg3_117_EXMPLR, Q(4)=>
      OutputImg3_116_EXMPLR, Q(3)=>OutputImg3_115_EXMPLR, Q(2)=>
      OutputImg3_114_EXMPLR, Q(1)=>OutputImg3_113_EXMPLR, Q(0)=>
      OutputImg3_112_EXMPLR);
   loop3_7_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_127, D(14)=>
      ImgReg4IN_126, D(13)=>ImgReg4IN_125, D(12)=>ImgReg4IN_124, D(11)=>
      ImgReg4IN_123, D(10)=>ImgReg4IN_122, D(9)=>ImgReg4IN_121, D(8)=>
      ImgReg4IN_120, D(7)=>ImgReg4IN_119, D(6)=>ImgReg4IN_118, D(5)=>
      ImgReg4IN_117, D(4)=>ImgReg4IN_116, D(3)=>ImgReg4IN_115, D(2)=>
      ImgReg4IN_114, D(1)=>ImgReg4IN_113, D(0)=>ImgReg4IN_112, CLK=>nx23874, 
      RST=>RST, EN=>nx23760, Q(15)=>OutputImg4_127_EXMPLR, Q(14)=>
      OutputImg4_126_EXMPLR, Q(13)=>OutputImg4_125_EXMPLR, Q(12)=>
      OutputImg4_124_EXMPLR, Q(11)=>OutputImg4_123_EXMPLR, Q(10)=>
      OutputImg4_122_EXMPLR, Q(9)=>OutputImg4_121_EXMPLR, Q(8)=>
      OutputImg4_120_EXMPLR, Q(7)=>OutputImg4_119_EXMPLR, Q(6)=>
      OutputImg4_118_EXMPLR, Q(5)=>OutputImg4_117_EXMPLR, Q(4)=>
      OutputImg4_116_EXMPLR, Q(3)=>OutputImg4_115_EXMPLR, Q(2)=>
      OutputImg4_114_EXMPLR, Q(1)=>OutputImg4_113_EXMPLR, Q(0)=>
      OutputImg4_112_EXMPLR);
   loop3_7_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_127, D(14)=>
      ImgReg5IN_126, D(13)=>ImgReg5IN_125, D(12)=>ImgReg5IN_124, D(11)=>
      ImgReg5IN_123, D(10)=>ImgReg5IN_122, D(9)=>ImgReg5IN_121, D(8)=>
      ImgReg5IN_120, D(7)=>ImgReg5IN_119, D(6)=>ImgReg5IN_118, D(5)=>
      ImgReg5IN_117, D(4)=>ImgReg5IN_116, D(3)=>ImgReg5IN_115, D(2)=>
      ImgReg5IN_114, D(1)=>ImgReg5IN_113, D(0)=>ImgReg5IN_112, CLK=>nx23876, 
      RST=>RST, EN=>nx23770, Q(15)=>OutputImg5_127_EXMPLR, Q(14)=>
      OutputImg5_126_EXMPLR, Q(13)=>OutputImg5_125_EXMPLR, Q(12)=>
      OutputImg5_124_EXMPLR, Q(11)=>OutputImg5_123_EXMPLR, Q(10)=>
      OutputImg5_122_EXMPLR, Q(9)=>OutputImg5_121_EXMPLR, Q(8)=>
      OutputImg5_120_EXMPLR, Q(7)=>OutputImg5_119_EXMPLR, Q(6)=>
      OutputImg5_118_EXMPLR, Q(5)=>OutputImg5_117_EXMPLR, Q(4)=>
      OutputImg5_116_EXMPLR, Q(3)=>OutputImg5_115_EXMPLR, Q(2)=>
      OutputImg5_114_EXMPLR, Q(1)=>OutputImg5_113_EXMPLR, Q(0)=>
      OutputImg5_112_EXMPLR);
   loop3_8_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_159_EXMPLR, D(14)=>OutputImg0_158_EXMPLR, D(13)=>
      OutputImg0_157_EXMPLR, D(12)=>OutputImg0_156_EXMPLR, D(11)=>
      OutputImg0_155_EXMPLR, D(10)=>OutputImg0_154_EXMPLR, D(9)=>
      OutputImg0_153_EXMPLR, D(8)=>OutputImg0_152_EXMPLR, D(7)=>
      OutputImg0_151_EXMPLR, D(6)=>OutputImg0_150_EXMPLR, D(5)=>
      OutputImg0_149_EXMPLR, D(4)=>OutputImg0_148_EXMPLR, D(3)=>
      OutputImg0_147_EXMPLR, D(2)=>OutputImg0_146_EXMPLR, D(1)=>
      OutputImg0_145_EXMPLR, D(0)=>OutputImg0_144_EXMPLR, EN=>nx23678, F(15)
      =>ImgReg0IN_143, F(14)=>ImgReg0IN_142, F(13)=>ImgReg0IN_141, F(12)=>
      ImgReg0IN_140, F(11)=>ImgReg0IN_139, F(10)=>ImgReg0IN_138, F(9)=>
      ImgReg0IN_137, F(8)=>ImgReg0IN_136, F(7)=>ImgReg0IN_135, F(6)=>
      ImgReg0IN_134, F(5)=>ImgReg0IN_133, F(4)=>ImgReg0IN_132, F(3)=>
      ImgReg0IN_131, F(2)=>ImgReg0IN_130, F(1)=>ImgReg0IN_129, F(0)=>
      ImgReg0IN_128);
   loop3_8_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_159_EXMPLR, D(14)=>OutputImg1_158_EXMPLR, D(13)=>
      OutputImg1_157_EXMPLR, D(12)=>OutputImg1_156_EXMPLR, D(11)=>
      OutputImg1_155_EXMPLR, D(10)=>OutputImg1_154_EXMPLR, D(9)=>
      OutputImg1_153_EXMPLR, D(8)=>OutputImg1_152_EXMPLR, D(7)=>
      OutputImg1_151_EXMPLR, D(6)=>OutputImg1_150_EXMPLR, D(5)=>
      OutputImg1_149_EXMPLR, D(4)=>OutputImg1_148_EXMPLR, D(3)=>
      OutputImg1_147_EXMPLR, D(2)=>OutputImg1_146_EXMPLR, D(1)=>
      OutputImg1_145_EXMPLR, D(0)=>OutputImg1_144_EXMPLR, EN=>nx23680, F(15)
      =>ImgReg1IN_143, F(14)=>ImgReg1IN_142, F(13)=>ImgReg1IN_141, F(12)=>
      ImgReg1IN_140, F(11)=>ImgReg1IN_139, F(10)=>ImgReg1IN_138, F(9)=>
      ImgReg1IN_137, F(8)=>ImgReg1IN_136, F(7)=>ImgReg1IN_135, F(6)=>
      ImgReg1IN_134, F(5)=>ImgReg1IN_133, F(4)=>ImgReg1IN_132, F(3)=>
      ImgReg1IN_131, F(2)=>ImgReg1IN_130, F(1)=>ImgReg1IN_129, F(0)=>
      ImgReg1IN_128);
   loop3_8_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_159_EXMPLR, D(14)=>OutputImg2_158_EXMPLR, D(13)=>
      OutputImg2_157_EXMPLR, D(12)=>OutputImg2_156_EXMPLR, D(11)=>
      OutputImg2_155_EXMPLR, D(10)=>OutputImg2_154_EXMPLR, D(9)=>
      OutputImg2_153_EXMPLR, D(8)=>OutputImg2_152_EXMPLR, D(7)=>
      OutputImg2_151_EXMPLR, D(6)=>OutputImg2_150_EXMPLR, D(5)=>
      OutputImg2_149_EXMPLR, D(4)=>OutputImg2_148_EXMPLR, D(3)=>
      OutputImg2_147_EXMPLR, D(2)=>OutputImg2_146_EXMPLR, D(1)=>
      OutputImg2_145_EXMPLR, D(0)=>OutputImg2_144_EXMPLR, EN=>nx23680, F(15)
      =>ImgReg2IN_143, F(14)=>ImgReg2IN_142, F(13)=>ImgReg2IN_141, F(12)=>
      ImgReg2IN_140, F(11)=>ImgReg2IN_139, F(10)=>ImgReg2IN_138, F(9)=>
      ImgReg2IN_137, F(8)=>ImgReg2IN_136, F(7)=>ImgReg2IN_135, F(6)=>
      ImgReg2IN_134, F(5)=>ImgReg2IN_133, F(4)=>ImgReg2IN_132, F(3)=>
      ImgReg2IN_131, F(2)=>ImgReg2IN_130, F(1)=>ImgReg2IN_129, F(0)=>
      ImgReg2IN_128);
   loop3_8_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_159_EXMPLR, D(14)=>OutputImg3_158_EXMPLR, D(13)=>
      OutputImg3_157_EXMPLR, D(12)=>OutputImg3_156_EXMPLR, D(11)=>
      OutputImg3_155_EXMPLR, D(10)=>OutputImg3_154_EXMPLR, D(9)=>
      OutputImg3_153_EXMPLR, D(8)=>OutputImg3_152_EXMPLR, D(7)=>
      OutputImg3_151_EXMPLR, D(6)=>OutputImg3_150_EXMPLR, D(5)=>
      OutputImg3_149_EXMPLR, D(4)=>OutputImg3_148_EXMPLR, D(3)=>
      OutputImg3_147_EXMPLR, D(2)=>OutputImg3_146_EXMPLR, D(1)=>
      OutputImg3_145_EXMPLR, D(0)=>OutputImg3_144_EXMPLR, EN=>nx23680, F(15)
      =>ImgReg3IN_143, F(14)=>ImgReg3IN_142, F(13)=>ImgReg3IN_141, F(12)=>
      ImgReg3IN_140, F(11)=>ImgReg3IN_139, F(10)=>ImgReg3IN_138, F(9)=>
      ImgReg3IN_137, F(8)=>ImgReg3IN_136, F(7)=>ImgReg3IN_135, F(6)=>
      ImgReg3IN_134, F(5)=>ImgReg3IN_133, F(4)=>ImgReg3IN_132, F(3)=>
      ImgReg3IN_131, F(2)=>ImgReg3IN_130, F(1)=>ImgReg3IN_129, F(0)=>
      ImgReg3IN_128);
   loop3_8_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_159_EXMPLR, D(14)=>OutputImg4_158_EXMPLR, D(13)=>
      OutputImg4_157_EXMPLR, D(12)=>OutputImg4_156_EXMPLR, D(11)=>
      OutputImg4_155_EXMPLR, D(10)=>OutputImg4_154_EXMPLR, D(9)=>
      OutputImg4_153_EXMPLR, D(8)=>OutputImg4_152_EXMPLR, D(7)=>
      OutputImg4_151_EXMPLR, D(6)=>OutputImg4_150_EXMPLR, D(5)=>
      OutputImg4_149_EXMPLR, D(4)=>OutputImg4_148_EXMPLR, D(3)=>
      OutputImg4_147_EXMPLR, D(2)=>OutputImg4_146_EXMPLR, D(1)=>
      OutputImg4_145_EXMPLR, D(0)=>OutputImg4_144_EXMPLR, EN=>nx23680, F(15)
      =>ImgReg4IN_143, F(14)=>ImgReg4IN_142, F(13)=>ImgReg4IN_141, F(12)=>
      ImgReg4IN_140, F(11)=>ImgReg4IN_139, F(10)=>ImgReg4IN_138, F(9)=>
      ImgReg4IN_137, F(8)=>ImgReg4IN_136, F(7)=>ImgReg4IN_135, F(6)=>
      ImgReg4IN_134, F(5)=>ImgReg4IN_133, F(4)=>ImgReg4IN_132, F(3)=>
      ImgReg4IN_131, F(2)=>ImgReg4IN_130, F(1)=>ImgReg4IN_129, F(0)=>
      ImgReg4IN_128);
   loop3_8_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_159_EXMPLR, D(14)=>OutputImg5_158_EXMPLR, D(13)=>
      OutputImg5_157_EXMPLR, D(12)=>OutputImg5_156_EXMPLR, D(11)=>
      OutputImg5_155_EXMPLR, D(10)=>OutputImg5_154_EXMPLR, D(9)=>
      OutputImg5_153_EXMPLR, D(8)=>OutputImg5_152_EXMPLR, D(7)=>
      OutputImg5_151_EXMPLR, D(6)=>OutputImg5_150_EXMPLR, D(5)=>
      OutputImg5_149_EXMPLR, D(4)=>OutputImg5_148_EXMPLR, D(3)=>
      OutputImg5_147_EXMPLR, D(2)=>OutputImg5_146_EXMPLR, D(1)=>
      OutputImg5_145_EXMPLR, D(0)=>OutputImg5_144_EXMPLR, EN=>nx23680, F(15)
      =>ImgReg5IN_143, F(14)=>ImgReg5IN_142, F(13)=>ImgReg5IN_141, F(12)=>
      ImgReg5IN_140, F(11)=>ImgReg5IN_139, F(10)=>ImgReg5IN_138, F(9)=>
      ImgReg5IN_137, F(8)=>ImgReg5IN_136, F(7)=>ImgReg5IN_135, F(6)=>
      ImgReg5IN_134, F(5)=>ImgReg5IN_133, F(4)=>ImgReg5IN_132, F(3)=>
      ImgReg5IN_131, F(2)=>ImgReg5IN_130, F(1)=>ImgReg5IN_129, F(0)=>
      ImgReg5IN_128);
   loop3_8_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(143), D(14)
      =>DATA(142), D(13)=>DATA(141), D(12)=>DATA(140), D(11)=>DATA(139), 
      D(10)=>DATA(138), D(9)=>DATA(137), D(8)=>DATA(136), D(7)=>DATA(135), 
      D(6)=>DATA(134), D(5)=>DATA(133), D(4)=>DATA(132), D(3)=>DATA(131), 
      D(2)=>DATA(130), D(1)=>DATA(129), D(0)=>DATA(128), EN=>nx23656, F(15)
      =>ImgReg0IN_143, F(14)=>ImgReg0IN_142, F(13)=>ImgReg0IN_141, F(12)=>
      ImgReg0IN_140, F(11)=>ImgReg0IN_139, F(10)=>ImgReg0IN_138, F(9)=>
      ImgReg0IN_137, F(8)=>ImgReg0IN_136, F(7)=>ImgReg0IN_135, F(6)=>
      ImgReg0IN_134, F(5)=>ImgReg0IN_133, F(4)=>ImgReg0IN_132, F(3)=>
      ImgReg0IN_131, F(2)=>ImgReg0IN_130, F(1)=>ImgReg0IN_129, F(0)=>
      ImgReg0IN_128);
   loop3_8_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(143), D(14)
      =>DATA(142), D(13)=>DATA(141), D(12)=>DATA(140), D(11)=>DATA(139), 
      D(10)=>DATA(138), D(9)=>DATA(137), D(8)=>DATA(136), D(7)=>DATA(135), 
      D(6)=>DATA(134), D(5)=>DATA(133), D(4)=>DATA(132), D(3)=>DATA(131), 
      D(2)=>DATA(130), D(1)=>DATA(129), D(0)=>DATA(128), EN=>nx23644, F(15)
      =>ImgReg1IN_143, F(14)=>ImgReg1IN_142, F(13)=>ImgReg1IN_141, F(12)=>
      ImgReg1IN_140, F(11)=>ImgReg1IN_139, F(10)=>ImgReg1IN_138, F(9)=>
      ImgReg1IN_137, F(8)=>ImgReg1IN_136, F(7)=>ImgReg1IN_135, F(6)=>
      ImgReg1IN_134, F(5)=>ImgReg1IN_133, F(4)=>ImgReg1IN_132, F(3)=>
      ImgReg1IN_131, F(2)=>ImgReg1IN_130, F(1)=>ImgReg1IN_129, F(0)=>
      ImgReg1IN_128);
   loop3_8_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(143), D(14)
      =>DATA(142), D(13)=>DATA(141), D(12)=>DATA(140), D(11)=>DATA(139), 
      D(10)=>DATA(138), D(9)=>DATA(137), D(8)=>DATA(136), D(7)=>DATA(135), 
      D(6)=>DATA(134), D(5)=>DATA(133), D(4)=>DATA(132), D(3)=>DATA(131), 
      D(2)=>DATA(130), D(1)=>DATA(129), D(0)=>DATA(128), EN=>nx23632, F(15)
      =>ImgReg2IN_143, F(14)=>ImgReg2IN_142, F(13)=>ImgReg2IN_141, F(12)=>
      ImgReg2IN_140, F(11)=>ImgReg2IN_139, F(10)=>ImgReg2IN_138, F(9)=>
      ImgReg2IN_137, F(8)=>ImgReg2IN_136, F(7)=>ImgReg2IN_135, F(6)=>
      ImgReg2IN_134, F(5)=>ImgReg2IN_133, F(4)=>ImgReg2IN_132, F(3)=>
      ImgReg2IN_131, F(2)=>ImgReg2IN_130, F(1)=>ImgReg2IN_129, F(0)=>
      ImgReg2IN_128);
   loop3_8_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(143), D(14)
      =>DATA(142), D(13)=>DATA(141), D(12)=>DATA(140), D(11)=>DATA(139), 
      D(10)=>DATA(138), D(9)=>DATA(137), D(8)=>DATA(136), D(7)=>DATA(135), 
      D(6)=>DATA(134), D(5)=>DATA(133), D(4)=>DATA(132), D(3)=>DATA(131), 
      D(2)=>DATA(130), D(1)=>DATA(129), D(0)=>DATA(128), EN=>nx23620, F(15)
      =>ImgReg3IN_143, F(14)=>ImgReg3IN_142, F(13)=>ImgReg3IN_141, F(12)=>
      ImgReg3IN_140, F(11)=>ImgReg3IN_139, F(10)=>ImgReg3IN_138, F(9)=>
      ImgReg3IN_137, F(8)=>ImgReg3IN_136, F(7)=>ImgReg3IN_135, F(6)=>
      ImgReg3IN_134, F(5)=>ImgReg3IN_133, F(4)=>ImgReg3IN_132, F(3)=>
      ImgReg3IN_131, F(2)=>ImgReg3IN_130, F(1)=>ImgReg3IN_129, F(0)=>
      ImgReg3IN_128);
   loop3_8_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(143), D(14)
      =>DATA(142), D(13)=>DATA(141), D(12)=>DATA(140), D(11)=>DATA(139), 
      D(10)=>DATA(138), D(9)=>DATA(137), D(8)=>DATA(136), D(7)=>DATA(135), 
      D(6)=>DATA(134), D(5)=>DATA(133), D(4)=>DATA(132), D(3)=>DATA(131), 
      D(2)=>DATA(130), D(1)=>DATA(129), D(0)=>DATA(128), EN=>nx23608, F(15)
      =>ImgReg4IN_143, F(14)=>ImgReg4IN_142, F(13)=>ImgReg4IN_141, F(12)=>
      ImgReg4IN_140, F(11)=>ImgReg4IN_139, F(10)=>ImgReg4IN_138, F(9)=>
      ImgReg4IN_137, F(8)=>ImgReg4IN_136, F(7)=>ImgReg4IN_135, F(6)=>
      ImgReg4IN_134, F(5)=>ImgReg4IN_133, F(4)=>ImgReg4IN_132, F(3)=>
      ImgReg4IN_131, F(2)=>ImgReg4IN_130, F(1)=>ImgReg4IN_129, F(0)=>
      ImgReg4IN_128);
   loop3_8_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(143), D(14)
      =>DATA(142), D(13)=>DATA(141), D(12)=>DATA(140), D(11)=>DATA(139), 
      D(10)=>DATA(138), D(9)=>DATA(137), D(8)=>DATA(136), D(7)=>DATA(135), 
      D(6)=>DATA(134), D(5)=>DATA(133), D(4)=>DATA(132), D(3)=>DATA(131), 
      D(2)=>DATA(130), D(1)=>DATA(129), D(0)=>DATA(128), EN=>nx23596, F(15)
      =>ImgReg5IN_143, F(14)=>ImgReg5IN_142, F(13)=>ImgReg5IN_141, F(12)=>
      ImgReg5IN_140, F(11)=>ImgReg5IN_139, F(10)=>ImgReg5IN_138, F(9)=>
      ImgReg5IN_137, F(8)=>ImgReg5IN_136, F(7)=>ImgReg5IN_135, F(6)=>
      ImgReg5IN_134, F(5)=>ImgReg5IN_133, F(4)=>ImgReg5IN_132, F(3)=>
      ImgReg5IN_131, F(2)=>ImgReg5IN_130, F(1)=>ImgReg5IN_129, F(0)=>
      ImgReg5IN_128);
   loop3_8_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_143_EXMPLR, D(14)=>OutputImg1_142_EXMPLR, D(13)=>
      OutputImg1_141_EXMPLR, D(12)=>OutputImg1_140_EXMPLR, D(11)=>
      OutputImg1_139_EXMPLR, D(10)=>OutputImg1_138_EXMPLR, D(9)=>
      OutputImg1_137_EXMPLR, D(8)=>OutputImg1_136_EXMPLR, D(7)=>
      OutputImg1_135_EXMPLR, D(6)=>OutputImg1_134_EXMPLR, D(5)=>
      OutputImg1_133_EXMPLR, D(4)=>OutputImg1_132_EXMPLR, D(3)=>
      OutputImg1_131_EXMPLR, D(2)=>OutputImg1_130_EXMPLR, D(1)=>
      OutputImg1_129_EXMPLR, D(0)=>OutputImg1_128_EXMPLR, EN=>nx23796, F(15)
      =>ImgReg0IN_143, F(14)=>ImgReg0IN_142, F(13)=>ImgReg0IN_141, F(12)=>
      ImgReg0IN_140, F(11)=>ImgReg0IN_139, F(10)=>ImgReg0IN_138, F(9)=>
      ImgReg0IN_137, F(8)=>ImgReg0IN_136, F(7)=>ImgReg0IN_135, F(6)=>
      ImgReg0IN_134, F(5)=>ImgReg0IN_133, F(4)=>ImgReg0IN_132, F(3)=>
      ImgReg0IN_131, F(2)=>ImgReg0IN_130, F(1)=>ImgReg0IN_129, F(0)=>
      ImgReg0IN_128);
   loop3_8_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_143_EXMPLR, D(14)=>OutputImg2_142_EXMPLR, D(13)=>
      OutputImg2_141_EXMPLR, D(12)=>OutputImg2_140_EXMPLR, D(11)=>
      OutputImg2_139_EXMPLR, D(10)=>OutputImg2_138_EXMPLR, D(9)=>
      OutputImg2_137_EXMPLR, D(8)=>OutputImg2_136_EXMPLR, D(7)=>
      OutputImg2_135_EXMPLR, D(6)=>OutputImg2_134_EXMPLR, D(5)=>
      OutputImg2_133_EXMPLR, D(4)=>OutputImg2_132_EXMPLR, D(3)=>
      OutputImg2_131_EXMPLR, D(2)=>OutputImg2_130_EXMPLR, D(1)=>
      OutputImg2_129_EXMPLR, D(0)=>OutputImg2_128_EXMPLR, EN=>nx23796, F(15)
      =>ImgReg1IN_143, F(14)=>ImgReg1IN_142, F(13)=>ImgReg1IN_141, F(12)=>
      ImgReg1IN_140, F(11)=>ImgReg1IN_139, F(10)=>ImgReg1IN_138, F(9)=>
      ImgReg1IN_137, F(8)=>ImgReg1IN_136, F(7)=>ImgReg1IN_135, F(6)=>
      ImgReg1IN_134, F(5)=>ImgReg1IN_133, F(4)=>ImgReg1IN_132, F(3)=>
      ImgReg1IN_131, F(2)=>ImgReg1IN_130, F(1)=>ImgReg1IN_129, F(0)=>
      ImgReg1IN_128);
   loop3_8_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_143_EXMPLR, D(14)=>OutputImg3_142_EXMPLR, D(13)=>
      OutputImg3_141_EXMPLR, D(12)=>OutputImg3_140_EXMPLR, D(11)=>
      OutputImg3_139_EXMPLR, D(10)=>OutputImg3_138_EXMPLR, D(9)=>
      OutputImg3_137_EXMPLR, D(8)=>OutputImg3_136_EXMPLR, D(7)=>
      OutputImg3_135_EXMPLR, D(6)=>OutputImg3_134_EXMPLR, D(5)=>
      OutputImg3_133_EXMPLR, D(4)=>OutputImg3_132_EXMPLR, D(3)=>
      OutputImg3_131_EXMPLR, D(2)=>OutputImg3_130_EXMPLR, D(1)=>
      OutputImg3_129_EXMPLR, D(0)=>OutputImg3_128_EXMPLR, EN=>nx23798, F(15)
      =>ImgReg2IN_143, F(14)=>ImgReg2IN_142, F(13)=>ImgReg2IN_141, F(12)=>
      ImgReg2IN_140, F(11)=>ImgReg2IN_139, F(10)=>ImgReg2IN_138, F(9)=>
      ImgReg2IN_137, F(8)=>ImgReg2IN_136, F(7)=>ImgReg2IN_135, F(6)=>
      ImgReg2IN_134, F(5)=>ImgReg2IN_133, F(4)=>ImgReg2IN_132, F(3)=>
      ImgReg2IN_131, F(2)=>ImgReg2IN_130, F(1)=>ImgReg2IN_129, F(0)=>
      ImgReg2IN_128);
   loop3_8_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_143_EXMPLR, D(14)=>OutputImg4_142_EXMPLR, D(13)=>
      OutputImg4_141_EXMPLR, D(12)=>OutputImg4_140_EXMPLR, D(11)=>
      OutputImg4_139_EXMPLR, D(10)=>OutputImg4_138_EXMPLR, D(9)=>
      OutputImg4_137_EXMPLR, D(8)=>OutputImg4_136_EXMPLR, D(7)=>
      OutputImg4_135_EXMPLR, D(6)=>OutputImg4_134_EXMPLR, D(5)=>
      OutputImg4_133_EXMPLR, D(4)=>OutputImg4_132_EXMPLR, D(3)=>
      OutputImg4_131_EXMPLR, D(2)=>OutputImg4_130_EXMPLR, D(1)=>
      OutputImg4_129_EXMPLR, D(0)=>OutputImg4_128_EXMPLR, EN=>nx23798, F(15)
      =>ImgReg3IN_143, F(14)=>ImgReg3IN_142, F(13)=>ImgReg3IN_141, F(12)=>
      ImgReg3IN_140, F(11)=>ImgReg3IN_139, F(10)=>ImgReg3IN_138, F(9)=>
      ImgReg3IN_137, F(8)=>ImgReg3IN_136, F(7)=>ImgReg3IN_135, F(6)=>
      ImgReg3IN_134, F(5)=>ImgReg3IN_133, F(4)=>ImgReg3IN_132, F(3)=>
      ImgReg3IN_131, F(2)=>ImgReg3IN_130, F(1)=>ImgReg3IN_129, F(0)=>
      ImgReg3IN_128);
   loop3_8_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_143_EXMPLR, D(14)=>OutputImg5_142_EXMPLR, D(13)=>
      OutputImg5_141_EXMPLR, D(12)=>OutputImg5_140_EXMPLR, D(11)=>
      OutputImg5_139_EXMPLR, D(10)=>OutputImg5_138_EXMPLR, D(9)=>
      OutputImg5_137_EXMPLR, D(8)=>OutputImg5_136_EXMPLR, D(7)=>
      OutputImg5_135_EXMPLR, D(6)=>OutputImg5_134_EXMPLR, D(5)=>
      OutputImg5_133_EXMPLR, D(4)=>OutputImg5_132_EXMPLR, D(3)=>
      OutputImg5_131_EXMPLR, D(2)=>OutputImg5_130_EXMPLR, D(1)=>
      OutputImg5_129_EXMPLR, D(0)=>OutputImg5_128_EXMPLR, EN=>nx23798, F(15)
      =>ImgReg4IN_143, F(14)=>ImgReg4IN_142, F(13)=>ImgReg4IN_141, F(12)=>
      ImgReg4IN_140, F(11)=>ImgReg4IN_139, F(10)=>ImgReg4IN_138, F(9)=>
      ImgReg4IN_137, F(8)=>ImgReg4IN_136, F(7)=>ImgReg4IN_135, F(6)=>
      ImgReg4IN_134, F(5)=>ImgReg4IN_133, F(4)=>ImgReg4IN_132, F(3)=>
      ImgReg4IN_131, F(2)=>ImgReg4IN_130, F(1)=>ImgReg4IN_129, F(0)=>
      ImgReg4IN_128);
   loop3_8_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_143, D(14)=>
      ImgReg0IN_142, D(13)=>ImgReg0IN_141, D(12)=>ImgReg0IN_140, D(11)=>
      ImgReg0IN_139, D(10)=>ImgReg0IN_138, D(9)=>ImgReg0IN_137, D(8)=>
      ImgReg0IN_136, D(7)=>ImgReg0IN_135, D(6)=>ImgReg0IN_134, D(5)=>
      ImgReg0IN_133, D(4)=>ImgReg0IN_132, D(3)=>ImgReg0IN_131, D(2)=>
      ImgReg0IN_130, D(1)=>ImgReg0IN_129, D(0)=>ImgReg0IN_128, CLK=>nx23876, 
      RST=>RST, EN=>nx23720, Q(15)=>OutputImg0_143_EXMPLR, Q(14)=>
      OutputImg0_142_EXMPLR, Q(13)=>OutputImg0_141_EXMPLR, Q(12)=>
      OutputImg0_140_EXMPLR, Q(11)=>OutputImg0_139_EXMPLR, Q(10)=>
      OutputImg0_138_EXMPLR, Q(9)=>OutputImg0_137_EXMPLR, Q(8)=>
      OutputImg0_136_EXMPLR, Q(7)=>OutputImg0_135_EXMPLR, Q(6)=>
      OutputImg0_134_EXMPLR, Q(5)=>OutputImg0_133_EXMPLR, Q(4)=>
      OutputImg0_132_EXMPLR, Q(3)=>OutputImg0_131_EXMPLR, Q(2)=>
      OutputImg0_130_EXMPLR, Q(1)=>OutputImg0_129_EXMPLR, Q(0)=>
      OutputImg0_128_EXMPLR);
   loop3_8_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_143, D(14)=>
      ImgReg1IN_142, D(13)=>ImgReg1IN_141, D(12)=>ImgReg1IN_140, D(11)=>
      ImgReg1IN_139, D(10)=>ImgReg1IN_138, D(9)=>ImgReg1IN_137, D(8)=>
      ImgReg1IN_136, D(7)=>ImgReg1IN_135, D(6)=>ImgReg1IN_134, D(5)=>
      ImgReg1IN_133, D(4)=>ImgReg1IN_132, D(3)=>ImgReg1IN_131, D(2)=>
      ImgReg1IN_130, D(1)=>ImgReg1IN_129, D(0)=>ImgReg1IN_128, CLK=>nx23878, 
      RST=>RST, EN=>nx23730, Q(15)=>OutputImg1_143_EXMPLR, Q(14)=>
      OutputImg1_142_EXMPLR, Q(13)=>OutputImg1_141_EXMPLR, Q(12)=>
      OutputImg1_140_EXMPLR, Q(11)=>OutputImg1_139_EXMPLR, Q(10)=>
      OutputImg1_138_EXMPLR, Q(9)=>OutputImg1_137_EXMPLR, Q(8)=>
      OutputImg1_136_EXMPLR, Q(7)=>OutputImg1_135_EXMPLR, Q(6)=>
      OutputImg1_134_EXMPLR, Q(5)=>OutputImg1_133_EXMPLR, Q(4)=>
      OutputImg1_132_EXMPLR, Q(3)=>OutputImg1_131_EXMPLR, Q(2)=>
      OutputImg1_130_EXMPLR, Q(1)=>OutputImg1_129_EXMPLR, Q(0)=>
      OutputImg1_128_EXMPLR);
   loop3_8_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_143, D(14)=>
      ImgReg2IN_142, D(13)=>ImgReg2IN_141, D(12)=>ImgReg2IN_140, D(11)=>
      ImgReg2IN_139, D(10)=>ImgReg2IN_138, D(9)=>ImgReg2IN_137, D(8)=>
      ImgReg2IN_136, D(7)=>ImgReg2IN_135, D(6)=>ImgReg2IN_134, D(5)=>
      ImgReg2IN_133, D(4)=>ImgReg2IN_132, D(3)=>ImgReg2IN_131, D(2)=>
      ImgReg2IN_130, D(1)=>ImgReg2IN_129, D(0)=>ImgReg2IN_128, CLK=>nx23878, 
      RST=>RST, EN=>nx23740, Q(15)=>OutputImg2_143_EXMPLR, Q(14)=>
      OutputImg2_142_EXMPLR, Q(13)=>OutputImg2_141_EXMPLR, Q(12)=>
      OutputImg2_140_EXMPLR, Q(11)=>OutputImg2_139_EXMPLR, Q(10)=>
      OutputImg2_138_EXMPLR, Q(9)=>OutputImg2_137_EXMPLR, Q(8)=>
      OutputImg2_136_EXMPLR, Q(7)=>OutputImg2_135_EXMPLR, Q(6)=>
      OutputImg2_134_EXMPLR, Q(5)=>OutputImg2_133_EXMPLR, Q(4)=>
      OutputImg2_132_EXMPLR, Q(3)=>OutputImg2_131_EXMPLR, Q(2)=>
      OutputImg2_130_EXMPLR, Q(1)=>OutputImg2_129_EXMPLR, Q(0)=>
      OutputImg2_128_EXMPLR);
   loop3_8_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_143, D(14)=>
      ImgReg3IN_142, D(13)=>ImgReg3IN_141, D(12)=>ImgReg3IN_140, D(11)=>
      ImgReg3IN_139, D(10)=>ImgReg3IN_138, D(9)=>ImgReg3IN_137, D(8)=>
      ImgReg3IN_136, D(7)=>ImgReg3IN_135, D(6)=>ImgReg3IN_134, D(5)=>
      ImgReg3IN_133, D(4)=>ImgReg3IN_132, D(3)=>ImgReg3IN_131, D(2)=>
      ImgReg3IN_130, D(1)=>ImgReg3IN_129, D(0)=>ImgReg3IN_128, CLK=>nx23880, 
      RST=>RST, EN=>nx23750, Q(15)=>OutputImg3_143_EXMPLR, Q(14)=>
      OutputImg3_142_EXMPLR, Q(13)=>OutputImg3_141_EXMPLR, Q(12)=>
      OutputImg3_140_EXMPLR, Q(11)=>OutputImg3_139_EXMPLR, Q(10)=>
      OutputImg3_138_EXMPLR, Q(9)=>OutputImg3_137_EXMPLR, Q(8)=>
      OutputImg3_136_EXMPLR, Q(7)=>OutputImg3_135_EXMPLR, Q(6)=>
      OutputImg3_134_EXMPLR, Q(5)=>OutputImg3_133_EXMPLR, Q(4)=>
      OutputImg3_132_EXMPLR, Q(3)=>OutputImg3_131_EXMPLR, Q(2)=>
      OutputImg3_130_EXMPLR, Q(1)=>OutputImg3_129_EXMPLR, Q(0)=>
      OutputImg3_128_EXMPLR);
   loop3_8_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_143, D(14)=>
      ImgReg4IN_142, D(13)=>ImgReg4IN_141, D(12)=>ImgReg4IN_140, D(11)=>
      ImgReg4IN_139, D(10)=>ImgReg4IN_138, D(9)=>ImgReg4IN_137, D(8)=>
      ImgReg4IN_136, D(7)=>ImgReg4IN_135, D(6)=>ImgReg4IN_134, D(5)=>
      ImgReg4IN_133, D(4)=>ImgReg4IN_132, D(3)=>ImgReg4IN_131, D(2)=>
      ImgReg4IN_130, D(1)=>ImgReg4IN_129, D(0)=>ImgReg4IN_128, CLK=>nx23880, 
      RST=>RST, EN=>nx23760, Q(15)=>OutputImg4_143_EXMPLR, Q(14)=>
      OutputImg4_142_EXMPLR, Q(13)=>OutputImg4_141_EXMPLR, Q(12)=>
      OutputImg4_140_EXMPLR, Q(11)=>OutputImg4_139_EXMPLR, Q(10)=>
      OutputImg4_138_EXMPLR, Q(9)=>OutputImg4_137_EXMPLR, Q(8)=>
      OutputImg4_136_EXMPLR, Q(7)=>OutputImg4_135_EXMPLR, Q(6)=>
      OutputImg4_134_EXMPLR, Q(5)=>OutputImg4_133_EXMPLR, Q(4)=>
      OutputImg4_132_EXMPLR, Q(3)=>OutputImg4_131_EXMPLR, Q(2)=>
      OutputImg4_130_EXMPLR, Q(1)=>OutputImg4_129_EXMPLR, Q(0)=>
      OutputImg4_128_EXMPLR);
   loop3_8_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_143, D(14)=>
      ImgReg5IN_142, D(13)=>ImgReg5IN_141, D(12)=>ImgReg5IN_140, D(11)=>
      ImgReg5IN_139, D(10)=>ImgReg5IN_138, D(9)=>ImgReg5IN_137, D(8)=>
      ImgReg5IN_136, D(7)=>ImgReg5IN_135, D(6)=>ImgReg5IN_134, D(5)=>
      ImgReg5IN_133, D(4)=>ImgReg5IN_132, D(3)=>ImgReg5IN_131, D(2)=>
      ImgReg5IN_130, D(1)=>ImgReg5IN_129, D(0)=>ImgReg5IN_128, CLK=>nx23882, 
      RST=>RST, EN=>nx23770, Q(15)=>OutputImg5_143_EXMPLR, Q(14)=>
      OutputImg5_142_EXMPLR, Q(13)=>OutputImg5_141_EXMPLR, Q(12)=>
      OutputImg5_140_EXMPLR, Q(11)=>OutputImg5_139_EXMPLR, Q(10)=>
      OutputImg5_138_EXMPLR, Q(9)=>OutputImg5_137_EXMPLR, Q(8)=>
      OutputImg5_136_EXMPLR, Q(7)=>OutputImg5_135_EXMPLR, Q(6)=>
      OutputImg5_134_EXMPLR, Q(5)=>OutputImg5_133_EXMPLR, Q(4)=>
      OutputImg5_132_EXMPLR, Q(3)=>OutputImg5_131_EXMPLR, Q(2)=>
      OutputImg5_130_EXMPLR, Q(1)=>OutputImg5_129_EXMPLR, Q(0)=>
      OutputImg5_128_EXMPLR);
   loop3_9_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_175_EXMPLR, D(14)=>OutputImg0_174_EXMPLR, D(13)=>
      OutputImg0_173_EXMPLR, D(12)=>OutputImg0_172_EXMPLR, D(11)=>
      OutputImg0_171_EXMPLR, D(10)=>OutputImg0_170_EXMPLR, D(9)=>
      OutputImg0_169_EXMPLR, D(8)=>OutputImg0_168_EXMPLR, D(7)=>
      OutputImg0_167_EXMPLR, D(6)=>OutputImg0_166_EXMPLR, D(5)=>
      OutputImg0_165_EXMPLR, D(4)=>OutputImg0_164_EXMPLR, D(3)=>
      OutputImg0_163_EXMPLR, D(2)=>OutputImg0_162_EXMPLR, D(1)=>
      OutputImg0_161_EXMPLR, D(0)=>OutputImg0_160_EXMPLR, EN=>nx23680, F(15)
      =>ImgReg0IN_159, F(14)=>ImgReg0IN_158, F(13)=>ImgReg0IN_157, F(12)=>
      ImgReg0IN_156, F(11)=>ImgReg0IN_155, F(10)=>ImgReg0IN_154, F(9)=>
      ImgReg0IN_153, F(8)=>ImgReg0IN_152, F(7)=>ImgReg0IN_151, F(6)=>
      ImgReg0IN_150, F(5)=>ImgReg0IN_149, F(4)=>ImgReg0IN_148, F(3)=>
      ImgReg0IN_147, F(2)=>ImgReg0IN_146, F(1)=>ImgReg0IN_145, F(0)=>
      ImgReg0IN_144);
   loop3_9_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_175_EXMPLR, D(14)=>OutputImg1_174_EXMPLR, D(13)=>
      OutputImg1_173_EXMPLR, D(12)=>OutputImg1_172_EXMPLR, D(11)=>
      OutputImg1_171_EXMPLR, D(10)=>OutputImg1_170_EXMPLR, D(9)=>
      OutputImg1_169_EXMPLR, D(8)=>OutputImg1_168_EXMPLR, D(7)=>
      OutputImg1_167_EXMPLR, D(6)=>OutputImg1_166_EXMPLR, D(5)=>
      OutputImg1_165_EXMPLR, D(4)=>OutputImg1_164_EXMPLR, D(3)=>
      OutputImg1_163_EXMPLR, D(2)=>OutputImg1_162_EXMPLR, D(1)=>
      OutputImg1_161_EXMPLR, D(0)=>OutputImg1_160_EXMPLR, EN=>nx23680, F(15)
      =>ImgReg1IN_159, F(14)=>ImgReg1IN_158, F(13)=>ImgReg1IN_157, F(12)=>
      ImgReg1IN_156, F(11)=>ImgReg1IN_155, F(10)=>ImgReg1IN_154, F(9)=>
      ImgReg1IN_153, F(8)=>ImgReg1IN_152, F(7)=>ImgReg1IN_151, F(6)=>
      ImgReg1IN_150, F(5)=>ImgReg1IN_149, F(4)=>ImgReg1IN_148, F(3)=>
      ImgReg1IN_147, F(2)=>ImgReg1IN_146, F(1)=>ImgReg1IN_145, F(0)=>
      ImgReg1IN_144);
   loop3_9_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_175_EXMPLR, D(14)=>OutputImg2_174_EXMPLR, D(13)=>
      OutputImg2_173_EXMPLR, D(12)=>OutputImg2_172_EXMPLR, D(11)=>
      OutputImg2_171_EXMPLR, D(10)=>OutputImg2_170_EXMPLR, D(9)=>
      OutputImg2_169_EXMPLR, D(8)=>OutputImg2_168_EXMPLR, D(7)=>
      OutputImg2_167_EXMPLR, D(6)=>OutputImg2_166_EXMPLR, D(5)=>
      OutputImg2_165_EXMPLR, D(4)=>OutputImg2_164_EXMPLR, D(3)=>
      OutputImg2_163_EXMPLR, D(2)=>OutputImg2_162_EXMPLR, D(1)=>
      OutputImg2_161_EXMPLR, D(0)=>OutputImg2_160_EXMPLR, EN=>nx23682, F(15)
      =>ImgReg2IN_159, F(14)=>ImgReg2IN_158, F(13)=>ImgReg2IN_157, F(12)=>
      ImgReg2IN_156, F(11)=>ImgReg2IN_155, F(10)=>ImgReg2IN_154, F(9)=>
      ImgReg2IN_153, F(8)=>ImgReg2IN_152, F(7)=>ImgReg2IN_151, F(6)=>
      ImgReg2IN_150, F(5)=>ImgReg2IN_149, F(4)=>ImgReg2IN_148, F(3)=>
      ImgReg2IN_147, F(2)=>ImgReg2IN_146, F(1)=>ImgReg2IN_145, F(0)=>
      ImgReg2IN_144);
   loop3_9_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_175_EXMPLR, D(14)=>OutputImg3_174_EXMPLR, D(13)=>
      OutputImg3_173_EXMPLR, D(12)=>OutputImg3_172_EXMPLR, D(11)=>
      OutputImg3_171_EXMPLR, D(10)=>OutputImg3_170_EXMPLR, D(9)=>
      OutputImg3_169_EXMPLR, D(8)=>OutputImg3_168_EXMPLR, D(7)=>
      OutputImg3_167_EXMPLR, D(6)=>OutputImg3_166_EXMPLR, D(5)=>
      OutputImg3_165_EXMPLR, D(4)=>OutputImg3_164_EXMPLR, D(3)=>
      OutputImg3_163_EXMPLR, D(2)=>OutputImg3_162_EXMPLR, D(1)=>
      OutputImg3_161_EXMPLR, D(0)=>OutputImg3_160_EXMPLR, EN=>nx23682, F(15)
      =>ImgReg3IN_159, F(14)=>ImgReg3IN_158, F(13)=>ImgReg3IN_157, F(12)=>
      ImgReg3IN_156, F(11)=>ImgReg3IN_155, F(10)=>ImgReg3IN_154, F(9)=>
      ImgReg3IN_153, F(8)=>ImgReg3IN_152, F(7)=>ImgReg3IN_151, F(6)=>
      ImgReg3IN_150, F(5)=>ImgReg3IN_149, F(4)=>ImgReg3IN_148, F(3)=>
      ImgReg3IN_147, F(2)=>ImgReg3IN_146, F(1)=>ImgReg3IN_145, F(0)=>
      ImgReg3IN_144);
   loop3_9_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_175_EXMPLR, D(14)=>OutputImg4_174_EXMPLR, D(13)=>
      OutputImg4_173_EXMPLR, D(12)=>OutputImg4_172_EXMPLR, D(11)=>
      OutputImg4_171_EXMPLR, D(10)=>OutputImg4_170_EXMPLR, D(9)=>
      OutputImg4_169_EXMPLR, D(8)=>OutputImg4_168_EXMPLR, D(7)=>
      OutputImg4_167_EXMPLR, D(6)=>OutputImg4_166_EXMPLR, D(5)=>
      OutputImg4_165_EXMPLR, D(4)=>OutputImg4_164_EXMPLR, D(3)=>
      OutputImg4_163_EXMPLR, D(2)=>OutputImg4_162_EXMPLR, D(1)=>
      OutputImg4_161_EXMPLR, D(0)=>OutputImg4_160_EXMPLR, EN=>nx23682, F(15)
      =>ImgReg4IN_159, F(14)=>ImgReg4IN_158, F(13)=>ImgReg4IN_157, F(12)=>
      ImgReg4IN_156, F(11)=>ImgReg4IN_155, F(10)=>ImgReg4IN_154, F(9)=>
      ImgReg4IN_153, F(8)=>ImgReg4IN_152, F(7)=>ImgReg4IN_151, F(6)=>
      ImgReg4IN_150, F(5)=>ImgReg4IN_149, F(4)=>ImgReg4IN_148, F(3)=>
      ImgReg4IN_147, F(2)=>ImgReg4IN_146, F(1)=>ImgReg4IN_145, F(0)=>
      ImgReg4IN_144);
   loop3_9_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_175_EXMPLR, D(14)=>OutputImg5_174_EXMPLR, D(13)=>
      OutputImg5_173_EXMPLR, D(12)=>OutputImg5_172_EXMPLR, D(11)=>
      OutputImg5_171_EXMPLR, D(10)=>OutputImg5_170_EXMPLR, D(9)=>
      OutputImg5_169_EXMPLR, D(8)=>OutputImg5_168_EXMPLR, D(7)=>
      OutputImg5_167_EXMPLR, D(6)=>OutputImg5_166_EXMPLR, D(5)=>
      OutputImg5_165_EXMPLR, D(4)=>OutputImg5_164_EXMPLR, D(3)=>
      OutputImg5_163_EXMPLR, D(2)=>OutputImg5_162_EXMPLR, D(1)=>
      OutputImg5_161_EXMPLR, D(0)=>OutputImg5_160_EXMPLR, EN=>nx23682, F(15)
      =>ImgReg5IN_159, F(14)=>ImgReg5IN_158, F(13)=>ImgReg5IN_157, F(12)=>
      ImgReg5IN_156, F(11)=>ImgReg5IN_155, F(10)=>ImgReg5IN_154, F(9)=>
      ImgReg5IN_153, F(8)=>ImgReg5IN_152, F(7)=>ImgReg5IN_151, F(6)=>
      ImgReg5IN_150, F(5)=>ImgReg5IN_149, F(4)=>ImgReg5IN_148, F(3)=>
      ImgReg5IN_147, F(2)=>ImgReg5IN_146, F(1)=>ImgReg5IN_145, F(0)=>
      ImgReg5IN_144);
   loop3_9_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(159), D(14)
      =>DATA(158), D(13)=>DATA(157), D(12)=>DATA(156), D(11)=>DATA(155), 
      D(10)=>DATA(154), D(9)=>DATA(153), D(8)=>DATA(152), D(7)=>DATA(151), 
      D(6)=>DATA(150), D(5)=>DATA(149), D(4)=>DATA(148), D(3)=>DATA(147), 
      D(2)=>DATA(146), D(1)=>DATA(145), D(0)=>DATA(144), EN=>nx23656, F(15)
      =>ImgReg0IN_159, F(14)=>ImgReg0IN_158, F(13)=>ImgReg0IN_157, F(12)=>
      ImgReg0IN_156, F(11)=>ImgReg0IN_155, F(10)=>ImgReg0IN_154, F(9)=>
      ImgReg0IN_153, F(8)=>ImgReg0IN_152, F(7)=>ImgReg0IN_151, F(6)=>
      ImgReg0IN_150, F(5)=>ImgReg0IN_149, F(4)=>ImgReg0IN_148, F(3)=>
      ImgReg0IN_147, F(2)=>ImgReg0IN_146, F(1)=>ImgReg0IN_145, F(0)=>
      ImgReg0IN_144);
   loop3_9_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(159), D(14)
      =>DATA(158), D(13)=>DATA(157), D(12)=>DATA(156), D(11)=>DATA(155), 
      D(10)=>DATA(154), D(9)=>DATA(153), D(8)=>DATA(152), D(7)=>DATA(151), 
      D(6)=>DATA(150), D(5)=>DATA(149), D(4)=>DATA(148), D(3)=>DATA(147), 
      D(2)=>DATA(146), D(1)=>DATA(145), D(0)=>DATA(144), EN=>nx23644, F(15)
      =>ImgReg1IN_159, F(14)=>ImgReg1IN_158, F(13)=>ImgReg1IN_157, F(12)=>
      ImgReg1IN_156, F(11)=>ImgReg1IN_155, F(10)=>ImgReg1IN_154, F(9)=>
      ImgReg1IN_153, F(8)=>ImgReg1IN_152, F(7)=>ImgReg1IN_151, F(6)=>
      ImgReg1IN_150, F(5)=>ImgReg1IN_149, F(4)=>ImgReg1IN_148, F(3)=>
      ImgReg1IN_147, F(2)=>ImgReg1IN_146, F(1)=>ImgReg1IN_145, F(0)=>
      ImgReg1IN_144);
   loop3_9_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(159), D(14)
      =>DATA(158), D(13)=>DATA(157), D(12)=>DATA(156), D(11)=>DATA(155), 
      D(10)=>DATA(154), D(9)=>DATA(153), D(8)=>DATA(152), D(7)=>DATA(151), 
      D(6)=>DATA(150), D(5)=>DATA(149), D(4)=>DATA(148), D(3)=>DATA(147), 
      D(2)=>DATA(146), D(1)=>DATA(145), D(0)=>DATA(144), EN=>nx23632, F(15)
      =>ImgReg2IN_159, F(14)=>ImgReg2IN_158, F(13)=>ImgReg2IN_157, F(12)=>
      ImgReg2IN_156, F(11)=>ImgReg2IN_155, F(10)=>ImgReg2IN_154, F(9)=>
      ImgReg2IN_153, F(8)=>ImgReg2IN_152, F(7)=>ImgReg2IN_151, F(6)=>
      ImgReg2IN_150, F(5)=>ImgReg2IN_149, F(4)=>ImgReg2IN_148, F(3)=>
      ImgReg2IN_147, F(2)=>ImgReg2IN_146, F(1)=>ImgReg2IN_145, F(0)=>
      ImgReg2IN_144);
   loop3_9_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(159), D(14)
      =>DATA(158), D(13)=>DATA(157), D(12)=>DATA(156), D(11)=>DATA(155), 
      D(10)=>DATA(154), D(9)=>DATA(153), D(8)=>DATA(152), D(7)=>DATA(151), 
      D(6)=>DATA(150), D(5)=>DATA(149), D(4)=>DATA(148), D(3)=>DATA(147), 
      D(2)=>DATA(146), D(1)=>DATA(145), D(0)=>DATA(144), EN=>nx23620, F(15)
      =>ImgReg3IN_159, F(14)=>ImgReg3IN_158, F(13)=>ImgReg3IN_157, F(12)=>
      ImgReg3IN_156, F(11)=>ImgReg3IN_155, F(10)=>ImgReg3IN_154, F(9)=>
      ImgReg3IN_153, F(8)=>ImgReg3IN_152, F(7)=>ImgReg3IN_151, F(6)=>
      ImgReg3IN_150, F(5)=>ImgReg3IN_149, F(4)=>ImgReg3IN_148, F(3)=>
      ImgReg3IN_147, F(2)=>ImgReg3IN_146, F(1)=>ImgReg3IN_145, F(0)=>
      ImgReg3IN_144);
   loop3_9_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(159), D(14)
      =>DATA(158), D(13)=>DATA(157), D(12)=>DATA(156), D(11)=>DATA(155), 
      D(10)=>DATA(154), D(9)=>DATA(153), D(8)=>DATA(152), D(7)=>DATA(151), 
      D(6)=>DATA(150), D(5)=>DATA(149), D(4)=>DATA(148), D(3)=>DATA(147), 
      D(2)=>DATA(146), D(1)=>DATA(145), D(0)=>DATA(144), EN=>nx23608, F(15)
      =>ImgReg4IN_159, F(14)=>ImgReg4IN_158, F(13)=>ImgReg4IN_157, F(12)=>
      ImgReg4IN_156, F(11)=>ImgReg4IN_155, F(10)=>ImgReg4IN_154, F(9)=>
      ImgReg4IN_153, F(8)=>ImgReg4IN_152, F(7)=>ImgReg4IN_151, F(6)=>
      ImgReg4IN_150, F(5)=>ImgReg4IN_149, F(4)=>ImgReg4IN_148, F(3)=>
      ImgReg4IN_147, F(2)=>ImgReg4IN_146, F(1)=>ImgReg4IN_145, F(0)=>
      ImgReg4IN_144);
   loop3_9_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(159), D(14)
      =>DATA(158), D(13)=>DATA(157), D(12)=>DATA(156), D(11)=>DATA(155), 
      D(10)=>DATA(154), D(9)=>DATA(153), D(8)=>DATA(152), D(7)=>DATA(151), 
      D(6)=>DATA(150), D(5)=>DATA(149), D(4)=>DATA(148), D(3)=>DATA(147), 
      D(2)=>DATA(146), D(1)=>DATA(145), D(0)=>DATA(144), EN=>nx23596, F(15)
      =>ImgReg5IN_159, F(14)=>ImgReg5IN_158, F(13)=>ImgReg5IN_157, F(12)=>
      ImgReg5IN_156, F(11)=>ImgReg5IN_155, F(10)=>ImgReg5IN_154, F(9)=>
      ImgReg5IN_153, F(8)=>ImgReg5IN_152, F(7)=>ImgReg5IN_151, F(6)=>
      ImgReg5IN_150, F(5)=>ImgReg5IN_149, F(4)=>ImgReg5IN_148, F(3)=>
      ImgReg5IN_147, F(2)=>ImgReg5IN_146, F(1)=>ImgReg5IN_145, F(0)=>
      ImgReg5IN_144);
   loop3_9_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_159_EXMPLR, D(14)=>OutputImg1_158_EXMPLR, D(13)=>
      OutputImg1_157_EXMPLR, D(12)=>OutputImg1_156_EXMPLR, D(11)=>
      OutputImg1_155_EXMPLR, D(10)=>OutputImg1_154_EXMPLR, D(9)=>
      OutputImg1_153_EXMPLR, D(8)=>OutputImg1_152_EXMPLR, D(7)=>
      OutputImg1_151_EXMPLR, D(6)=>OutputImg1_150_EXMPLR, D(5)=>
      OutputImg1_149_EXMPLR, D(4)=>OutputImg1_148_EXMPLR, D(3)=>
      OutputImg1_147_EXMPLR, D(2)=>OutputImg1_146_EXMPLR, D(1)=>
      OutputImg1_145_EXMPLR, D(0)=>OutputImg1_144_EXMPLR, EN=>nx23798, F(15)
      =>ImgReg0IN_159, F(14)=>ImgReg0IN_158, F(13)=>ImgReg0IN_157, F(12)=>
      ImgReg0IN_156, F(11)=>ImgReg0IN_155, F(10)=>ImgReg0IN_154, F(9)=>
      ImgReg0IN_153, F(8)=>ImgReg0IN_152, F(7)=>ImgReg0IN_151, F(6)=>
      ImgReg0IN_150, F(5)=>ImgReg0IN_149, F(4)=>ImgReg0IN_148, F(3)=>
      ImgReg0IN_147, F(2)=>ImgReg0IN_146, F(1)=>ImgReg0IN_145, F(0)=>
      ImgReg0IN_144);
   loop3_9_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_159_EXMPLR, D(14)=>OutputImg2_158_EXMPLR, D(13)=>
      OutputImg2_157_EXMPLR, D(12)=>OutputImg2_156_EXMPLR, D(11)=>
      OutputImg2_155_EXMPLR, D(10)=>OutputImg2_154_EXMPLR, D(9)=>
      OutputImg2_153_EXMPLR, D(8)=>OutputImg2_152_EXMPLR, D(7)=>
      OutputImg2_151_EXMPLR, D(6)=>OutputImg2_150_EXMPLR, D(5)=>
      OutputImg2_149_EXMPLR, D(4)=>OutputImg2_148_EXMPLR, D(3)=>
      OutputImg2_147_EXMPLR, D(2)=>OutputImg2_146_EXMPLR, D(1)=>
      OutputImg2_145_EXMPLR, D(0)=>OutputImg2_144_EXMPLR, EN=>nx23798, F(15)
      =>ImgReg1IN_159, F(14)=>ImgReg1IN_158, F(13)=>ImgReg1IN_157, F(12)=>
      ImgReg1IN_156, F(11)=>ImgReg1IN_155, F(10)=>ImgReg1IN_154, F(9)=>
      ImgReg1IN_153, F(8)=>ImgReg1IN_152, F(7)=>ImgReg1IN_151, F(6)=>
      ImgReg1IN_150, F(5)=>ImgReg1IN_149, F(4)=>ImgReg1IN_148, F(3)=>
      ImgReg1IN_147, F(2)=>ImgReg1IN_146, F(1)=>ImgReg1IN_145, F(0)=>
      ImgReg1IN_144);
   loop3_9_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_159_EXMPLR, D(14)=>OutputImg3_158_EXMPLR, D(13)=>
      OutputImg3_157_EXMPLR, D(12)=>OutputImg3_156_EXMPLR, D(11)=>
      OutputImg3_155_EXMPLR, D(10)=>OutputImg3_154_EXMPLR, D(9)=>
      OutputImg3_153_EXMPLR, D(8)=>OutputImg3_152_EXMPLR, D(7)=>
      OutputImg3_151_EXMPLR, D(6)=>OutputImg3_150_EXMPLR, D(5)=>
      OutputImg3_149_EXMPLR, D(4)=>OutputImg3_148_EXMPLR, D(3)=>
      OutputImg3_147_EXMPLR, D(2)=>OutputImg3_146_EXMPLR, D(1)=>
      OutputImg3_145_EXMPLR, D(0)=>OutputImg3_144_EXMPLR, EN=>nx23798, F(15)
      =>ImgReg2IN_159, F(14)=>ImgReg2IN_158, F(13)=>ImgReg2IN_157, F(12)=>
      ImgReg2IN_156, F(11)=>ImgReg2IN_155, F(10)=>ImgReg2IN_154, F(9)=>
      ImgReg2IN_153, F(8)=>ImgReg2IN_152, F(7)=>ImgReg2IN_151, F(6)=>
      ImgReg2IN_150, F(5)=>ImgReg2IN_149, F(4)=>ImgReg2IN_148, F(3)=>
      ImgReg2IN_147, F(2)=>ImgReg2IN_146, F(1)=>ImgReg2IN_145, F(0)=>
      ImgReg2IN_144);
   loop3_9_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_159_EXMPLR, D(14)=>OutputImg4_158_EXMPLR, D(13)=>
      OutputImg4_157_EXMPLR, D(12)=>OutputImg4_156_EXMPLR, D(11)=>
      OutputImg4_155_EXMPLR, D(10)=>OutputImg4_154_EXMPLR, D(9)=>
      OutputImg4_153_EXMPLR, D(8)=>OutputImg4_152_EXMPLR, D(7)=>
      OutputImg4_151_EXMPLR, D(6)=>OutputImg4_150_EXMPLR, D(5)=>
      OutputImg4_149_EXMPLR, D(4)=>OutputImg4_148_EXMPLR, D(3)=>
      OutputImg4_147_EXMPLR, D(2)=>OutputImg4_146_EXMPLR, D(1)=>
      OutputImg4_145_EXMPLR, D(0)=>OutputImg4_144_EXMPLR, EN=>nx23798, F(15)
      =>ImgReg3IN_159, F(14)=>ImgReg3IN_158, F(13)=>ImgReg3IN_157, F(12)=>
      ImgReg3IN_156, F(11)=>ImgReg3IN_155, F(10)=>ImgReg3IN_154, F(9)=>
      ImgReg3IN_153, F(8)=>ImgReg3IN_152, F(7)=>ImgReg3IN_151, F(6)=>
      ImgReg3IN_150, F(5)=>ImgReg3IN_149, F(4)=>ImgReg3IN_148, F(3)=>
      ImgReg3IN_147, F(2)=>ImgReg3IN_146, F(1)=>ImgReg3IN_145, F(0)=>
      ImgReg3IN_144);
   loop3_9_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_159_EXMPLR, D(14)=>OutputImg5_158_EXMPLR, D(13)=>
      OutputImg5_157_EXMPLR, D(12)=>OutputImg5_156_EXMPLR, D(11)=>
      OutputImg5_155_EXMPLR, D(10)=>OutputImg5_154_EXMPLR, D(9)=>
      OutputImg5_153_EXMPLR, D(8)=>OutputImg5_152_EXMPLR, D(7)=>
      OutputImg5_151_EXMPLR, D(6)=>OutputImg5_150_EXMPLR, D(5)=>
      OutputImg5_149_EXMPLR, D(4)=>OutputImg5_148_EXMPLR, D(3)=>
      OutputImg5_147_EXMPLR, D(2)=>OutputImg5_146_EXMPLR, D(1)=>
      OutputImg5_145_EXMPLR, D(0)=>OutputImg5_144_EXMPLR, EN=>nx23800, F(15)
      =>ImgReg4IN_159, F(14)=>ImgReg4IN_158, F(13)=>ImgReg4IN_157, F(12)=>
      ImgReg4IN_156, F(11)=>ImgReg4IN_155, F(10)=>ImgReg4IN_154, F(9)=>
      ImgReg4IN_153, F(8)=>ImgReg4IN_152, F(7)=>ImgReg4IN_151, F(6)=>
      ImgReg4IN_150, F(5)=>ImgReg4IN_149, F(4)=>ImgReg4IN_148, F(3)=>
      ImgReg4IN_147, F(2)=>ImgReg4IN_146, F(1)=>ImgReg4IN_145, F(0)=>
      ImgReg4IN_144);
   loop3_9_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_159, D(14)=>
      ImgReg0IN_158, D(13)=>ImgReg0IN_157, D(12)=>ImgReg0IN_156, D(11)=>
      ImgReg0IN_155, D(10)=>ImgReg0IN_154, D(9)=>ImgReg0IN_153, D(8)=>
      ImgReg0IN_152, D(7)=>ImgReg0IN_151, D(6)=>ImgReg0IN_150, D(5)=>
      ImgReg0IN_149, D(4)=>ImgReg0IN_148, D(3)=>ImgReg0IN_147, D(2)=>
      ImgReg0IN_146, D(1)=>ImgReg0IN_145, D(0)=>ImgReg0IN_144, CLK=>nx23882, 
      RST=>RST, EN=>nx23720, Q(15)=>OutputImg0_159_EXMPLR, Q(14)=>
      OutputImg0_158_EXMPLR, Q(13)=>OutputImg0_157_EXMPLR, Q(12)=>
      OutputImg0_156_EXMPLR, Q(11)=>OutputImg0_155_EXMPLR, Q(10)=>
      OutputImg0_154_EXMPLR, Q(9)=>OutputImg0_153_EXMPLR, Q(8)=>
      OutputImg0_152_EXMPLR, Q(7)=>OutputImg0_151_EXMPLR, Q(6)=>
      OutputImg0_150_EXMPLR, Q(5)=>OutputImg0_149_EXMPLR, Q(4)=>
      OutputImg0_148_EXMPLR, Q(3)=>OutputImg0_147_EXMPLR, Q(2)=>
      OutputImg0_146_EXMPLR, Q(1)=>OutputImg0_145_EXMPLR, Q(0)=>
      OutputImg0_144_EXMPLR);
   loop3_9_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_159, D(14)=>
      ImgReg1IN_158, D(13)=>ImgReg1IN_157, D(12)=>ImgReg1IN_156, D(11)=>
      ImgReg1IN_155, D(10)=>ImgReg1IN_154, D(9)=>ImgReg1IN_153, D(8)=>
      ImgReg1IN_152, D(7)=>ImgReg1IN_151, D(6)=>ImgReg1IN_150, D(5)=>
      ImgReg1IN_149, D(4)=>ImgReg1IN_148, D(3)=>ImgReg1IN_147, D(2)=>
      ImgReg1IN_146, D(1)=>ImgReg1IN_145, D(0)=>ImgReg1IN_144, CLK=>nx23884, 
      RST=>RST, EN=>nx23730, Q(15)=>OutputImg1_159_EXMPLR, Q(14)=>
      OutputImg1_158_EXMPLR, Q(13)=>OutputImg1_157_EXMPLR, Q(12)=>
      OutputImg1_156_EXMPLR, Q(11)=>OutputImg1_155_EXMPLR, Q(10)=>
      OutputImg1_154_EXMPLR, Q(9)=>OutputImg1_153_EXMPLR, Q(8)=>
      OutputImg1_152_EXMPLR, Q(7)=>OutputImg1_151_EXMPLR, Q(6)=>
      OutputImg1_150_EXMPLR, Q(5)=>OutputImg1_149_EXMPLR, Q(4)=>
      OutputImg1_148_EXMPLR, Q(3)=>OutputImg1_147_EXMPLR, Q(2)=>
      OutputImg1_146_EXMPLR, Q(1)=>OutputImg1_145_EXMPLR, Q(0)=>
      OutputImg1_144_EXMPLR);
   loop3_9_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_159, D(14)=>
      ImgReg2IN_158, D(13)=>ImgReg2IN_157, D(12)=>ImgReg2IN_156, D(11)=>
      ImgReg2IN_155, D(10)=>ImgReg2IN_154, D(9)=>ImgReg2IN_153, D(8)=>
      ImgReg2IN_152, D(7)=>ImgReg2IN_151, D(6)=>ImgReg2IN_150, D(5)=>
      ImgReg2IN_149, D(4)=>ImgReg2IN_148, D(3)=>ImgReg2IN_147, D(2)=>
      ImgReg2IN_146, D(1)=>ImgReg2IN_145, D(0)=>ImgReg2IN_144, CLK=>nx23884, 
      RST=>RST, EN=>nx23740, Q(15)=>OutputImg2_159_EXMPLR, Q(14)=>
      OutputImg2_158_EXMPLR, Q(13)=>OutputImg2_157_EXMPLR, Q(12)=>
      OutputImg2_156_EXMPLR, Q(11)=>OutputImg2_155_EXMPLR, Q(10)=>
      OutputImg2_154_EXMPLR, Q(9)=>OutputImg2_153_EXMPLR, Q(8)=>
      OutputImg2_152_EXMPLR, Q(7)=>OutputImg2_151_EXMPLR, Q(6)=>
      OutputImg2_150_EXMPLR, Q(5)=>OutputImg2_149_EXMPLR, Q(4)=>
      OutputImg2_148_EXMPLR, Q(3)=>OutputImg2_147_EXMPLR, Q(2)=>
      OutputImg2_146_EXMPLR, Q(1)=>OutputImg2_145_EXMPLR, Q(0)=>
      OutputImg2_144_EXMPLR);
   loop3_9_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_159, D(14)=>
      ImgReg3IN_158, D(13)=>ImgReg3IN_157, D(12)=>ImgReg3IN_156, D(11)=>
      ImgReg3IN_155, D(10)=>ImgReg3IN_154, D(9)=>ImgReg3IN_153, D(8)=>
      ImgReg3IN_152, D(7)=>ImgReg3IN_151, D(6)=>ImgReg3IN_150, D(5)=>
      ImgReg3IN_149, D(4)=>ImgReg3IN_148, D(3)=>ImgReg3IN_147, D(2)=>
      ImgReg3IN_146, D(1)=>ImgReg3IN_145, D(0)=>ImgReg3IN_144, CLK=>nx23886, 
      RST=>RST, EN=>nx23750, Q(15)=>OutputImg3_159_EXMPLR, Q(14)=>
      OutputImg3_158_EXMPLR, Q(13)=>OutputImg3_157_EXMPLR, Q(12)=>
      OutputImg3_156_EXMPLR, Q(11)=>OutputImg3_155_EXMPLR, Q(10)=>
      OutputImg3_154_EXMPLR, Q(9)=>OutputImg3_153_EXMPLR, Q(8)=>
      OutputImg3_152_EXMPLR, Q(7)=>OutputImg3_151_EXMPLR, Q(6)=>
      OutputImg3_150_EXMPLR, Q(5)=>OutputImg3_149_EXMPLR, Q(4)=>
      OutputImg3_148_EXMPLR, Q(3)=>OutputImg3_147_EXMPLR, Q(2)=>
      OutputImg3_146_EXMPLR, Q(1)=>OutputImg3_145_EXMPLR, Q(0)=>
      OutputImg3_144_EXMPLR);
   loop3_9_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_159, D(14)=>
      ImgReg4IN_158, D(13)=>ImgReg4IN_157, D(12)=>ImgReg4IN_156, D(11)=>
      ImgReg4IN_155, D(10)=>ImgReg4IN_154, D(9)=>ImgReg4IN_153, D(8)=>
      ImgReg4IN_152, D(7)=>ImgReg4IN_151, D(6)=>ImgReg4IN_150, D(5)=>
      ImgReg4IN_149, D(4)=>ImgReg4IN_148, D(3)=>ImgReg4IN_147, D(2)=>
      ImgReg4IN_146, D(1)=>ImgReg4IN_145, D(0)=>ImgReg4IN_144, CLK=>nx23886, 
      RST=>RST, EN=>nx23760, Q(15)=>OutputImg4_159_EXMPLR, Q(14)=>
      OutputImg4_158_EXMPLR, Q(13)=>OutputImg4_157_EXMPLR, Q(12)=>
      OutputImg4_156_EXMPLR, Q(11)=>OutputImg4_155_EXMPLR, Q(10)=>
      OutputImg4_154_EXMPLR, Q(9)=>OutputImg4_153_EXMPLR, Q(8)=>
      OutputImg4_152_EXMPLR, Q(7)=>OutputImg4_151_EXMPLR, Q(6)=>
      OutputImg4_150_EXMPLR, Q(5)=>OutputImg4_149_EXMPLR, Q(4)=>
      OutputImg4_148_EXMPLR, Q(3)=>OutputImg4_147_EXMPLR, Q(2)=>
      OutputImg4_146_EXMPLR, Q(1)=>OutputImg4_145_EXMPLR, Q(0)=>
      OutputImg4_144_EXMPLR);
   loop3_9_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_159, D(14)=>
      ImgReg5IN_158, D(13)=>ImgReg5IN_157, D(12)=>ImgReg5IN_156, D(11)=>
      ImgReg5IN_155, D(10)=>ImgReg5IN_154, D(9)=>ImgReg5IN_153, D(8)=>
      ImgReg5IN_152, D(7)=>ImgReg5IN_151, D(6)=>ImgReg5IN_150, D(5)=>
      ImgReg5IN_149, D(4)=>ImgReg5IN_148, D(3)=>ImgReg5IN_147, D(2)=>
      ImgReg5IN_146, D(1)=>ImgReg5IN_145, D(0)=>ImgReg5IN_144, CLK=>nx23888, 
      RST=>RST, EN=>nx23770, Q(15)=>OutputImg5_159_EXMPLR, Q(14)=>
      OutputImg5_158_EXMPLR, Q(13)=>OutputImg5_157_EXMPLR, Q(12)=>
      OutputImg5_156_EXMPLR, Q(11)=>OutputImg5_155_EXMPLR, Q(10)=>
      OutputImg5_154_EXMPLR, Q(9)=>OutputImg5_153_EXMPLR, Q(8)=>
      OutputImg5_152_EXMPLR, Q(7)=>OutputImg5_151_EXMPLR, Q(6)=>
      OutputImg5_150_EXMPLR, Q(5)=>OutputImg5_149_EXMPLR, Q(4)=>
      OutputImg5_148_EXMPLR, Q(3)=>OutputImg5_147_EXMPLR, Q(2)=>
      OutputImg5_146_EXMPLR, Q(1)=>OutputImg5_145_EXMPLR, Q(0)=>
      OutputImg5_144_EXMPLR);
   loop3_10_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_191_EXMPLR, D(14)=>OutputImg0_190_EXMPLR, D(13)=>
      OutputImg0_189_EXMPLR, D(12)=>OutputImg0_188_EXMPLR, D(11)=>
      OutputImg0_187_EXMPLR, D(10)=>OutputImg0_186_EXMPLR, D(9)=>
      OutputImg0_185_EXMPLR, D(8)=>OutputImg0_184_EXMPLR, D(7)=>
      OutputImg0_183_EXMPLR, D(6)=>OutputImg0_182_EXMPLR, D(5)=>
      OutputImg0_181_EXMPLR, D(4)=>OutputImg0_180_EXMPLR, D(3)=>
      OutputImg0_179_EXMPLR, D(2)=>OutputImg0_178_EXMPLR, D(1)=>
      OutputImg0_177_EXMPLR, D(0)=>OutputImg0_176_EXMPLR, EN=>nx23682, F(15)
      =>ImgReg0IN_175, F(14)=>ImgReg0IN_174, F(13)=>ImgReg0IN_173, F(12)=>
      ImgReg0IN_172, F(11)=>ImgReg0IN_171, F(10)=>ImgReg0IN_170, F(9)=>
      ImgReg0IN_169, F(8)=>ImgReg0IN_168, F(7)=>ImgReg0IN_167, F(6)=>
      ImgReg0IN_166, F(5)=>ImgReg0IN_165, F(4)=>ImgReg0IN_164, F(3)=>
      ImgReg0IN_163, F(2)=>ImgReg0IN_162, F(1)=>ImgReg0IN_161, F(0)=>
      ImgReg0IN_160);
   loop3_10_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_191_EXMPLR, D(14)=>OutputImg1_190_EXMPLR, D(13)=>
      OutputImg1_189_EXMPLR, D(12)=>OutputImg1_188_EXMPLR, D(11)=>
      OutputImg1_187_EXMPLR, D(10)=>OutputImg1_186_EXMPLR, D(9)=>
      OutputImg1_185_EXMPLR, D(8)=>OutputImg1_184_EXMPLR, D(7)=>
      OutputImg1_183_EXMPLR, D(6)=>OutputImg1_182_EXMPLR, D(5)=>
      OutputImg1_181_EXMPLR, D(4)=>OutputImg1_180_EXMPLR, D(3)=>
      OutputImg1_179_EXMPLR, D(2)=>OutputImg1_178_EXMPLR, D(1)=>
      OutputImg1_177_EXMPLR, D(0)=>OutputImg1_176_EXMPLR, EN=>nx23682, F(15)
      =>ImgReg1IN_175, F(14)=>ImgReg1IN_174, F(13)=>ImgReg1IN_173, F(12)=>
      ImgReg1IN_172, F(11)=>ImgReg1IN_171, F(10)=>ImgReg1IN_170, F(9)=>
      ImgReg1IN_169, F(8)=>ImgReg1IN_168, F(7)=>ImgReg1IN_167, F(6)=>
      ImgReg1IN_166, F(5)=>ImgReg1IN_165, F(4)=>ImgReg1IN_164, F(3)=>
      ImgReg1IN_163, F(2)=>ImgReg1IN_162, F(1)=>ImgReg1IN_161, F(0)=>
      ImgReg1IN_160);
   loop3_10_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_191_EXMPLR, D(14)=>OutputImg2_190_EXMPLR, D(13)=>
      OutputImg2_189_EXMPLR, D(12)=>OutputImg2_188_EXMPLR, D(11)=>
      OutputImg2_187_EXMPLR, D(10)=>OutputImg2_186_EXMPLR, D(9)=>
      OutputImg2_185_EXMPLR, D(8)=>OutputImg2_184_EXMPLR, D(7)=>
      OutputImg2_183_EXMPLR, D(6)=>OutputImg2_182_EXMPLR, D(5)=>
      OutputImg2_181_EXMPLR, D(4)=>OutputImg2_180_EXMPLR, D(3)=>
      OutputImg2_179_EXMPLR, D(2)=>OutputImg2_178_EXMPLR, D(1)=>
      OutputImg2_177_EXMPLR, D(0)=>OutputImg2_176_EXMPLR, EN=>nx23682, F(15)
      =>ImgReg2IN_175, F(14)=>ImgReg2IN_174, F(13)=>ImgReg2IN_173, F(12)=>
      ImgReg2IN_172, F(11)=>ImgReg2IN_171, F(10)=>ImgReg2IN_170, F(9)=>
      ImgReg2IN_169, F(8)=>ImgReg2IN_168, F(7)=>ImgReg2IN_167, F(6)=>
      ImgReg2IN_166, F(5)=>ImgReg2IN_165, F(4)=>ImgReg2IN_164, F(3)=>
      ImgReg2IN_163, F(2)=>ImgReg2IN_162, F(1)=>ImgReg2IN_161, F(0)=>
      ImgReg2IN_160);
   loop3_10_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_191_EXMPLR, D(14)=>OutputImg3_190_EXMPLR, D(13)=>
      OutputImg3_189_EXMPLR, D(12)=>OutputImg3_188_EXMPLR, D(11)=>
      OutputImg3_187_EXMPLR, D(10)=>OutputImg3_186_EXMPLR, D(9)=>
      OutputImg3_185_EXMPLR, D(8)=>OutputImg3_184_EXMPLR, D(7)=>
      OutputImg3_183_EXMPLR, D(6)=>OutputImg3_182_EXMPLR, D(5)=>
      OutputImg3_181_EXMPLR, D(4)=>OutputImg3_180_EXMPLR, D(3)=>
      OutputImg3_179_EXMPLR, D(2)=>OutputImg3_178_EXMPLR, D(1)=>
      OutputImg3_177_EXMPLR, D(0)=>OutputImg3_176_EXMPLR, EN=>nx23684, F(15)
      =>ImgReg3IN_175, F(14)=>ImgReg3IN_174, F(13)=>ImgReg3IN_173, F(12)=>
      ImgReg3IN_172, F(11)=>ImgReg3IN_171, F(10)=>ImgReg3IN_170, F(9)=>
      ImgReg3IN_169, F(8)=>ImgReg3IN_168, F(7)=>ImgReg3IN_167, F(6)=>
      ImgReg3IN_166, F(5)=>ImgReg3IN_165, F(4)=>ImgReg3IN_164, F(3)=>
      ImgReg3IN_163, F(2)=>ImgReg3IN_162, F(1)=>ImgReg3IN_161, F(0)=>
      ImgReg3IN_160);
   loop3_10_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_191_EXMPLR, D(14)=>OutputImg4_190_EXMPLR, D(13)=>
      OutputImg4_189_EXMPLR, D(12)=>OutputImg4_188_EXMPLR, D(11)=>
      OutputImg4_187_EXMPLR, D(10)=>OutputImg4_186_EXMPLR, D(9)=>
      OutputImg4_185_EXMPLR, D(8)=>OutputImg4_184_EXMPLR, D(7)=>
      OutputImg4_183_EXMPLR, D(6)=>OutputImg4_182_EXMPLR, D(5)=>
      OutputImg4_181_EXMPLR, D(4)=>OutputImg4_180_EXMPLR, D(3)=>
      OutputImg4_179_EXMPLR, D(2)=>OutputImg4_178_EXMPLR, D(1)=>
      OutputImg4_177_EXMPLR, D(0)=>OutputImg4_176_EXMPLR, EN=>nx23684, F(15)
      =>ImgReg4IN_175, F(14)=>ImgReg4IN_174, F(13)=>ImgReg4IN_173, F(12)=>
      ImgReg4IN_172, F(11)=>ImgReg4IN_171, F(10)=>ImgReg4IN_170, F(9)=>
      ImgReg4IN_169, F(8)=>ImgReg4IN_168, F(7)=>ImgReg4IN_167, F(6)=>
      ImgReg4IN_166, F(5)=>ImgReg4IN_165, F(4)=>ImgReg4IN_164, F(3)=>
      ImgReg4IN_163, F(2)=>ImgReg4IN_162, F(1)=>ImgReg4IN_161, F(0)=>
      ImgReg4IN_160);
   loop3_10_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_191_EXMPLR, D(14)=>OutputImg5_190_EXMPLR, D(13)=>
      OutputImg5_189_EXMPLR, D(12)=>OutputImg5_188_EXMPLR, D(11)=>
      OutputImg5_187_EXMPLR, D(10)=>OutputImg5_186_EXMPLR, D(9)=>
      OutputImg5_185_EXMPLR, D(8)=>OutputImg5_184_EXMPLR, D(7)=>
      OutputImg5_183_EXMPLR, D(6)=>OutputImg5_182_EXMPLR, D(5)=>
      OutputImg5_181_EXMPLR, D(4)=>OutputImg5_180_EXMPLR, D(3)=>
      OutputImg5_179_EXMPLR, D(2)=>OutputImg5_178_EXMPLR, D(1)=>
      OutputImg5_177_EXMPLR, D(0)=>OutputImg5_176_EXMPLR, EN=>nx23684, F(15)
      =>ImgReg5IN_175, F(14)=>ImgReg5IN_174, F(13)=>ImgReg5IN_173, F(12)=>
      ImgReg5IN_172, F(11)=>ImgReg5IN_171, F(10)=>ImgReg5IN_170, F(9)=>
      ImgReg5IN_169, F(8)=>ImgReg5IN_168, F(7)=>ImgReg5IN_167, F(6)=>
      ImgReg5IN_166, F(5)=>ImgReg5IN_165, F(4)=>ImgReg5IN_164, F(3)=>
      ImgReg5IN_163, F(2)=>ImgReg5IN_162, F(1)=>ImgReg5IN_161, F(0)=>
      ImgReg5IN_160);
   loop3_10_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(175), 
      D(14)=>DATA(174), D(13)=>DATA(173), D(12)=>DATA(172), D(11)=>DATA(171), 
      D(10)=>DATA(170), D(9)=>DATA(169), D(8)=>DATA(168), D(7)=>DATA(167), 
      D(6)=>DATA(166), D(5)=>DATA(165), D(4)=>DATA(164), D(3)=>DATA(163), 
      D(2)=>DATA(162), D(1)=>DATA(161), D(0)=>DATA(160), EN=>nx23656, F(15)
      =>ImgReg0IN_175, F(14)=>ImgReg0IN_174, F(13)=>ImgReg0IN_173, F(12)=>
      ImgReg0IN_172, F(11)=>ImgReg0IN_171, F(10)=>ImgReg0IN_170, F(9)=>
      ImgReg0IN_169, F(8)=>ImgReg0IN_168, F(7)=>ImgReg0IN_167, F(6)=>
      ImgReg0IN_166, F(5)=>ImgReg0IN_165, F(4)=>ImgReg0IN_164, F(3)=>
      ImgReg0IN_163, F(2)=>ImgReg0IN_162, F(1)=>ImgReg0IN_161, F(0)=>
      ImgReg0IN_160);
   loop3_10_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(175), 
      D(14)=>DATA(174), D(13)=>DATA(173), D(12)=>DATA(172), D(11)=>DATA(171), 
      D(10)=>DATA(170), D(9)=>DATA(169), D(8)=>DATA(168), D(7)=>DATA(167), 
      D(6)=>DATA(166), D(5)=>DATA(165), D(4)=>DATA(164), D(3)=>DATA(163), 
      D(2)=>DATA(162), D(1)=>DATA(161), D(0)=>DATA(160), EN=>nx23644, F(15)
      =>ImgReg1IN_175, F(14)=>ImgReg1IN_174, F(13)=>ImgReg1IN_173, F(12)=>
      ImgReg1IN_172, F(11)=>ImgReg1IN_171, F(10)=>ImgReg1IN_170, F(9)=>
      ImgReg1IN_169, F(8)=>ImgReg1IN_168, F(7)=>ImgReg1IN_167, F(6)=>
      ImgReg1IN_166, F(5)=>ImgReg1IN_165, F(4)=>ImgReg1IN_164, F(3)=>
      ImgReg1IN_163, F(2)=>ImgReg1IN_162, F(1)=>ImgReg1IN_161, F(0)=>
      ImgReg1IN_160);
   loop3_10_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(175), 
      D(14)=>DATA(174), D(13)=>DATA(173), D(12)=>DATA(172), D(11)=>DATA(171), 
      D(10)=>DATA(170), D(9)=>DATA(169), D(8)=>DATA(168), D(7)=>DATA(167), 
      D(6)=>DATA(166), D(5)=>DATA(165), D(4)=>DATA(164), D(3)=>DATA(163), 
      D(2)=>DATA(162), D(1)=>DATA(161), D(0)=>DATA(160), EN=>nx23632, F(15)
      =>ImgReg2IN_175, F(14)=>ImgReg2IN_174, F(13)=>ImgReg2IN_173, F(12)=>
      ImgReg2IN_172, F(11)=>ImgReg2IN_171, F(10)=>ImgReg2IN_170, F(9)=>
      ImgReg2IN_169, F(8)=>ImgReg2IN_168, F(7)=>ImgReg2IN_167, F(6)=>
      ImgReg2IN_166, F(5)=>ImgReg2IN_165, F(4)=>ImgReg2IN_164, F(3)=>
      ImgReg2IN_163, F(2)=>ImgReg2IN_162, F(1)=>ImgReg2IN_161, F(0)=>
      ImgReg2IN_160);
   loop3_10_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(175), 
      D(14)=>DATA(174), D(13)=>DATA(173), D(12)=>DATA(172), D(11)=>DATA(171), 
      D(10)=>DATA(170), D(9)=>DATA(169), D(8)=>DATA(168), D(7)=>DATA(167), 
      D(6)=>DATA(166), D(5)=>DATA(165), D(4)=>DATA(164), D(3)=>DATA(163), 
      D(2)=>DATA(162), D(1)=>DATA(161), D(0)=>DATA(160), EN=>nx23620, F(15)
      =>ImgReg3IN_175, F(14)=>ImgReg3IN_174, F(13)=>ImgReg3IN_173, F(12)=>
      ImgReg3IN_172, F(11)=>ImgReg3IN_171, F(10)=>ImgReg3IN_170, F(9)=>
      ImgReg3IN_169, F(8)=>ImgReg3IN_168, F(7)=>ImgReg3IN_167, F(6)=>
      ImgReg3IN_166, F(5)=>ImgReg3IN_165, F(4)=>ImgReg3IN_164, F(3)=>
      ImgReg3IN_163, F(2)=>ImgReg3IN_162, F(1)=>ImgReg3IN_161, F(0)=>
      ImgReg3IN_160);
   loop3_10_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(175), 
      D(14)=>DATA(174), D(13)=>DATA(173), D(12)=>DATA(172), D(11)=>DATA(171), 
      D(10)=>DATA(170), D(9)=>DATA(169), D(8)=>DATA(168), D(7)=>DATA(167), 
      D(6)=>DATA(166), D(5)=>DATA(165), D(4)=>DATA(164), D(3)=>DATA(163), 
      D(2)=>DATA(162), D(1)=>DATA(161), D(0)=>DATA(160), EN=>nx23608, F(15)
      =>ImgReg4IN_175, F(14)=>ImgReg4IN_174, F(13)=>ImgReg4IN_173, F(12)=>
      ImgReg4IN_172, F(11)=>ImgReg4IN_171, F(10)=>ImgReg4IN_170, F(9)=>
      ImgReg4IN_169, F(8)=>ImgReg4IN_168, F(7)=>ImgReg4IN_167, F(6)=>
      ImgReg4IN_166, F(5)=>ImgReg4IN_165, F(4)=>ImgReg4IN_164, F(3)=>
      ImgReg4IN_163, F(2)=>ImgReg4IN_162, F(1)=>ImgReg4IN_161, F(0)=>
      ImgReg4IN_160);
   loop3_10_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(175), 
      D(14)=>DATA(174), D(13)=>DATA(173), D(12)=>DATA(172), D(11)=>DATA(171), 
      D(10)=>DATA(170), D(9)=>DATA(169), D(8)=>DATA(168), D(7)=>DATA(167), 
      D(6)=>DATA(166), D(5)=>DATA(165), D(4)=>DATA(164), D(3)=>DATA(163), 
      D(2)=>DATA(162), D(1)=>DATA(161), D(0)=>DATA(160), EN=>nx23596, F(15)
      =>ImgReg5IN_175, F(14)=>ImgReg5IN_174, F(13)=>ImgReg5IN_173, F(12)=>
      ImgReg5IN_172, F(11)=>ImgReg5IN_171, F(10)=>ImgReg5IN_170, F(9)=>
      ImgReg5IN_169, F(8)=>ImgReg5IN_168, F(7)=>ImgReg5IN_167, F(6)=>
      ImgReg5IN_166, F(5)=>ImgReg5IN_165, F(4)=>ImgReg5IN_164, F(3)=>
      ImgReg5IN_163, F(2)=>ImgReg5IN_162, F(1)=>ImgReg5IN_161, F(0)=>
      ImgReg5IN_160);
   loop3_10_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_175_EXMPLR, D(14)=>OutputImg1_174_EXMPLR, D(13)=>
      OutputImg1_173_EXMPLR, D(12)=>OutputImg1_172_EXMPLR, D(11)=>
      OutputImg1_171_EXMPLR, D(10)=>OutputImg1_170_EXMPLR, D(9)=>
      OutputImg1_169_EXMPLR, D(8)=>OutputImg1_168_EXMPLR, D(7)=>
      OutputImg1_167_EXMPLR, D(6)=>OutputImg1_166_EXMPLR, D(5)=>
      OutputImg1_165_EXMPLR, D(4)=>OutputImg1_164_EXMPLR, D(3)=>
      OutputImg1_163_EXMPLR, D(2)=>OutputImg1_162_EXMPLR, D(1)=>
      OutputImg1_161_EXMPLR, D(0)=>OutputImg1_160_EXMPLR, EN=>nx23800, F(15)
      =>ImgReg0IN_175, F(14)=>ImgReg0IN_174, F(13)=>ImgReg0IN_173, F(12)=>
      ImgReg0IN_172, F(11)=>ImgReg0IN_171, F(10)=>ImgReg0IN_170, F(9)=>
      ImgReg0IN_169, F(8)=>ImgReg0IN_168, F(7)=>ImgReg0IN_167, F(6)=>
      ImgReg0IN_166, F(5)=>ImgReg0IN_165, F(4)=>ImgReg0IN_164, F(3)=>
      ImgReg0IN_163, F(2)=>ImgReg0IN_162, F(1)=>ImgReg0IN_161, F(0)=>
      ImgReg0IN_160);
   loop3_10_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_175_EXMPLR, D(14)=>OutputImg2_174_EXMPLR, D(13)=>
      OutputImg2_173_EXMPLR, D(12)=>OutputImg2_172_EXMPLR, D(11)=>
      OutputImg2_171_EXMPLR, D(10)=>OutputImg2_170_EXMPLR, D(9)=>
      OutputImg2_169_EXMPLR, D(8)=>OutputImg2_168_EXMPLR, D(7)=>
      OutputImg2_167_EXMPLR, D(6)=>OutputImg2_166_EXMPLR, D(5)=>
      OutputImg2_165_EXMPLR, D(4)=>OutputImg2_164_EXMPLR, D(3)=>
      OutputImg2_163_EXMPLR, D(2)=>OutputImg2_162_EXMPLR, D(1)=>
      OutputImg2_161_EXMPLR, D(0)=>OutputImg2_160_EXMPLR, EN=>nx23800, F(15)
      =>ImgReg1IN_175, F(14)=>ImgReg1IN_174, F(13)=>ImgReg1IN_173, F(12)=>
      ImgReg1IN_172, F(11)=>ImgReg1IN_171, F(10)=>ImgReg1IN_170, F(9)=>
      ImgReg1IN_169, F(8)=>ImgReg1IN_168, F(7)=>ImgReg1IN_167, F(6)=>
      ImgReg1IN_166, F(5)=>ImgReg1IN_165, F(4)=>ImgReg1IN_164, F(3)=>
      ImgReg1IN_163, F(2)=>ImgReg1IN_162, F(1)=>ImgReg1IN_161, F(0)=>
      ImgReg1IN_160);
   loop3_10_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_175_EXMPLR, D(14)=>OutputImg3_174_EXMPLR, D(13)=>
      OutputImg3_173_EXMPLR, D(12)=>OutputImg3_172_EXMPLR, D(11)=>
      OutputImg3_171_EXMPLR, D(10)=>OutputImg3_170_EXMPLR, D(9)=>
      OutputImg3_169_EXMPLR, D(8)=>OutputImg3_168_EXMPLR, D(7)=>
      OutputImg3_167_EXMPLR, D(6)=>OutputImg3_166_EXMPLR, D(5)=>
      OutputImg3_165_EXMPLR, D(4)=>OutputImg3_164_EXMPLR, D(3)=>
      OutputImg3_163_EXMPLR, D(2)=>OutputImg3_162_EXMPLR, D(1)=>
      OutputImg3_161_EXMPLR, D(0)=>OutputImg3_160_EXMPLR, EN=>nx23800, F(15)
      =>ImgReg2IN_175, F(14)=>ImgReg2IN_174, F(13)=>ImgReg2IN_173, F(12)=>
      ImgReg2IN_172, F(11)=>ImgReg2IN_171, F(10)=>ImgReg2IN_170, F(9)=>
      ImgReg2IN_169, F(8)=>ImgReg2IN_168, F(7)=>ImgReg2IN_167, F(6)=>
      ImgReg2IN_166, F(5)=>ImgReg2IN_165, F(4)=>ImgReg2IN_164, F(3)=>
      ImgReg2IN_163, F(2)=>ImgReg2IN_162, F(1)=>ImgReg2IN_161, F(0)=>
      ImgReg2IN_160);
   loop3_10_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_175_EXMPLR, D(14)=>OutputImg4_174_EXMPLR, D(13)=>
      OutputImg4_173_EXMPLR, D(12)=>OutputImg4_172_EXMPLR, D(11)=>
      OutputImg4_171_EXMPLR, D(10)=>OutputImg4_170_EXMPLR, D(9)=>
      OutputImg4_169_EXMPLR, D(8)=>OutputImg4_168_EXMPLR, D(7)=>
      OutputImg4_167_EXMPLR, D(6)=>OutputImg4_166_EXMPLR, D(5)=>
      OutputImg4_165_EXMPLR, D(4)=>OutputImg4_164_EXMPLR, D(3)=>
      OutputImg4_163_EXMPLR, D(2)=>OutputImg4_162_EXMPLR, D(1)=>
      OutputImg4_161_EXMPLR, D(0)=>OutputImg4_160_EXMPLR, EN=>nx23800, F(15)
      =>ImgReg3IN_175, F(14)=>ImgReg3IN_174, F(13)=>ImgReg3IN_173, F(12)=>
      ImgReg3IN_172, F(11)=>ImgReg3IN_171, F(10)=>ImgReg3IN_170, F(9)=>
      ImgReg3IN_169, F(8)=>ImgReg3IN_168, F(7)=>ImgReg3IN_167, F(6)=>
      ImgReg3IN_166, F(5)=>ImgReg3IN_165, F(4)=>ImgReg3IN_164, F(3)=>
      ImgReg3IN_163, F(2)=>ImgReg3IN_162, F(1)=>ImgReg3IN_161, F(0)=>
      ImgReg3IN_160);
   loop3_10_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_175_EXMPLR, D(14)=>OutputImg5_174_EXMPLR, D(13)=>
      OutputImg5_173_EXMPLR, D(12)=>OutputImg5_172_EXMPLR, D(11)=>
      OutputImg5_171_EXMPLR, D(10)=>OutputImg5_170_EXMPLR, D(9)=>
      OutputImg5_169_EXMPLR, D(8)=>OutputImg5_168_EXMPLR, D(7)=>
      OutputImg5_167_EXMPLR, D(6)=>OutputImg5_166_EXMPLR, D(5)=>
      OutputImg5_165_EXMPLR, D(4)=>OutputImg5_164_EXMPLR, D(3)=>
      OutputImg5_163_EXMPLR, D(2)=>OutputImg5_162_EXMPLR, D(1)=>
      OutputImg5_161_EXMPLR, D(0)=>OutputImg5_160_EXMPLR, EN=>nx23800, F(15)
      =>ImgReg4IN_175, F(14)=>ImgReg4IN_174, F(13)=>ImgReg4IN_173, F(12)=>
      ImgReg4IN_172, F(11)=>ImgReg4IN_171, F(10)=>ImgReg4IN_170, F(9)=>
      ImgReg4IN_169, F(8)=>ImgReg4IN_168, F(7)=>ImgReg4IN_167, F(6)=>
      ImgReg4IN_166, F(5)=>ImgReg4IN_165, F(4)=>ImgReg4IN_164, F(3)=>
      ImgReg4IN_163, F(2)=>ImgReg4IN_162, F(1)=>ImgReg4IN_161, F(0)=>
      ImgReg4IN_160);
   loop3_10_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_175, D(14)=>
      ImgReg0IN_174, D(13)=>ImgReg0IN_173, D(12)=>ImgReg0IN_172, D(11)=>
      ImgReg0IN_171, D(10)=>ImgReg0IN_170, D(9)=>ImgReg0IN_169, D(8)=>
      ImgReg0IN_168, D(7)=>ImgReg0IN_167, D(6)=>ImgReg0IN_166, D(5)=>
      ImgReg0IN_165, D(4)=>ImgReg0IN_164, D(3)=>ImgReg0IN_163, D(2)=>
      ImgReg0IN_162, D(1)=>ImgReg0IN_161, D(0)=>ImgReg0IN_160, CLK=>nx23888, 
      RST=>RST, EN=>nx23720, Q(15)=>OutputImg0_175_EXMPLR, Q(14)=>
      OutputImg0_174_EXMPLR, Q(13)=>OutputImg0_173_EXMPLR, Q(12)=>
      OutputImg0_172_EXMPLR, Q(11)=>OutputImg0_171_EXMPLR, Q(10)=>
      OutputImg0_170_EXMPLR, Q(9)=>OutputImg0_169_EXMPLR, Q(8)=>
      OutputImg0_168_EXMPLR, Q(7)=>OutputImg0_167_EXMPLR, Q(6)=>
      OutputImg0_166_EXMPLR, Q(5)=>OutputImg0_165_EXMPLR, Q(4)=>
      OutputImg0_164_EXMPLR, Q(3)=>OutputImg0_163_EXMPLR, Q(2)=>
      OutputImg0_162_EXMPLR, Q(1)=>OutputImg0_161_EXMPLR, Q(0)=>
      OutputImg0_160_EXMPLR);
   loop3_10_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_175, D(14)=>
      ImgReg1IN_174, D(13)=>ImgReg1IN_173, D(12)=>ImgReg1IN_172, D(11)=>
      ImgReg1IN_171, D(10)=>ImgReg1IN_170, D(9)=>ImgReg1IN_169, D(8)=>
      ImgReg1IN_168, D(7)=>ImgReg1IN_167, D(6)=>ImgReg1IN_166, D(5)=>
      ImgReg1IN_165, D(4)=>ImgReg1IN_164, D(3)=>ImgReg1IN_163, D(2)=>
      ImgReg1IN_162, D(1)=>ImgReg1IN_161, D(0)=>ImgReg1IN_160, CLK=>nx23890, 
      RST=>RST, EN=>nx23730, Q(15)=>OutputImg1_175_EXMPLR, Q(14)=>
      OutputImg1_174_EXMPLR, Q(13)=>OutputImg1_173_EXMPLR, Q(12)=>
      OutputImg1_172_EXMPLR, Q(11)=>OutputImg1_171_EXMPLR, Q(10)=>
      OutputImg1_170_EXMPLR, Q(9)=>OutputImg1_169_EXMPLR, Q(8)=>
      OutputImg1_168_EXMPLR, Q(7)=>OutputImg1_167_EXMPLR, Q(6)=>
      OutputImg1_166_EXMPLR, Q(5)=>OutputImg1_165_EXMPLR, Q(4)=>
      OutputImg1_164_EXMPLR, Q(3)=>OutputImg1_163_EXMPLR, Q(2)=>
      OutputImg1_162_EXMPLR, Q(1)=>OutputImg1_161_EXMPLR, Q(0)=>
      OutputImg1_160_EXMPLR);
   loop3_10_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_175, D(14)=>
      ImgReg2IN_174, D(13)=>ImgReg2IN_173, D(12)=>ImgReg2IN_172, D(11)=>
      ImgReg2IN_171, D(10)=>ImgReg2IN_170, D(9)=>ImgReg2IN_169, D(8)=>
      ImgReg2IN_168, D(7)=>ImgReg2IN_167, D(6)=>ImgReg2IN_166, D(5)=>
      ImgReg2IN_165, D(4)=>ImgReg2IN_164, D(3)=>ImgReg2IN_163, D(2)=>
      ImgReg2IN_162, D(1)=>ImgReg2IN_161, D(0)=>ImgReg2IN_160, CLK=>nx23890, 
      RST=>RST, EN=>nx23740, Q(15)=>OutputImg2_175_EXMPLR, Q(14)=>
      OutputImg2_174_EXMPLR, Q(13)=>OutputImg2_173_EXMPLR, Q(12)=>
      OutputImg2_172_EXMPLR, Q(11)=>OutputImg2_171_EXMPLR, Q(10)=>
      OutputImg2_170_EXMPLR, Q(9)=>OutputImg2_169_EXMPLR, Q(8)=>
      OutputImg2_168_EXMPLR, Q(7)=>OutputImg2_167_EXMPLR, Q(6)=>
      OutputImg2_166_EXMPLR, Q(5)=>OutputImg2_165_EXMPLR, Q(4)=>
      OutputImg2_164_EXMPLR, Q(3)=>OutputImg2_163_EXMPLR, Q(2)=>
      OutputImg2_162_EXMPLR, Q(1)=>OutputImg2_161_EXMPLR, Q(0)=>
      OutputImg2_160_EXMPLR);
   loop3_10_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_175, D(14)=>
      ImgReg3IN_174, D(13)=>ImgReg3IN_173, D(12)=>ImgReg3IN_172, D(11)=>
      ImgReg3IN_171, D(10)=>ImgReg3IN_170, D(9)=>ImgReg3IN_169, D(8)=>
      ImgReg3IN_168, D(7)=>ImgReg3IN_167, D(6)=>ImgReg3IN_166, D(5)=>
      ImgReg3IN_165, D(4)=>ImgReg3IN_164, D(3)=>ImgReg3IN_163, D(2)=>
      ImgReg3IN_162, D(1)=>ImgReg3IN_161, D(0)=>ImgReg3IN_160, CLK=>nx23892, 
      RST=>RST, EN=>nx23750, Q(15)=>OutputImg3_175_EXMPLR, Q(14)=>
      OutputImg3_174_EXMPLR, Q(13)=>OutputImg3_173_EXMPLR, Q(12)=>
      OutputImg3_172_EXMPLR, Q(11)=>OutputImg3_171_EXMPLR, Q(10)=>
      OutputImg3_170_EXMPLR, Q(9)=>OutputImg3_169_EXMPLR, Q(8)=>
      OutputImg3_168_EXMPLR, Q(7)=>OutputImg3_167_EXMPLR, Q(6)=>
      OutputImg3_166_EXMPLR, Q(5)=>OutputImg3_165_EXMPLR, Q(4)=>
      OutputImg3_164_EXMPLR, Q(3)=>OutputImg3_163_EXMPLR, Q(2)=>
      OutputImg3_162_EXMPLR, Q(1)=>OutputImg3_161_EXMPLR, Q(0)=>
      OutputImg3_160_EXMPLR);
   loop3_10_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_175, D(14)=>
      ImgReg4IN_174, D(13)=>ImgReg4IN_173, D(12)=>ImgReg4IN_172, D(11)=>
      ImgReg4IN_171, D(10)=>ImgReg4IN_170, D(9)=>ImgReg4IN_169, D(8)=>
      ImgReg4IN_168, D(7)=>ImgReg4IN_167, D(6)=>ImgReg4IN_166, D(5)=>
      ImgReg4IN_165, D(4)=>ImgReg4IN_164, D(3)=>ImgReg4IN_163, D(2)=>
      ImgReg4IN_162, D(1)=>ImgReg4IN_161, D(0)=>ImgReg4IN_160, CLK=>nx23892, 
      RST=>RST, EN=>nx23760, Q(15)=>OutputImg4_175_EXMPLR, Q(14)=>
      OutputImg4_174_EXMPLR, Q(13)=>OutputImg4_173_EXMPLR, Q(12)=>
      OutputImg4_172_EXMPLR, Q(11)=>OutputImg4_171_EXMPLR, Q(10)=>
      OutputImg4_170_EXMPLR, Q(9)=>OutputImg4_169_EXMPLR, Q(8)=>
      OutputImg4_168_EXMPLR, Q(7)=>OutputImg4_167_EXMPLR, Q(6)=>
      OutputImg4_166_EXMPLR, Q(5)=>OutputImg4_165_EXMPLR, Q(4)=>
      OutputImg4_164_EXMPLR, Q(3)=>OutputImg4_163_EXMPLR, Q(2)=>
      OutputImg4_162_EXMPLR, Q(1)=>OutputImg4_161_EXMPLR, Q(0)=>
      OutputImg4_160_EXMPLR);
   loop3_10_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_175, D(14)=>
      ImgReg5IN_174, D(13)=>ImgReg5IN_173, D(12)=>ImgReg5IN_172, D(11)=>
      ImgReg5IN_171, D(10)=>ImgReg5IN_170, D(9)=>ImgReg5IN_169, D(8)=>
      ImgReg5IN_168, D(7)=>ImgReg5IN_167, D(6)=>ImgReg5IN_166, D(5)=>
      ImgReg5IN_165, D(4)=>ImgReg5IN_164, D(3)=>ImgReg5IN_163, D(2)=>
      ImgReg5IN_162, D(1)=>ImgReg5IN_161, D(0)=>ImgReg5IN_160, CLK=>nx23894, 
      RST=>RST, EN=>nx23770, Q(15)=>OutputImg5_175_EXMPLR, Q(14)=>
      OutputImg5_174_EXMPLR, Q(13)=>OutputImg5_173_EXMPLR, Q(12)=>
      OutputImg5_172_EXMPLR, Q(11)=>OutputImg5_171_EXMPLR, Q(10)=>
      OutputImg5_170_EXMPLR, Q(9)=>OutputImg5_169_EXMPLR, Q(8)=>
      OutputImg5_168_EXMPLR, Q(7)=>OutputImg5_167_EXMPLR, Q(6)=>
      OutputImg5_166_EXMPLR, Q(5)=>OutputImg5_165_EXMPLR, Q(4)=>
      OutputImg5_164_EXMPLR, Q(3)=>OutputImg5_163_EXMPLR, Q(2)=>
      OutputImg5_162_EXMPLR, Q(1)=>OutputImg5_161_EXMPLR, Q(0)=>
      OutputImg5_160_EXMPLR);
   loop3_11_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_207_EXMPLR, D(14)=>OutputImg0_206_EXMPLR, D(13)=>
      OutputImg0_205_EXMPLR, D(12)=>OutputImg0_204_EXMPLR, D(11)=>
      OutputImg0_203_EXMPLR, D(10)=>OutputImg0_202_EXMPLR, D(9)=>
      OutputImg0_201_EXMPLR, D(8)=>OutputImg0_200_EXMPLR, D(7)=>
      OutputImg0_199_EXMPLR, D(6)=>OutputImg0_198_EXMPLR, D(5)=>
      OutputImg0_197_EXMPLR, D(4)=>OutputImg0_196_EXMPLR, D(3)=>
      OutputImg0_195_EXMPLR, D(2)=>OutputImg0_194_EXMPLR, D(1)=>
      OutputImg0_193_EXMPLR, D(0)=>OutputImg0_192_EXMPLR, EN=>nx23684, F(15)
      =>ImgReg0IN_191, F(14)=>ImgReg0IN_190, F(13)=>ImgReg0IN_189, F(12)=>
      ImgReg0IN_188, F(11)=>ImgReg0IN_187, F(10)=>ImgReg0IN_186, F(9)=>
      ImgReg0IN_185, F(8)=>ImgReg0IN_184, F(7)=>ImgReg0IN_183, F(6)=>
      ImgReg0IN_182, F(5)=>ImgReg0IN_181, F(4)=>ImgReg0IN_180, F(3)=>
      ImgReg0IN_179, F(2)=>ImgReg0IN_178, F(1)=>ImgReg0IN_177, F(0)=>
      ImgReg0IN_176);
   loop3_11_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_207_EXMPLR, D(14)=>OutputImg1_206_EXMPLR, D(13)=>
      OutputImg1_205_EXMPLR, D(12)=>OutputImg1_204_EXMPLR, D(11)=>
      OutputImg1_203_EXMPLR, D(10)=>OutputImg1_202_EXMPLR, D(9)=>
      OutputImg1_201_EXMPLR, D(8)=>OutputImg1_200_EXMPLR, D(7)=>
      OutputImg1_199_EXMPLR, D(6)=>OutputImg1_198_EXMPLR, D(5)=>
      OutputImg1_197_EXMPLR, D(4)=>OutputImg1_196_EXMPLR, D(3)=>
      OutputImg1_195_EXMPLR, D(2)=>OutputImg1_194_EXMPLR, D(1)=>
      OutputImg1_193_EXMPLR, D(0)=>OutputImg1_192_EXMPLR, EN=>nx23684, F(15)
      =>ImgReg1IN_191, F(14)=>ImgReg1IN_190, F(13)=>ImgReg1IN_189, F(12)=>
      ImgReg1IN_188, F(11)=>ImgReg1IN_187, F(10)=>ImgReg1IN_186, F(9)=>
      ImgReg1IN_185, F(8)=>ImgReg1IN_184, F(7)=>ImgReg1IN_183, F(6)=>
      ImgReg1IN_182, F(5)=>ImgReg1IN_181, F(4)=>ImgReg1IN_180, F(3)=>
      ImgReg1IN_179, F(2)=>ImgReg1IN_178, F(1)=>ImgReg1IN_177, F(0)=>
      ImgReg1IN_176);
   loop3_11_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_207_EXMPLR, D(14)=>OutputImg2_206_EXMPLR, D(13)=>
      OutputImg2_205_EXMPLR, D(12)=>OutputImg2_204_EXMPLR, D(11)=>
      OutputImg2_203_EXMPLR, D(10)=>OutputImg2_202_EXMPLR, D(9)=>
      OutputImg2_201_EXMPLR, D(8)=>OutputImg2_200_EXMPLR, D(7)=>
      OutputImg2_199_EXMPLR, D(6)=>OutputImg2_198_EXMPLR, D(5)=>
      OutputImg2_197_EXMPLR, D(4)=>OutputImg2_196_EXMPLR, D(3)=>
      OutputImg2_195_EXMPLR, D(2)=>OutputImg2_194_EXMPLR, D(1)=>
      OutputImg2_193_EXMPLR, D(0)=>OutputImg2_192_EXMPLR, EN=>nx23684, F(15)
      =>ImgReg2IN_191, F(14)=>ImgReg2IN_190, F(13)=>ImgReg2IN_189, F(12)=>
      ImgReg2IN_188, F(11)=>ImgReg2IN_187, F(10)=>ImgReg2IN_186, F(9)=>
      ImgReg2IN_185, F(8)=>ImgReg2IN_184, F(7)=>ImgReg2IN_183, F(6)=>
      ImgReg2IN_182, F(5)=>ImgReg2IN_181, F(4)=>ImgReg2IN_180, F(3)=>
      ImgReg2IN_179, F(2)=>ImgReg2IN_178, F(1)=>ImgReg2IN_177, F(0)=>
      ImgReg2IN_176);
   loop3_11_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_207_EXMPLR, D(14)=>OutputImg3_206_EXMPLR, D(13)=>
      OutputImg3_205_EXMPLR, D(12)=>OutputImg3_204_EXMPLR, D(11)=>
      OutputImg3_203_EXMPLR, D(10)=>OutputImg3_202_EXMPLR, D(9)=>
      OutputImg3_201_EXMPLR, D(8)=>OutputImg3_200_EXMPLR, D(7)=>
      OutputImg3_199_EXMPLR, D(6)=>OutputImg3_198_EXMPLR, D(5)=>
      OutputImg3_197_EXMPLR, D(4)=>OutputImg3_196_EXMPLR, D(3)=>
      OutputImg3_195_EXMPLR, D(2)=>OutputImg3_194_EXMPLR, D(1)=>
      OutputImg3_193_EXMPLR, D(0)=>OutputImg3_192_EXMPLR, EN=>nx23684, F(15)
      =>ImgReg3IN_191, F(14)=>ImgReg3IN_190, F(13)=>ImgReg3IN_189, F(12)=>
      ImgReg3IN_188, F(11)=>ImgReg3IN_187, F(10)=>ImgReg3IN_186, F(9)=>
      ImgReg3IN_185, F(8)=>ImgReg3IN_184, F(7)=>ImgReg3IN_183, F(6)=>
      ImgReg3IN_182, F(5)=>ImgReg3IN_181, F(4)=>ImgReg3IN_180, F(3)=>
      ImgReg3IN_179, F(2)=>ImgReg3IN_178, F(1)=>ImgReg3IN_177, F(0)=>
      ImgReg3IN_176);
   loop3_11_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_207_EXMPLR, D(14)=>OutputImg4_206_EXMPLR, D(13)=>
      OutputImg4_205_EXMPLR, D(12)=>OutputImg4_204_EXMPLR, D(11)=>
      OutputImg4_203_EXMPLR, D(10)=>OutputImg4_202_EXMPLR, D(9)=>
      OutputImg4_201_EXMPLR, D(8)=>OutputImg4_200_EXMPLR, D(7)=>
      OutputImg4_199_EXMPLR, D(6)=>OutputImg4_198_EXMPLR, D(5)=>
      OutputImg4_197_EXMPLR, D(4)=>OutputImg4_196_EXMPLR, D(3)=>
      OutputImg4_195_EXMPLR, D(2)=>OutputImg4_194_EXMPLR, D(1)=>
      OutputImg4_193_EXMPLR, D(0)=>OutputImg4_192_EXMPLR, EN=>nx23686, F(15)
      =>ImgReg4IN_191, F(14)=>ImgReg4IN_190, F(13)=>ImgReg4IN_189, F(12)=>
      ImgReg4IN_188, F(11)=>ImgReg4IN_187, F(10)=>ImgReg4IN_186, F(9)=>
      ImgReg4IN_185, F(8)=>ImgReg4IN_184, F(7)=>ImgReg4IN_183, F(6)=>
      ImgReg4IN_182, F(5)=>ImgReg4IN_181, F(4)=>ImgReg4IN_180, F(3)=>
      ImgReg4IN_179, F(2)=>ImgReg4IN_178, F(1)=>ImgReg4IN_177, F(0)=>
      ImgReg4IN_176);
   loop3_11_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_207_EXMPLR, D(14)=>OutputImg5_206_EXMPLR, D(13)=>
      OutputImg5_205_EXMPLR, D(12)=>OutputImg5_204_EXMPLR, D(11)=>
      OutputImg5_203_EXMPLR, D(10)=>OutputImg5_202_EXMPLR, D(9)=>
      OutputImg5_201_EXMPLR, D(8)=>OutputImg5_200_EXMPLR, D(7)=>
      OutputImg5_199_EXMPLR, D(6)=>OutputImg5_198_EXMPLR, D(5)=>
      OutputImg5_197_EXMPLR, D(4)=>OutputImg5_196_EXMPLR, D(3)=>
      OutputImg5_195_EXMPLR, D(2)=>OutputImg5_194_EXMPLR, D(1)=>
      OutputImg5_193_EXMPLR, D(0)=>OutputImg5_192_EXMPLR, EN=>nx23686, F(15)
      =>ImgReg5IN_191, F(14)=>ImgReg5IN_190, F(13)=>ImgReg5IN_189, F(12)=>
      ImgReg5IN_188, F(11)=>ImgReg5IN_187, F(10)=>ImgReg5IN_186, F(9)=>
      ImgReg5IN_185, F(8)=>ImgReg5IN_184, F(7)=>ImgReg5IN_183, F(6)=>
      ImgReg5IN_182, F(5)=>ImgReg5IN_181, F(4)=>ImgReg5IN_180, F(3)=>
      ImgReg5IN_179, F(2)=>ImgReg5IN_178, F(1)=>ImgReg5IN_177, F(0)=>
      ImgReg5IN_176);
   loop3_11_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(191), 
      D(14)=>DATA(190), D(13)=>DATA(189), D(12)=>DATA(188), D(11)=>DATA(187), 
      D(10)=>DATA(186), D(9)=>DATA(185), D(8)=>DATA(184), D(7)=>DATA(183), 
      D(6)=>DATA(182), D(5)=>DATA(181), D(4)=>DATA(180), D(3)=>DATA(179), 
      D(2)=>DATA(178), D(1)=>DATA(177), D(0)=>DATA(176), EN=>nx23656, F(15)
      =>ImgReg0IN_191, F(14)=>ImgReg0IN_190, F(13)=>ImgReg0IN_189, F(12)=>
      ImgReg0IN_188, F(11)=>ImgReg0IN_187, F(10)=>ImgReg0IN_186, F(9)=>
      ImgReg0IN_185, F(8)=>ImgReg0IN_184, F(7)=>ImgReg0IN_183, F(6)=>
      ImgReg0IN_182, F(5)=>ImgReg0IN_181, F(4)=>ImgReg0IN_180, F(3)=>
      ImgReg0IN_179, F(2)=>ImgReg0IN_178, F(1)=>ImgReg0IN_177, F(0)=>
      ImgReg0IN_176);
   loop3_11_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(191), 
      D(14)=>DATA(190), D(13)=>DATA(189), D(12)=>DATA(188), D(11)=>DATA(187), 
      D(10)=>DATA(186), D(9)=>DATA(185), D(8)=>DATA(184), D(7)=>DATA(183), 
      D(6)=>DATA(182), D(5)=>DATA(181), D(4)=>DATA(180), D(3)=>DATA(179), 
      D(2)=>DATA(178), D(1)=>DATA(177), D(0)=>DATA(176), EN=>nx23644, F(15)
      =>ImgReg1IN_191, F(14)=>ImgReg1IN_190, F(13)=>ImgReg1IN_189, F(12)=>
      ImgReg1IN_188, F(11)=>ImgReg1IN_187, F(10)=>ImgReg1IN_186, F(9)=>
      ImgReg1IN_185, F(8)=>ImgReg1IN_184, F(7)=>ImgReg1IN_183, F(6)=>
      ImgReg1IN_182, F(5)=>ImgReg1IN_181, F(4)=>ImgReg1IN_180, F(3)=>
      ImgReg1IN_179, F(2)=>ImgReg1IN_178, F(1)=>ImgReg1IN_177, F(0)=>
      ImgReg1IN_176);
   loop3_11_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(191), 
      D(14)=>DATA(190), D(13)=>DATA(189), D(12)=>DATA(188), D(11)=>DATA(187), 
      D(10)=>DATA(186), D(9)=>DATA(185), D(8)=>DATA(184), D(7)=>DATA(183), 
      D(6)=>DATA(182), D(5)=>DATA(181), D(4)=>DATA(180), D(3)=>DATA(179), 
      D(2)=>DATA(178), D(1)=>DATA(177), D(0)=>DATA(176), EN=>nx23632, F(15)
      =>ImgReg2IN_191, F(14)=>ImgReg2IN_190, F(13)=>ImgReg2IN_189, F(12)=>
      ImgReg2IN_188, F(11)=>ImgReg2IN_187, F(10)=>ImgReg2IN_186, F(9)=>
      ImgReg2IN_185, F(8)=>ImgReg2IN_184, F(7)=>ImgReg2IN_183, F(6)=>
      ImgReg2IN_182, F(5)=>ImgReg2IN_181, F(4)=>ImgReg2IN_180, F(3)=>
      ImgReg2IN_179, F(2)=>ImgReg2IN_178, F(1)=>ImgReg2IN_177, F(0)=>
      ImgReg2IN_176);
   loop3_11_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(191), 
      D(14)=>DATA(190), D(13)=>DATA(189), D(12)=>DATA(188), D(11)=>DATA(187), 
      D(10)=>DATA(186), D(9)=>DATA(185), D(8)=>DATA(184), D(7)=>DATA(183), 
      D(6)=>DATA(182), D(5)=>DATA(181), D(4)=>DATA(180), D(3)=>DATA(179), 
      D(2)=>DATA(178), D(1)=>DATA(177), D(0)=>DATA(176), EN=>nx23620, F(15)
      =>ImgReg3IN_191, F(14)=>ImgReg3IN_190, F(13)=>ImgReg3IN_189, F(12)=>
      ImgReg3IN_188, F(11)=>ImgReg3IN_187, F(10)=>ImgReg3IN_186, F(9)=>
      ImgReg3IN_185, F(8)=>ImgReg3IN_184, F(7)=>ImgReg3IN_183, F(6)=>
      ImgReg3IN_182, F(5)=>ImgReg3IN_181, F(4)=>ImgReg3IN_180, F(3)=>
      ImgReg3IN_179, F(2)=>ImgReg3IN_178, F(1)=>ImgReg3IN_177, F(0)=>
      ImgReg3IN_176);
   loop3_11_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(191), 
      D(14)=>DATA(190), D(13)=>DATA(189), D(12)=>DATA(188), D(11)=>DATA(187), 
      D(10)=>DATA(186), D(9)=>DATA(185), D(8)=>DATA(184), D(7)=>DATA(183), 
      D(6)=>DATA(182), D(5)=>DATA(181), D(4)=>DATA(180), D(3)=>DATA(179), 
      D(2)=>DATA(178), D(1)=>DATA(177), D(0)=>DATA(176), EN=>nx23608, F(15)
      =>ImgReg4IN_191, F(14)=>ImgReg4IN_190, F(13)=>ImgReg4IN_189, F(12)=>
      ImgReg4IN_188, F(11)=>ImgReg4IN_187, F(10)=>ImgReg4IN_186, F(9)=>
      ImgReg4IN_185, F(8)=>ImgReg4IN_184, F(7)=>ImgReg4IN_183, F(6)=>
      ImgReg4IN_182, F(5)=>ImgReg4IN_181, F(4)=>ImgReg4IN_180, F(3)=>
      ImgReg4IN_179, F(2)=>ImgReg4IN_178, F(1)=>ImgReg4IN_177, F(0)=>
      ImgReg4IN_176);
   loop3_11_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(191), 
      D(14)=>DATA(190), D(13)=>DATA(189), D(12)=>DATA(188), D(11)=>DATA(187), 
      D(10)=>DATA(186), D(9)=>DATA(185), D(8)=>DATA(184), D(7)=>DATA(183), 
      D(6)=>DATA(182), D(5)=>DATA(181), D(4)=>DATA(180), D(3)=>DATA(179), 
      D(2)=>DATA(178), D(1)=>DATA(177), D(0)=>DATA(176), EN=>nx23596, F(15)
      =>ImgReg5IN_191, F(14)=>ImgReg5IN_190, F(13)=>ImgReg5IN_189, F(12)=>
      ImgReg5IN_188, F(11)=>ImgReg5IN_187, F(10)=>ImgReg5IN_186, F(9)=>
      ImgReg5IN_185, F(8)=>ImgReg5IN_184, F(7)=>ImgReg5IN_183, F(6)=>
      ImgReg5IN_182, F(5)=>ImgReg5IN_181, F(4)=>ImgReg5IN_180, F(3)=>
      ImgReg5IN_179, F(2)=>ImgReg5IN_178, F(1)=>ImgReg5IN_177, F(0)=>
      ImgReg5IN_176);
   loop3_11_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_191_EXMPLR, D(14)=>OutputImg1_190_EXMPLR, D(13)=>
      OutputImg1_189_EXMPLR, D(12)=>OutputImg1_188_EXMPLR, D(11)=>
      OutputImg1_187_EXMPLR, D(10)=>OutputImg1_186_EXMPLR, D(9)=>
      OutputImg1_185_EXMPLR, D(8)=>OutputImg1_184_EXMPLR, D(7)=>
      OutputImg1_183_EXMPLR, D(6)=>OutputImg1_182_EXMPLR, D(5)=>
      OutputImg1_181_EXMPLR, D(4)=>OutputImg1_180_EXMPLR, D(3)=>
      OutputImg1_179_EXMPLR, D(2)=>OutputImg1_178_EXMPLR, D(1)=>
      OutputImg1_177_EXMPLR, D(0)=>OutputImg1_176_EXMPLR, EN=>nx23800, F(15)
      =>ImgReg0IN_191, F(14)=>ImgReg0IN_190, F(13)=>ImgReg0IN_189, F(12)=>
      ImgReg0IN_188, F(11)=>ImgReg0IN_187, F(10)=>ImgReg0IN_186, F(9)=>
      ImgReg0IN_185, F(8)=>ImgReg0IN_184, F(7)=>ImgReg0IN_183, F(6)=>
      ImgReg0IN_182, F(5)=>ImgReg0IN_181, F(4)=>ImgReg0IN_180, F(3)=>
      ImgReg0IN_179, F(2)=>ImgReg0IN_178, F(1)=>ImgReg0IN_177, F(0)=>
      ImgReg0IN_176);
   loop3_11_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_191_EXMPLR, D(14)=>OutputImg2_190_EXMPLR, D(13)=>
      OutputImg2_189_EXMPLR, D(12)=>OutputImg2_188_EXMPLR, D(11)=>
      OutputImg2_187_EXMPLR, D(10)=>OutputImg2_186_EXMPLR, D(9)=>
      OutputImg2_185_EXMPLR, D(8)=>OutputImg2_184_EXMPLR, D(7)=>
      OutputImg2_183_EXMPLR, D(6)=>OutputImg2_182_EXMPLR, D(5)=>
      OutputImg2_181_EXMPLR, D(4)=>OutputImg2_180_EXMPLR, D(3)=>
      OutputImg2_179_EXMPLR, D(2)=>OutputImg2_178_EXMPLR, D(1)=>
      OutputImg2_177_EXMPLR, D(0)=>OutputImg2_176_EXMPLR, EN=>nx23802, F(15)
      =>ImgReg1IN_191, F(14)=>ImgReg1IN_190, F(13)=>ImgReg1IN_189, F(12)=>
      ImgReg1IN_188, F(11)=>ImgReg1IN_187, F(10)=>ImgReg1IN_186, F(9)=>
      ImgReg1IN_185, F(8)=>ImgReg1IN_184, F(7)=>ImgReg1IN_183, F(6)=>
      ImgReg1IN_182, F(5)=>ImgReg1IN_181, F(4)=>ImgReg1IN_180, F(3)=>
      ImgReg1IN_179, F(2)=>ImgReg1IN_178, F(1)=>ImgReg1IN_177, F(0)=>
      ImgReg1IN_176);
   loop3_11_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_191_EXMPLR, D(14)=>OutputImg3_190_EXMPLR, D(13)=>
      OutputImg3_189_EXMPLR, D(12)=>OutputImg3_188_EXMPLR, D(11)=>
      OutputImg3_187_EXMPLR, D(10)=>OutputImg3_186_EXMPLR, D(9)=>
      OutputImg3_185_EXMPLR, D(8)=>OutputImg3_184_EXMPLR, D(7)=>
      OutputImg3_183_EXMPLR, D(6)=>OutputImg3_182_EXMPLR, D(5)=>
      OutputImg3_181_EXMPLR, D(4)=>OutputImg3_180_EXMPLR, D(3)=>
      OutputImg3_179_EXMPLR, D(2)=>OutputImg3_178_EXMPLR, D(1)=>
      OutputImg3_177_EXMPLR, D(0)=>OutputImg3_176_EXMPLR, EN=>nx23802, F(15)
      =>ImgReg2IN_191, F(14)=>ImgReg2IN_190, F(13)=>ImgReg2IN_189, F(12)=>
      ImgReg2IN_188, F(11)=>ImgReg2IN_187, F(10)=>ImgReg2IN_186, F(9)=>
      ImgReg2IN_185, F(8)=>ImgReg2IN_184, F(7)=>ImgReg2IN_183, F(6)=>
      ImgReg2IN_182, F(5)=>ImgReg2IN_181, F(4)=>ImgReg2IN_180, F(3)=>
      ImgReg2IN_179, F(2)=>ImgReg2IN_178, F(1)=>ImgReg2IN_177, F(0)=>
      ImgReg2IN_176);
   loop3_11_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_191_EXMPLR, D(14)=>OutputImg4_190_EXMPLR, D(13)=>
      OutputImg4_189_EXMPLR, D(12)=>OutputImg4_188_EXMPLR, D(11)=>
      OutputImg4_187_EXMPLR, D(10)=>OutputImg4_186_EXMPLR, D(9)=>
      OutputImg4_185_EXMPLR, D(8)=>OutputImg4_184_EXMPLR, D(7)=>
      OutputImg4_183_EXMPLR, D(6)=>OutputImg4_182_EXMPLR, D(5)=>
      OutputImg4_181_EXMPLR, D(4)=>OutputImg4_180_EXMPLR, D(3)=>
      OutputImg4_179_EXMPLR, D(2)=>OutputImg4_178_EXMPLR, D(1)=>
      OutputImg4_177_EXMPLR, D(0)=>OutputImg4_176_EXMPLR, EN=>nx23802, F(15)
      =>ImgReg3IN_191, F(14)=>ImgReg3IN_190, F(13)=>ImgReg3IN_189, F(12)=>
      ImgReg3IN_188, F(11)=>ImgReg3IN_187, F(10)=>ImgReg3IN_186, F(9)=>
      ImgReg3IN_185, F(8)=>ImgReg3IN_184, F(7)=>ImgReg3IN_183, F(6)=>
      ImgReg3IN_182, F(5)=>ImgReg3IN_181, F(4)=>ImgReg3IN_180, F(3)=>
      ImgReg3IN_179, F(2)=>ImgReg3IN_178, F(1)=>ImgReg3IN_177, F(0)=>
      ImgReg3IN_176);
   loop3_11_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_191_EXMPLR, D(14)=>OutputImg5_190_EXMPLR, D(13)=>
      OutputImg5_189_EXMPLR, D(12)=>OutputImg5_188_EXMPLR, D(11)=>
      OutputImg5_187_EXMPLR, D(10)=>OutputImg5_186_EXMPLR, D(9)=>
      OutputImg5_185_EXMPLR, D(8)=>OutputImg5_184_EXMPLR, D(7)=>
      OutputImg5_183_EXMPLR, D(6)=>OutputImg5_182_EXMPLR, D(5)=>
      OutputImg5_181_EXMPLR, D(4)=>OutputImg5_180_EXMPLR, D(3)=>
      OutputImg5_179_EXMPLR, D(2)=>OutputImg5_178_EXMPLR, D(1)=>
      OutputImg5_177_EXMPLR, D(0)=>OutputImg5_176_EXMPLR, EN=>nx23802, F(15)
      =>ImgReg4IN_191, F(14)=>ImgReg4IN_190, F(13)=>ImgReg4IN_189, F(12)=>
      ImgReg4IN_188, F(11)=>ImgReg4IN_187, F(10)=>ImgReg4IN_186, F(9)=>
      ImgReg4IN_185, F(8)=>ImgReg4IN_184, F(7)=>ImgReg4IN_183, F(6)=>
      ImgReg4IN_182, F(5)=>ImgReg4IN_181, F(4)=>ImgReg4IN_180, F(3)=>
      ImgReg4IN_179, F(2)=>ImgReg4IN_178, F(1)=>ImgReg4IN_177, F(0)=>
      ImgReg4IN_176);
   loop3_11_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_191, D(14)=>
      ImgReg0IN_190, D(13)=>ImgReg0IN_189, D(12)=>ImgReg0IN_188, D(11)=>
      ImgReg0IN_187, D(10)=>ImgReg0IN_186, D(9)=>ImgReg0IN_185, D(8)=>
      ImgReg0IN_184, D(7)=>ImgReg0IN_183, D(6)=>ImgReg0IN_182, D(5)=>
      ImgReg0IN_181, D(4)=>ImgReg0IN_180, D(3)=>ImgReg0IN_179, D(2)=>
      ImgReg0IN_178, D(1)=>ImgReg0IN_177, D(0)=>ImgReg0IN_176, CLK=>nx23894, 
      RST=>RST, EN=>nx23720, Q(15)=>OutputImg0_191_EXMPLR, Q(14)=>
      OutputImg0_190_EXMPLR, Q(13)=>OutputImg0_189_EXMPLR, Q(12)=>
      OutputImg0_188_EXMPLR, Q(11)=>OutputImg0_187_EXMPLR, Q(10)=>
      OutputImg0_186_EXMPLR, Q(9)=>OutputImg0_185_EXMPLR, Q(8)=>
      OutputImg0_184_EXMPLR, Q(7)=>OutputImg0_183_EXMPLR, Q(6)=>
      OutputImg0_182_EXMPLR, Q(5)=>OutputImg0_181_EXMPLR, Q(4)=>
      OutputImg0_180_EXMPLR, Q(3)=>OutputImg0_179_EXMPLR, Q(2)=>
      OutputImg0_178_EXMPLR, Q(1)=>OutputImg0_177_EXMPLR, Q(0)=>
      OutputImg0_176_EXMPLR);
   loop3_11_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_191, D(14)=>
      ImgReg1IN_190, D(13)=>ImgReg1IN_189, D(12)=>ImgReg1IN_188, D(11)=>
      ImgReg1IN_187, D(10)=>ImgReg1IN_186, D(9)=>ImgReg1IN_185, D(8)=>
      ImgReg1IN_184, D(7)=>ImgReg1IN_183, D(6)=>ImgReg1IN_182, D(5)=>
      ImgReg1IN_181, D(4)=>ImgReg1IN_180, D(3)=>ImgReg1IN_179, D(2)=>
      ImgReg1IN_178, D(1)=>ImgReg1IN_177, D(0)=>ImgReg1IN_176, CLK=>nx23896, 
      RST=>RST, EN=>nx23730, Q(15)=>OutputImg1_191_EXMPLR, Q(14)=>
      OutputImg1_190_EXMPLR, Q(13)=>OutputImg1_189_EXMPLR, Q(12)=>
      OutputImg1_188_EXMPLR, Q(11)=>OutputImg1_187_EXMPLR, Q(10)=>
      OutputImg1_186_EXMPLR, Q(9)=>OutputImg1_185_EXMPLR, Q(8)=>
      OutputImg1_184_EXMPLR, Q(7)=>OutputImg1_183_EXMPLR, Q(6)=>
      OutputImg1_182_EXMPLR, Q(5)=>OutputImg1_181_EXMPLR, Q(4)=>
      OutputImg1_180_EXMPLR, Q(3)=>OutputImg1_179_EXMPLR, Q(2)=>
      OutputImg1_178_EXMPLR, Q(1)=>OutputImg1_177_EXMPLR, Q(0)=>
      OutputImg1_176_EXMPLR);
   loop3_11_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_191, D(14)=>
      ImgReg2IN_190, D(13)=>ImgReg2IN_189, D(12)=>ImgReg2IN_188, D(11)=>
      ImgReg2IN_187, D(10)=>ImgReg2IN_186, D(9)=>ImgReg2IN_185, D(8)=>
      ImgReg2IN_184, D(7)=>ImgReg2IN_183, D(6)=>ImgReg2IN_182, D(5)=>
      ImgReg2IN_181, D(4)=>ImgReg2IN_180, D(3)=>ImgReg2IN_179, D(2)=>
      ImgReg2IN_178, D(1)=>ImgReg2IN_177, D(0)=>ImgReg2IN_176, CLK=>nx23896, 
      RST=>RST, EN=>nx23740, Q(15)=>OutputImg2_191_EXMPLR, Q(14)=>
      OutputImg2_190_EXMPLR, Q(13)=>OutputImg2_189_EXMPLR, Q(12)=>
      OutputImg2_188_EXMPLR, Q(11)=>OutputImg2_187_EXMPLR, Q(10)=>
      OutputImg2_186_EXMPLR, Q(9)=>OutputImg2_185_EXMPLR, Q(8)=>
      OutputImg2_184_EXMPLR, Q(7)=>OutputImg2_183_EXMPLR, Q(6)=>
      OutputImg2_182_EXMPLR, Q(5)=>OutputImg2_181_EXMPLR, Q(4)=>
      OutputImg2_180_EXMPLR, Q(3)=>OutputImg2_179_EXMPLR, Q(2)=>
      OutputImg2_178_EXMPLR, Q(1)=>OutputImg2_177_EXMPLR, Q(0)=>
      OutputImg2_176_EXMPLR);
   loop3_11_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_191, D(14)=>
      ImgReg3IN_190, D(13)=>ImgReg3IN_189, D(12)=>ImgReg3IN_188, D(11)=>
      ImgReg3IN_187, D(10)=>ImgReg3IN_186, D(9)=>ImgReg3IN_185, D(8)=>
      ImgReg3IN_184, D(7)=>ImgReg3IN_183, D(6)=>ImgReg3IN_182, D(5)=>
      ImgReg3IN_181, D(4)=>ImgReg3IN_180, D(3)=>ImgReg3IN_179, D(2)=>
      ImgReg3IN_178, D(1)=>ImgReg3IN_177, D(0)=>ImgReg3IN_176, CLK=>nx23898, 
      RST=>RST, EN=>nx23750, Q(15)=>OutputImg3_191_EXMPLR, Q(14)=>
      OutputImg3_190_EXMPLR, Q(13)=>OutputImg3_189_EXMPLR, Q(12)=>
      OutputImg3_188_EXMPLR, Q(11)=>OutputImg3_187_EXMPLR, Q(10)=>
      OutputImg3_186_EXMPLR, Q(9)=>OutputImg3_185_EXMPLR, Q(8)=>
      OutputImg3_184_EXMPLR, Q(7)=>OutputImg3_183_EXMPLR, Q(6)=>
      OutputImg3_182_EXMPLR, Q(5)=>OutputImg3_181_EXMPLR, Q(4)=>
      OutputImg3_180_EXMPLR, Q(3)=>OutputImg3_179_EXMPLR, Q(2)=>
      OutputImg3_178_EXMPLR, Q(1)=>OutputImg3_177_EXMPLR, Q(0)=>
      OutputImg3_176_EXMPLR);
   loop3_11_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_191, D(14)=>
      ImgReg4IN_190, D(13)=>ImgReg4IN_189, D(12)=>ImgReg4IN_188, D(11)=>
      ImgReg4IN_187, D(10)=>ImgReg4IN_186, D(9)=>ImgReg4IN_185, D(8)=>
      ImgReg4IN_184, D(7)=>ImgReg4IN_183, D(6)=>ImgReg4IN_182, D(5)=>
      ImgReg4IN_181, D(4)=>ImgReg4IN_180, D(3)=>ImgReg4IN_179, D(2)=>
      ImgReg4IN_178, D(1)=>ImgReg4IN_177, D(0)=>ImgReg4IN_176, CLK=>nx23898, 
      RST=>RST, EN=>nx23760, Q(15)=>OutputImg4_191_EXMPLR, Q(14)=>
      OutputImg4_190_EXMPLR, Q(13)=>OutputImg4_189_EXMPLR, Q(12)=>
      OutputImg4_188_EXMPLR, Q(11)=>OutputImg4_187_EXMPLR, Q(10)=>
      OutputImg4_186_EXMPLR, Q(9)=>OutputImg4_185_EXMPLR, Q(8)=>
      OutputImg4_184_EXMPLR, Q(7)=>OutputImg4_183_EXMPLR, Q(6)=>
      OutputImg4_182_EXMPLR, Q(5)=>OutputImg4_181_EXMPLR, Q(4)=>
      OutputImg4_180_EXMPLR, Q(3)=>OutputImg4_179_EXMPLR, Q(2)=>
      OutputImg4_178_EXMPLR, Q(1)=>OutputImg4_177_EXMPLR, Q(0)=>
      OutputImg4_176_EXMPLR);
   loop3_11_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_191, D(14)=>
      ImgReg5IN_190, D(13)=>ImgReg5IN_189, D(12)=>ImgReg5IN_188, D(11)=>
      ImgReg5IN_187, D(10)=>ImgReg5IN_186, D(9)=>ImgReg5IN_185, D(8)=>
      ImgReg5IN_184, D(7)=>ImgReg5IN_183, D(6)=>ImgReg5IN_182, D(5)=>
      ImgReg5IN_181, D(4)=>ImgReg5IN_180, D(3)=>ImgReg5IN_179, D(2)=>
      ImgReg5IN_178, D(1)=>ImgReg5IN_177, D(0)=>ImgReg5IN_176, CLK=>nx23900, 
      RST=>RST, EN=>nx23770, Q(15)=>OutputImg5_191_EXMPLR, Q(14)=>
      OutputImg5_190_EXMPLR, Q(13)=>OutputImg5_189_EXMPLR, Q(12)=>
      OutputImg5_188_EXMPLR, Q(11)=>OutputImg5_187_EXMPLR, Q(10)=>
      OutputImg5_186_EXMPLR, Q(9)=>OutputImg5_185_EXMPLR, Q(8)=>
      OutputImg5_184_EXMPLR, Q(7)=>OutputImg5_183_EXMPLR, Q(6)=>
      OutputImg5_182_EXMPLR, Q(5)=>OutputImg5_181_EXMPLR, Q(4)=>
      OutputImg5_180_EXMPLR, Q(3)=>OutputImg5_179_EXMPLR, Q(2)=>
      OutputImg5_178_EXMPLR, Q(1)=>OutputImg5_177_EXMPLR, Q(0)=>
      OutputImg5_176_EXMPLR);
   loop3_12_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_223_EXMPLR, D(14)=>OutputImg0_222_EXMPLR, D(13)=>
      OutputImg0_221_EXMPLR, D(12)=>OutputImg0_220_EXMPLR, D(11)=>
      OutputImg0_219_EXMPLR, D(10)=>OutputImg0_218_EXMPLR, D(9)=>
      OutputImg0_217_EXMPLR, D(8)=>OutputImg0_216_EXMPLR, D(7)=>
      OutputImg0_215_EXMPLR, D(6)=>OutputImg0_214_EXMPLR, D(5)=>
      OutputImg0_213_EXMPLR, D(4)=>OutputImg0_212_EXMPLR, D(3)=>
      OutputImg0_211_EXMPLR, D(2)=>OutputImg0_210_EXMPLR, D(1)=>
      OutputImg0_209_EXMPLR, D(0)=>OutputImg0_208_EXMPLR, EN=>nx23686, F(15)
      =>ImgReg0IN_207, F(14)=>ImgReg0IN_206, F(13)=>ImgReg0IN_205, F(12)=>
      ImgReg0IN_204, F(11)=>ImgReg0IN_203, F(10)=>ImgReg0IN_202, F(9)=>
      ImgReg0IN_201, F(8)=>ImgReg0IN_200, F(7)=>ImgReg0IN_199, F(6)=>
      ImgReg0IN_198, F(5)=>ImgReg0IN_197, F(4)=>ImgReg0IN_196, F(3)=>
      ImgReg0IN_195, F(2)=>ImgReg0IN_194, F(1)=>ImgReg0IN_193, F(0)=>
      ImgReg0IN_192);
   loop3_12_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_223_EXMPLR, D(14)=>OutputImg1_222_EXMPLR, D(13)=>
      OutputImg1_221_EXMPLR, D(12)=>OutputImg1_220_EXMPLR, D(11)=>
      OutputImg1_219_EXMPLR, D(10)=>OutputImg1_218_EXMPLR, D(9)=>
      OutputImg1_217_EXMPLR, D(8)=>OutputImg1_216_EXMPLR, D(7)=>
      OutputImg1_215_EXMPLR, D(6)=>OutputImg1_214_EXMPLR, D(5)=>
      OutputImg1_213_EXMPLR, D(4)=>OutputImg1_212_EXMPLR, D(3)=>
      OutputImg1_211_EXMPLR, D(2)=>OutputImg1_210_EXMPLR, D(1)=>
      OutputImg1_209_EXMPLR, D(0)=>OutputImg1_208_EXMPLR, EN=>nx23686, F(15)
      =>ImgReg1IN_207, F(14)=>ImgReg1IN_206, F(13)=>ImgReg1IN_205, F(12)=>
      ImgReg1IN_204, F(11)=>ImgReg1IN_203, F(10)=>ImgReg1IN_202, F(9)=>
      ImgReg1IN_201, F(8)=>ImgReg1IN_200, F(7)=>ImgReg1IN_199, F(6)=>
      ImgReg1IN_198, F(5)=>ImgReg1IN_197, F(4)=>ImgReg1IN_196, F(3)=>
      ImgReg1IN_195, F(2)=>ImgReg1IN_194, F(1)=>ImgReg1IN_193, F(0)=>
      ImgReg1IN_192);
   loop3_12_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_223_EXMPLR, D(14)=>OutputImg2_222_EXMPLR, D(13)=>
      OutputImg2_221_EXMPLR, D(12)=>OutputImg2_220_EXMPLR, D(11)=>
      OutputImg2_219_EXMPLR, D(10)=>OutputImg2_218_EXMPLR, D(9)=>
      OutputImg2_217_EXMPLR, D(8)=>OutputImg2_216_EXMPLR, D(7)=>
      OutputImg2_215_EXMPLR, D(6)=>OutputImg2_214_EXMPLR, D(5)=>
      OutputImg2_213_EXMPLR, D(4)=>OutputImg2_212_EXMPLR, D(3)=>
      OutputImg2_211_EXMPLR, D(2)=>OutputImg2_210_EXMPLR, D(1)=>
      OutputImg2_209_EXMPLR, D(0)=>OutputImg2_208_EXMPLR, EN=>nx23686, F(15)
      =>ImgReg2IN_207, F(14)=>ImgReg2IN_206, F(13)=>ImgReg2IN_205, F(12)=>
      ImgReg2IN_204, F(11)=>ImgReg2IN_203, F(10)=>ImgReg2IN_202, F(9)=>
      ImgReg2IN_201, F(8)=>ImgReg2IN_200, F(7)=>ImgReg2IN_199, F(6)=>
      ImgReg2IN_198, F(5)=>ImgReg2IN_197, F(4)=>ImgReg2IN_196, F(3)=>
      ImgReg2IN_195, F(2)=>ImgReg2IN_194, F(1)=>ImgReg2IN_193, F(0)=>
      ImgReg2IN_192);
   loop3_12_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_223_EXMPLR, D(14)=>OutputImg3_222_EXMPLR, D(13)=>
      OutputImg3_221_EXMPLR, D(12)=>OutputImg3_220_EXMPLR, D(11)=>
      OutputImg3_219_EXMPLR, D(10)=>OutputImg3_218_EXMPLR, D(9)=>
      OutputImg3_217_EXMPLR, D(8)=>OutputImg3_216_EXMPLR, D(7)=>
      OutputImg3_215_EXMPLR, D(6)=>OutputImg3_214_EXMPLR, D(5)=>
      OutputImg3_213_EXMPLR, D(4)=>OutputImg3_212_EXMPLR, D(3)=>
      OutputImg3_211_EXMPLR, D(2)=>OutputImg3_210_EXMPLR, D(1)=>
      OutputImg3_209_EXMPLR, D(0)=>OutputImg3_208_EXMPLR, EN=>nx23686, F(15)
      =>ImgReg3IN_207, F(14)=>ImgReg3IN_206, F(13)=>ImgReg3IN_205, F(12)=>
      ImgReg3IN_204, F(11)=>ImgReg3IN_203, F(10)=>ImgReg3IN_202, F(9)=>
      ImgReg3IN_201, F(8)=>ImgReg3IN_200, F(7)=>ImgReg3IN_199, F(6)=>
      ImgReg3IN_198, F(5)=>ImgReg3IN_197, F(4)=>ImgReg3IN_196, F(3)=>
      ImgReg3IN_195, F(2)=>ImgReg3IN_194, F(1)=>ImgReg3IN_193, F(0)=>
      ImgReg3IN_192);
   loop3_12_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_223_EXMPLR, D(14)=>OutputImg4_222_EXMPLR, D(13)=>
      OutputImg4_221_EXMPLR, D(12)=>OutputImg4_220_EXMPLR, D(11)=>
      OutputImg4_219_EXMPLR, D(10)=>OutputImg4_218_EXMPLR, D(9)=>
      OutputImg4_217_EXMPLR, D(8)=>OutputImg4_216_EXMPLR, D(7)=>
      OutputImg4_215_EXMPLR, D(6)=>OutputImg4_214_EXMPLR, D(5)=>
      OutputImg4_213_EXMPLR, D(4)=>OutputImg4_212_EXMPLR, D(3)=>
      OutputImg4_211_EXMPLR, D(2)=>OutputImg4_210_EXMPLR, D(1)=>
      OutputImg4_209_EXMPLR, D(0)=>OutputImg4_208_EXMPLR, EN=>nx23686, F(15)
      =>ImgReg4IN_207, F(14)=>ImgReg4IN_206, F(13)=>ImgReg4IN_205, F(12)=>
      ImgReg4IN_204, F(11)=>ImgReg4IN_203, F(10)=>ImgReg4IN_202, F(9)=>
      ImgReg4IN_201, F(8)=>ImgReg4IN_200, F(7)=>ImgReg4IN_199, F(6)=>
      ImgReg4IN_198, F(5)=>ImgReg4IN_197, F(4)=>ImgReg4IN_196, F(3)=>
      ImgReg4IN_195, F(2)=>ImgReg4IN_194, F(1)=>ImgReg4IN_193, F(0)=>
      ImgReg4IN_192);
   loop3_12_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_223_EXMPLR, D(14)=>OutputImg5_222_EXMPLR, D(13)=>
      OutputImg5_221_EXMPLR, D(12)=>OutputImg5_220_EXMPLR, D(11)=>
      OutputImg5_219_EXMPLR, D(10)=>OutputImg5_218_EXMPLR, D(9)=>
      OutputImg5_217_EXMPLR, D(8)=>OutputImg5_216_EXMPLR, D(7)=>
      OutputImg5_215_EXMPLR, D(6)=>OutputImg5_214_EXMPLR, D(5)=>
      OutputImg5_213_EXMPLR, D(4)=>OutputImg5_212_EXMPLR, D(3)=>
      OutputImg5_211_EXMPLR, D(2)=>OutputImg5_210_EXMPLR, D(1)=>
      OutputImg5_209_EXMPLR, D(0)=>OutputImg5_208_EXMPLR, EN=>nx23688, F(15)
      =>ImgReg5IN_207, F(14)=>ImgReg5IN_206, F(13)=>ImgReg5IN_205, F(12)=>
      ImgReg5IN_204, F(11)=>ImgReg5IN_203, F(10)=>ImgReg5IN_202, F(9)=>
      ImgReg5IN_201, F(8)=>ImgReg5IN_200, F(7)=>ImgReg5IN_199, F(6)=>
      ImgReg5IN_198, F(5)=>ImgReg5IN_197, F(4)=>ImgReg5IN_196, F(3)=>
      ImgReg5IN_195, F(2)=>ImgReg5IN_194, F(1)=>ImgReg5IN_193, F(0)=>
      ImgReg5IN_192);
   loop3_12_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(207), 
      D(14)=>DATA(206), D(13)=>DATA(205), D(12)=>DATA(204), D(11)=>DATA(203), 
      D(10)=>DATA(202), D(9)=>DATA(201), D(8)=>DATA(200), D(7)=>DATA(199), 
      D(6)=>DATA(198), D(5)=>DATA(197), D(4)=>DATA(196), D(3)=>DATA(195), 
      D(2)=>DATA(194), D(1)=>DATA(193), D(0)=>DATA(192), EN=>nx23656, F(15)
      =>ImgReg0IN_207, F(14)=>ImgReg0IN_206, F(13)=>ImgReg0IN_205, F(12)=>
      ImgReg0IN_204, F(11)=>ImgReg0IN_203, F(10)=>ImgReg0IN_202, F(9)=>
      ImgReg0IN_201, F(8)=>ImgReg0IN_200, F(7)=>ImgReg0IN_199, F(6)=>
      ImgReg0IN_198, F(5)=>ImgReg0IN_197, F(4)=>ImgReg0IN_196, F(3)=>
      ImgReg0IN_195, F(2)=>ImgReg0IN_194, F(1)=>ImgReg0IN_193, F(0)=>
      ImgReg0IN_192);
   loop3_12_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(207), 
      D(14)=>DATA(206), D(13)=>DATA(205), D(12)=>DATA(204), D(11)=>DATA(203), 
      D(10)=>DATA(202), D(9)=>DATA(201), D(8)=>DATA(200), D(7)=>DATA(199), 
      D(6)=>DATA(198), D(5)=>DATA(197), D(4)=>DATA(196), D(3)=>DATA(195), 
      D(2)=>DATA(194), D(1)=>DATA(193), D(0)=>DATA(192), EN=>nx23644, F(15)
      =>ImgReg1IN_207, F(14)=>ImgReg1IN_206, F(13)=>ImgReg1IN_205, F(12)=>
      ImgReg1IN_204, F(11)=>ImgReg1IN_203, F(10)=>ImgReg1IN_202, F(9)=>
      ImgReg1IN_201, F(8)=>ImgReg1IN_200, F(7)=>ImgReg1IN_199, F(6)=>
      ImgReg1IN_198, F(5)=>ImgReg1IN_197, F(4)=>ImgReg1IN_196, F(3)=>
      ImgReg1IN_195, F(2)=>ImgReg1IN_194, F(1)=>ImgReg1IN_193, F(0)=>
      ImgReg1IN_192);
   loop3_12_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(207), 
      D(14)=>DATA(206), D(13)=>DATA(205), D(12)=>DATA(204), D(11)=>DATA(203), 
      D(10)=>DATA(202), D(9)=>DATA(201), D(8)=>DATA(200), D(7)=>DATA(199), 
      D(6)=>DATA(198), D(5)=>DATA(197), D(4)=>DATA(196), D(3)=>DATA(195), 
      D(2)=>DATA(194), D(1)=>DATA(193), D(0)=>DATA(192), EN=>nx23632, F(15)
      =>ImgReg2IN_207, F(14)=>ImgReg2IN_206, F(13)=>ImgReg2IN_205, F(12)=>
      ImgReg2IN_204, F(11)=>ImgReg2IN_203, F(10)=>ImgReg2IN_202, F(9)=>
      ImgReg2IN_201, F(8)=>ImgReg2IN_200, F(7)=>ImgReg2IN_199, F(6)=>
      ImgReg2IN_198, F(5)=>ImgReg2IN_197, F(4)=>ImgReg2IN_196, F(3)=>
      ImgReg2IN_195, F(2)=>ImgReg2IN_194, F(1)=>ImgReg2IN_193, F(0)=>
      ImgReg2IN_192);
   loop3_12_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(207), 
      D(14)=>DATA(206), D(13)=>DATA(205), D(12)=>DATA(204), D(11)=>DATA(203), 
      D(10)=>DATA(202), D(9)=>DATA(201), D(8)=>DATA(200), D(7)=>DATA(199), 
      D(6)=>DATA(198), D(5)=>DATA(197), D(4)=>DATA(196), D(3)=>DATA(195), 
      D(2)=>DATA(194), D(1)=>DATA(193), D(0)=>DATA(192), EN=>nx23620, F(15)
      =>ImgReg3IN_207, F(14)=>ImgReg3IN_206, F(13)=>ImgReg3IN_205, F(12)=>
      ImgReg3IN_204, F(11)=>ImgReg3IN_203, F(10)=>ImgReg3IN_202, F(9)=>
      ImgReg3IN_201, F(8)=>ImgReg3IN_200, F(7)=>ImgReg3IN_199, F(6)=>
      ImgReg3IN_198, F(5)=>ImgReg3IN_197, F(4)=>ImgReg3IN_196, F(3)=>
      ImgReg3IN_195, F(2)=>ImgReg3IN_194, F(1)=>ImgReg3IN_193, F(0)=>
      ImgReg3IN_192);
   loop3_12_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(207), 
      D(14)=>DATA(206), D(13)=>DATA(205), D(12)=>DATA(204), D(11)=>DATA(203), 
      D(10)=>DATA(202), D(9)=>DATA(201), D(8)=>DATA(200), D(7)=>DATA(199), 
      D(6)=>DATA(198), D(5)=>DATA(197), D(4)=>DATA(196), D(3)=>DATA(195), 
      D(2)=>DATA(194), D(1)=>DATA(193), D(0)=>DATA(192), EN=>nx23608, F(15)
      =>ImgReg4IN_207, F(14)=>ImgReg4IN_206, F(13)=>ImgReg4IN_205, F(12)=>
      ImgReg4IN_204, F(11)=>ImgReg4IN_203, F(10)=>ImgReg4IN_202, F(9)=>
      ImgReg4IN_201, F(8)=>ImgReg4IN_200, F(7)=>ImgReg4IN_199, F(6)=>
      ImgReg4IN_198, F(5)=>ImgReg4IN_197, F(4)=>ImgReg4IN_196, F(3)=>
      ImgReg4IN_195, F(2)=>ImgReg4IN_194, F(1)=>ImgReg4IN_193, F(0)=>
      ImgReg4IN_192);
   loop3_12_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(207), 
      D(14)=>DATA(206), D(13)=>DATA(205), D(12)=>DATA(204), D(11)=>DATA(203), 
      D(10)=>DATA(202), D(9)=>DATA(201), D(8)=>DATA(200), D(7)=>DATA(199), 
      D(6)=>DATA(198), D(5)=>DATA(197), D(4)=>DATA(196), D(3)=>DATA(195), 
      D(2)=>DATA(194), D(1)=>DATA(193), D(0)=>DATA(192), EN=>nx23596, F(15)
      =>ImgReg5IN_207, F(14)=>ImgReg5IN_206, F(13)=>ImgReg5IN_205, F(12)=>
      ImgReg5IN_204, F(11)=>ImgReg5IN_203, F(10)=>ImgReg5IN_202, F(9)=>
      ImgReg5IN_201, F(8)=>ImgReg5IN_200, F(7)=>ImgReg5IN_199, F(6)=>
      ImgReg5IN_198, F(5)=>ImgReg5IN_197, F(4)=>ImgReg5IN_196, F(3)=>
      ImgReg5IN_195, F(2)=>ImgReg5IN_194, F(1)=>ImgReg5IN_193, F(0)=>
      ImgReg5IN_192);
   loop3_12_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_207_EXMPLR, D(14)=>OutputImg1_206_EXMPLR, D(13)=>
      OutputImg1_205_EXMPLR, D(12)=>OutputImg1_204_EXMPLR, D(11)=>
      OutputImg1_203_EXMPLR, D(10)=>OutputImg1_202_EXMPLR, D(9)=>
      OutputImg1_201_EXMPLR, D(8)=>OutputImg1_200_EXMPLR, D(7)=>
      OutputImg1_199_EXMPLR, D(6)=>OutputImg1_198_EXMPLR, D(5)=>
      OutputImg1_197_EXMPLR, D(4)=>OutputImg1_196_EXMPLR, D(3)=>
      OutputImg1_195_EXMPLR, D(2)=>OutputImg1_194_EXMPLR, D(1)=>
      OutputImg1_193_EXMPLR, D(0)=>OutputImg1_192_EXMPLR, EN=>nx23802, F(15)
      =>ImgReg0IN_207, F(14)=>ImgReg0IN_206, F(13)=>ImgReg0IN_205, F(12)=>
      ImgReg0IN_204, F(11)=>ImgReg0IN_203, F(10)=>ImgReg0IN_202, F(9)=>
      ImgReg0IN_201, F(8)=>ImgReg0IN_200, F(7)=>ImgReg0IN_199, F(6)=>
      ImgReg0IN_198, F(5)=>ImgReg0IN_197, F(4)=>ImgReg0IN_196, F(3)=>
      ImgReg0IN_195, F(2)=>ImgReg0IN_194, F(1)=>ImgReg0IN_193, F(0)=>
      ImgReg0IN_192);
   loop3_12_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_207_EXMPLR, D(14)=>OutputImg2_206_EXMPLR, D(13)=>
      OutputImg2_205_EXMPLR, D(12)=>OutputImg2_204_EXMPLR, D(11)=>
      OutputImg2_203_EXMPLR, D(10)=>OutputImg2_202_EXMPLR, D(9)=>
      OutputImg2_201_EXMPLR, D(8)=>OutputImg2_200_EXMPLR, D(7)=>
      OutputImg2_199_EXMPLR, D(6)=>OutputImg2_198_EXMPLR, D(5)=>
      OutputImg2_197_EXMPLR, D(4)=>OutputImg2_196_EXMPLR, D(3)=>
      OutputImg2_195_EXMPLR, D(2)=>OutputImg2_194_EXMPLR, D(1)=>
      OutputImg2_193_EXMPLR, D(0)=>OutputImg2_192_EXMPLR, EN=>nx23802, F(15)
      =>ImgReg1IN_207, F(14)=>ImgReg1IN_206, F(13)=>ImgReg1IN_205, F(12)=>
      ImgReg1IN_204, F(11)=>ImgReg1IN_203, F(10)=>ImgReg1IN_202, F(9)=>
      ImgReg1IN_201, F(8)=>ImgReg1IN_200, F(7)=>ImgReg1IN_199, F(6)=>
      ImgReg1IN_198, F(5)=>ImgReg1IN_197, F(4)=>ImgReg1IN_196, F(3)=>
      ImgReg1IN_195, F(2)=>ImgReg1IN_194, F(1)=>ImgReg1IN_193, F(0)=>
      ImgReg1IN_192);
   loop3_12_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_207_EXMPLR, D(14)=>OutputImg3_206_EXMPLR, D(13)=>
      OutputImg3_205_EXMPLR, D(12)=>OutputImg3_204_EXMPLR, D(11)=>
      OutputImg3_203_EXMPLR, D(10)=>OutputImg3_202_EXMPLR, D(9)=>
      OutputImg3_201_EXMPLR, D(8)=>OutputImg3_200_EXMPLR, D(7)=>
      OutputImg3_199_EXMPLR, D(6)=>OutputImg3_198_EXMPLR, D(5)=>
      OutputImg3_197_EXMPLR, D(4)=>OutputImg3_196_EXMPLR, D(3)=>
      OutputImg3_195_EXMPLR, D(2)=>OutputImg3_194_EXMPLR, D(1)=>
      OutputImg3_193_EXMPLR, D(0)=>OutputImg3_192_EXMPLR, EN=>nx23802, F(15)
      =>ImgReg2IN_207, F(14)=>ImgReg2IN_206, F(13)=>ImgReg2IN_205, F(12)=>
      ImgReg2IN_204, F(11)=>ImgReg2IN_203, F(10)=>ImgReg2IN_202, F(9)=>
      ImgReg2IN_201, F(8)=>ImgReg2IN_200, F(7)=>ImgReg2IN_199, F(6)=>
      ImgReg2IN_198, F(5)=>ImgReg2IN_197, F(4)=>ImgReg2IN_196, F(3)=>
      ImgReg2IN_195, F(2)=>ImgReg2IN_194, F(1)=>ImgReg2IN_193, F(0)=>
      ImgReg2IN_192);
   loop3_12_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_207_EXMPLR, D(14)=>OutputImg4_206_EXMPLR, D(13)=>
      OutputImg4_205_EXMPLR, D(12)=>OutputImg4_204_EXMPLR, D(11)=>
      OutputImg4_203_EXMPLR, D(10)=>OutputImg4_202_EXMPLR, D(9)=>
      OutputImg4_201_EXMPLR, D(8)=>OutputImg4_200_EXMPLR, D(7)=>
      OutputImg4_199_EXMPLR, D(6)=>OutputImg4_198_EXMPLR, D(5)=>
      OutputImg4_197_EXMPLR, D(4)=>OutputImg4_196_EXMPLR, D(3)=>
      OutputImg4_195_EXMPLR, D(2)=>OutputImg4_194_EXMPLR, D(1)=>
      OutputImg4_193_EXMPLR, D(0)=>OutputImg4_192_EXMPLR, EN=>nx23804, F(15)
      =>ImgReg3IN_207, F(14)=>ImgReg3IN_206, F(13)=>ImgReg3IN_205, F(12)=>
      ImgReg3IN_204, F(11)=>ImgReg3IN_203, F(10)=>ImgReg3IN_202, F(9)=>
      ImgReg3IN_201, F(8)=>ImgReg3IN_200, F(7)=>ImgReg3IN_199, F(6)=>
      ImgReg3IN_198, F(5)=>ImgReg3IN_197, F(4)=>ImgReg3IN_196, F(3)=>
      ImgReg3IN_195, F(2)=>ImgReg3IN_194, F(1)=>ImgReg3IN_193, F(0)=>
      ImgReg3IN_192);
   loop3_12_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_207_EXMPLR, D(14)=>OutputImg5_206_EXMPLR, D(13)=>
      OutputImg5_205_EXMPLR, D(12)=>OutputImg5_204_EXMPLR, D(11)=>
      OutputImg5_203_EXMPLR, D(10)=>OutputImg5_202_EXMPLR, D(9)=>
      OutputImg5_201_EXMPLR, D(8)=>OutputImg5_200_EXMPLR, D(7)=>
      OutputImg5_199_EXMPLR, D(6)=>OutputImg5_198_EXMPLR, D(5)=>
      OutputImg5_197_EXMPLR, D(4)=>OutputImg5_196_EXMPLR, D(3)=>
      OutputImg5_195_EXMPLR, D(2)=>OutputImg5_194_EXMPLR, D(1)=>
      OutputImg5_193_EXMPLR, D(0)=>OutputImg5_192_EXMPLR, EN=>nx23804, F(15)
      =>ImgReg4IN_207, F(14)=>ImgReg4IN_206, F(13)=>ImgReg4IN_205, F(12)=>
      ImgReg4IN_204, F(11)=>ImgReg4IN_203, F(10)=>ImgReg4IN_202, F(9)=>
      ImgReg4IN_201, F(8)=>ImgReg4IN_200, F(7)=>ImgReg4IN_199, F(6)=>
      ImgReg4IN_198, F(5)=>ImgReg4IN_197, F(4)=>ImgReg4IN_196, F(3)=>
      ImgReg4IN_195, F(2)=>ImgReg4IN_194, F(1)=>ImgReg4IN_193, F(0)=>
      ImgReg4IN_192);
   loop3_12_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_207, D(14)=>
      ImgReg0IN_206, D(13)=>ImgReg0IN_205, D(12)=>ImgReg0IN_204, D(11)=>
      ImgReg0IN_203, D(10)=>ImgReg0IN_202, D(9)=>ImgReg0IN_201, D(8)=>
      ImgReg0IN_200, D(7)=>ImgReg0IN_199, D(6)=>ImgReg0IN_198, D(5)=>
      ImgReg0IN_197, D(4)=>ImgReg0IN_196, D(3)=>ImgReg0IN_195, D(2)=>
      ImgReg0IN_194, D(1)=>ImgReg0IN_193, D(0)=>ImgReg0IN_192, CLK=>nx23900, 
      RST=>RST, EN=>nx23720, Q(15)=>OutputImg0_207_EXMPLR, Q(14)=>
      OutputImg0_206_EXMPLR, Q(13)=>OutputImg0_205_EXMPLR, Q(12)=>
      OutputImg0_204_EXMPLR, Q(11)=>OutputImg0_203_EXMPLR, Q(10)=>
      OutputImg0_202_EXMPLR, Q(9)=>OutputImg0_201_EXMPLR, Q(8)=>
      OutputImg0_200_EXMPLR, Q(7)=>OutputImg0_199_EXMPLR, Q(6)=>
      OutputImg0_198_EXMPLR, Q(5)=>OutputImg0_197_EXMPLR, Q(4)=>
      OutputImg0_196_EXMPLR, Q(3)=>OutputImg0_195_EXMPLR, Q(2)=>
      OutputImg0_194_EXMPLR, Q(1)=>OutputImg0_193_EXMPLR, Q(0)=>
      OutputImg0_192_EXMPLR);
   loop3_12_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_207, D(14)=>
      ImgReg1IN_206, D(13)=>ImgReg1IN_205, D(12)=>ImgReg1IN_204, D(11)=>
      ImgReg1IN_203, D(10)=>ImgReg1IN_202, D(9)=>ImgReg1IN_201, D(8)=>
      ImgReg1IN_200, D(7)=>ImgReg1IN_199, D(6)=>ImgReg1IN_198, D(5)=>
      ImgReg1IN_197, D(4)=>ImgReg1IN_196, D(3)=>ImgReg1IN_195, D(2)=>
      ImgReg1IN_194, D(1)=>ImgReg1IN_193, D(0)=>ImgReg1IN_192, CLK=>nx23902, 
      RST=>RST, EN=>nx23730, Q(15)=>OutputImg1_207_EXMPLR, Q(14)=>
      OutputImg1_206_EXMPLR, Q(13)=>OutputImg1_205_EXMPLR, Q(12)=>
      OutputImg1_204_EXMPLR, Q(11)=>OutputImg1_203_EXMPLR, Q(10)=>
      OutputImg1_202_EXMPLR, Q(9)=>OutputImg1_201_EXMPLR, Q(8)=>
      OutputImg1_200_EXMPLR, Q(7)=>OutputImg1_199_EXMPLR, Q(6)=>
      OutputImg1_198_EXMPLR, Q(5)=>OutputImg1_197_EXMPLR, Q(4)=>
      OutputImg1_196_EXMPLR, Q(3)=>OutputImg1_195_EXMPLR, Q(2)=>
      OutputImg1_194_EXMPLR, Q(1)=>OutputImg1_193_EXMPLR, Q(0)=>
      OutputImg1_192_EXMPLR);
   loop3_12_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_207, D(14)=>
      ImgReg2IN_206, D(13)=>ImgReg2IN_205, D(12)=>ImgReg2IN_204, D(11)=>
      ImgReg2IN_203, D(10)=>ImgReg2IN_202, D(9)=>ImgReg2IN_201, D(8)=>
      ImgReg2IN_200, D(7)=>ImgReg2IN_199, D(6)=>ImgReg2IN_198, D(5)=>
      ImgReg2IN_197, D(4)=>ImgReg2IN_196, D(3)=>ImgReg2IN_195, D(2)=>
      ImgReg2IN_194, D(1)=>ImgReg2IN_193, D(0)=>ImgReg2IN_192, CLK=>nx23902, 
      RST=>RST, EN=>nx23740, Q(15)=>OutputImg2_207_EXMPLR, Q(14)=>
      OutputImg2_206_EXMPLR, Q(13)=>OutputImg2_205_EXMPLR, Q(12)=>
      OutputImg2_204_EXMPLR, Q(11)=>OutputImg2_203_EXMPLR, Q(10)=>
      OutputImg2_202_EXMPLR, Q(9)=>OutputImg2_201_EXMPLR, Q(8)=>
      OutputImg2_200_EXMPLR, Q(7)=>OutputImg2_199_EXMPLR, Q(6)=>
      OutputImg2_198_EXMPLR, Q(5)=>OutputImg2_197_EXMPLR, Q(4)=>
      OutputImg2_196_EXMPLR, Q(3)=>OutputImg2_195_EXMPLR, Q(2)=>
      OutputImg2_194_EXMPLR, Q(1)=>OutputImg2_193_EXMPLR, Q(0)=>
      OutputImg2_192_EXMPLR);
   loop3_12_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_207, D(14)=>
      ImgReg3IN_206, D(13)=>ImgReg3IN_205, D(12)=>ImgReg3IN_204, D(11)=>
      ImgReg3IN_203, D(10)=>ImgReg3IN_202, D(9)=>ImgReg3IN_201, D(8)=>
      ImgReg3IN_200, D(7)=>ImgReg3IN_199, D(6)=>ImgReg3IN_198, D(5)=>
      ImgReg3IN_197, D(4)=>ImgReg3IN_196, D(3)=>ImgReg3IN_195, D(2)=>
      ImgReg3IN_194, D(1)=>ImgReg3IN_193, D(0)=>ImgReg3IN_192, CLK=>nx23904, 
      RST=>RST, EN=>nx23750, Q(15)=>OutputImg3_207_EXMPLR, Q(14)=>
      OutputImg3_206_EXMPLR, Q(13)=>OutputImg3_205_EXMPLR, Q(12)=>
      OutputImg3_204_EXMPLR, Q(11)=>OutputImg3_203_EXMPLR, Q(10)=>
      OutputImg3_202_EXMPLR, Q(9)=>OutputImg3_201_EXMPLR, Q(8)=>
      OutputImg3_200_EXMPLR, Q(7)=>OutputImg3_199_EXMPLR, Q(6)=>
      OutputImg3_198_EXMPLR, Q(5)=>OutputImg3_197_EXMPLR, Q(4)=>
      OutputImg3_196_EXMPLR, Q(3)=>OutputImg3_195_EXMPLR, Q(2)=>
      OutputImg3_194_EXMPLR, Q(1)=>OutputImg3_193_EXMPLR, Q(0)=>
      OutputImg3_192_EXMPLR);
   loop3_12_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_207, D(14)=>
      ImgReg4IN_206, D(13)=>ImgReg4IN_205, D(12)=>ImgReg4IN_204, D(11)=>
      ImgReg4IN_203, D(10)=>ImgReg4IN_202, D(9)=>ImgReg4IN_201, D(8)=>
      ImgReg4IN_200, D(7)=>ImgReg4IN_199, D(6)=>ImgReg4IN_198, D(5)=>
      ImgReg4IN_197, D(4)=>ImgReg4IN_196, D(3)=>ImgReg4IN_195, D(2)=>
      ImgReg4IN_194, D(1)=>ImgReg4IN_193, D(0)=>ImgReg4IN_192, CLK=>nx23904, 
      RST=>RST, EN=>nx23760, Q(15)=>OutputImg4_207_EXMPLR, Q(14)=>
      OutputImg4_206_EXMPLR, Q(13)=>OutputImg4_205_EXMPLR, Q(12)=>
      OutputImg4_204_EXMPLR, Q(11)=>OutputImg4_203_EXMPLR, Q(10)=>
      OutputImg4_202_EXMPLR, Q(9)=>OutputImg4_201_EXMPLR, Q(8)=>
      OutputImg4_200_EXMPLR, Q(7)=>OutputImg4_199_EXMPLR, Q(6)=>
      OutputImg4_198_EXMPLR, Q(5)=>OutputImg4_197_EXMPLR, Q(4)=>
      OutputImg4_196_EXMPLR, Q(3)=>OutputImg4_195_EXMPLR, Q(2)=>
      OutputImg4_194_EXMPLR, Q(1)=>OutputImg4_193_EXMPLR, Q(0)=>
      OutputImg4_192_EXMPLR);
   loop3_12_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_207, D(14)=>
      ImgReg5IN_206, D(13)=>ImgReg5IN_205, D(12)=>ImgReg5IN_204, D(11)=>
      ImgReg5IN_203, D(10)=>ImgReg5IN_202, D(9)=>ImgReg5IN_201, D(8)=>
      ImgReg5IN_200, D(7)=>ImgReg5IN_199, D(6)=>ImgReg5IN_198, D(5)=>
      ImgReg5IN_197, D(4)=>ImgReg5IN_196, D(3)=>ImgReg5IN_195, D(2)=>
      ImgReg5IN_194, D(1)=>ImgReg5IN_193, D(0)=>ImgReg5IN_192, CLK=>nx23906, 
      RST=>RST, EN=>nx23770, Q(15)=>OutputImg5_207_EXMPLR, Q(14)=>
      OutputImg5_206_EXMPLR, Q(13)=>OutputImg5_205_EXMPLR, Q(12)=>
      OutputImg5_204_EXMPLR, Q(11)=>OutputImg5_203_EXMPLR, Q(10)=>
      OutputImg5_202_EXMPLR, Q(9)=>OutputImg5_201_EXMPLR, Q(8)=>
      OutputImg5_200_EXMPLR, Q(7)=>OutputImg5_199_EXMPLR, Q(6)=>
      OutputImg5_198_EXMPLR, Q(5)=>OutputImg5_197_EXMPLR, Q(4)=>
      OutputImg5_196_EXMPLR, Q(3)=>OutputImg5_195_EXMPLR, Q(2)=>
      OutputImg5_194_EXMPLR, Q(1)=>OutputImg5_193_EXMPLR, Q(0)=>
      OutputImg5_192_EXMPLR);
   loop3_13_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_239_EXMPLR, D(14)=>OutputImg0_238_EXMPLR, D(13)=>
      OutputImg0_237_EXMPLR, D(12)=>OutputImg0_236_EXMPLR, D(11)=>
      OutputImg0_235_EXMPLR, D(10)=>OutputImg0_234_EXMPLR, D(9)=>
      OutputImg0_233_EXMPLR, D(8)=>OutputImg0_232_EXMPLR, D(7)=>
      OutputImg0_231_EXMPLR, D(6)=>OutputImg0_230_EXMPLR, D(5)=>
      OutputImg0_229_EXMPLR, D(4)=>OutputImg0_228_EXMPLR, D(3)=>
      OutputImg0_227_EXMPLR, D(2)=>OutputImg0_226_EXMPLR, D(1)=>
      OutputImg0_225_EXMPLR, D(0)=>OutputImg0_224_EXMPLR, EN=>nx23688, F(15)
      =>ImgReg0IN_223, F(14)=>ImgReg0IN_222, F(13)=>ImgReg0IN_221, F(12)=>
      ImgReg0IN_220, F(11)=>ImgReg0IN_219, F(10)=>ImgReg0IN_218, F(9)=>
      ImgReg0IN_217, F(8)=>ImgReg0IN_216, F(7)=>ImgReg0IN_215, F(6)=>
      ImgReg0IN_214, F(5)=>ImgReg0IN_213, F(4)=>ImgReg0IN_212, F(3)=>
      ImgReg0IN_211, F(2)=>ImgReg0IN_210, F(1)=>ImgReg0IN_209, F(0)=>
      ImgReg0IN_208);
   loop3_13_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_239_EXMPLR, D(14)=>OutputImg1_238_EXMPLR, D(13)=>
      OutputImg1_237_EXMPLR, D(12)=>OutputImg1_236_EXMPLR, D(11)=>
      OutputImg1_235_EXMPLR, D(10)=>OutputImg1_234_EXMPLR, D(9)=>
      OutputImg1_233_EXMPLR, D(8)=>OutputImg1_232_EXMPLR, D(7)=>
      OutputImg1_231_EXMPLR, D(6)=>OutputImg1_230_EXMPLR, D(5)=>
      OutputImg1_229_EXMPLR, D(4)=>OutputImg1_228_EXMPLR, D(3)=>
      OutputImg1_227_EXMPLR, D(2)=>OutputImg1_226_EXMPLR, D(1)=>
      OutputImg1_225_EXMPLR, D(0)=>OutputImg1_224_EXMPLR, EN=>nx23688, F(15)
      =>ImgReg1IN_223, F(14)=>ImgReg1IN_222, F(13)=>ImgReg1IN_221, F(12)=>
      ImgReg1IN_220, F(11)=>ImgReg1IN_219, F(10)=>ImgReg1IN_218, F(9)=>
      ImgReg1IN_217, F(8)=>ImgReg1IN_216, F(7)=>ImgReg1IN_215, F(6)=>
      ImgReg1IN_214, F(5)=>ImgReg1IN_213, F(4)=>ImgReg1IN_212, F(3)=>
      ImgReg1IN_211, F(2)=>ImgReg1IN_210, F(1)=>ImgReg1IN_209, F(0)=>
      ImgReg1IN_208);
   loop3_13_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_239_EXMPLR, D(14)=>OutputImg2_238_EXMPLR, D(13)=>
      OutputImg2_237_EXMPLR, D(12)=>OutputImg2_236_EXMPLR, D(11)=>
      OutputImg2_235_EXMPLR, D(10)=>OutputImg2_234_EXMPLR, D(9)=>
      OutputImg2_233_EXMPLR, D(8)=>OutputImg2_232_EXMPLR, D(7)=>
      OutputImg2_231_EXMPLR, D(6)=>OutputImg2_230_EXMPLR, D(5)=>
      OutputImg2_229_EXMPLR, D(4)=>OutputImg2_228_EXMPLR, D(3)=>
      OutputImg2_227_EXMPLR, D(2)=>OutputImg2_226_EXMPLR, D(1)=>
      OutputImg2_225_EXMPLR, D(0)=>OutputImg2_224_EXMPLR, EN=>nx23688, F(15)
      =>ImgReg2IN_223, F(14)=>ImgReg2IN_222, F(13)=>ImgReg2IN_221, F(12)=>
      ImgReg2IN_220, F(11)=>ImgReg2IN_219, F(10)=>ImgReg2IN_218, F(9)=>
      ImgReg2IN_217, F(8)=>ImgReg2IN_216, F(7)=>ImgReg2IN_215, F(6)=>
      ImgReg2IN_214, F(5)=>ImgReg2IN_213, F(4)=>ImgReg2IN_212, F(3)=>
      ImgReg2IN_211, F(2)=>ImgReg2IN_210, F(1)=>ImgReg2IN_209, F(0)=>
      ImgReg2IN_208);
   loop3_13_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_239_EXMPLR, D(14)=>OutputImg3_238_EXMPLR, D(13)=>
      OutputImg3_237_EXMPLR, D(12)=>OutputImg3_236_EXMPLR, D(11)=>
      OutputImg3_235_EXMPLR, D(10)=>OutputImg3_234_EXMPLR, D(9)=>
      OutputImg3_233_EXMPLR, D(8)=>OutputImg3_232_EXMPLR, D(7)=>
      OutputImg3_231_EXMPLR, D(6)=>OutputImg3_230_EXMPLR, D(5)=>
      OutputImg3_229_EXMPLR, D(4)=>OutputImg3_228_EXMPLR, D(3)=>
      OutputImg3_227_EXMPLR, D(2)=>OutputImg3_226_EXMPLR, D(1)=>
      OutputImg3_225_EXMPLR, D(0)=>OutputImg3_224_EXMPLR, EN=>nx23688, F(15)
      =>ImgReg3IN_223, F(14)=>ImgReg3IN_222, F(13)=>ImgReg3IN_221, F(12)=>
      ImgReg3IN_220, F(11)=>ImgReg3IN_219, F(10)=>ImgReg3IN_218, F(9)=>
      ImgReg3IN_217, F(8)=>ImgReg3IN_216, F(7)=>ImgReg3IN_215, F(6)=>
      ImgReg3IN_214, F(5)=>ImgReg3IN_213, F(4)=>ImgReg3IN_212, F(3)=>
      ImgReg3IN_211, F(2)=>ImgReg3IN_210, F(1)=>ImgReg3IN_209, F(0)=>
      ImgReg3IN_208);
   loop3_13_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_239_EXMPLR, D(14)=>OutputImg4_238_EXMPLR, D(13)=>
      OutputImg4_237_EXMPLR, D(12)=>OutputImg4_236_EXMPLR, D(11)=>
      OutputImg4_235_EXMPLR, D(10)=>OutputImg4_234_EXMPLR, D(9)=>
      OutputImg4_233_EXMPLR, D(8)=>OutputImg4_232_EXMPLR, D(7)=>
      OutputImg4_231_EXMPLR, D(6)=>OutputImg4_230_EXMPLR, D(5)=>
      OutputImg4_229_EXMPLR, D(4)=>OutputImg4_228_EXMPLR, D(3)=>
      OutputImg4_227_EXMPLR, D(2)=>OutputImg4_226_EXMPLR, D(1)=>
      OutputImg4_225_EXMPLR, D(0)=>OutputImg4_224_EXMPLR, EN=>nx23688, F(15)
      =>ImgReg4IN_223, F(14)=>ImgReg4IN_222, F(13)=>ImgReg4IN_221, F(12)=>
      ImgReg4IN_220, F(11)=>ImgReg4IN_219, F(10)=>ImgReg4IN_218, F(9)=>
      ImgReg4IN_217, F(8)=>ImgReg4IN_216, F(7)=>ImgReg4IN_215, F(6)=>
      ImgReg4IN_214, F(5)=>ImgReg4IN_213, F(4)=>ImgReg4IN_212, F(3)=>
      ImgReg4IN_211, F(2)=>ImgReg4IN_210, F(1)=>ImgReg4IN_209, F(0)=>
      ImgReg4IN_208);
   loop3_13_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_239_EXMPLR, D(14)=>OutputImg5_238_EXMPLR, D(13)=>
      OutputImg5_237_EXMPLR, D(12)=>OutputImg5_236_EXMPLR, D(11)=>
      OutputImg5_235_EXMPLR, D(10)=>OutputImg5_234_EXMPLR, D(9)=>
      OutputImg5_233_EXMPLR, D(8)=>OutputImg5_232_EXMPLR, D(7)=>
      OutputImg5_231_EXMPLR, D(6)=>OutputImg5_230_EXMPLR, D(5)=>
      OutputImg5_229_EXMPLR, D(4)=>OutputImg5_228_EXMPLR, D(3)=>
      OutputImg5_227_EXMPLR, D(2)=>OutputImg5_226_EXMPLR, D(1)=>
      OutputImg5_225_EXMPLR, D(0)=>OutputImg5_224_EXMPLR, EN=>nx23688, F(15)
      =>ImgReg5IN_223, F(14)=>ImgReg5IN_222, F(13)=>ImgReg5IN_221, F(12)=>
      ImgReg5IN_220, F(11)=>ImgReg5IN_219, F(10)=>ImgReg5IN_218, F(9)=>
      ImgReg5IN_217, F(8)=>ImgReg5IN_216, F(7)=>ImgReg5IN_215, F(6)=>
      ImgReg5IN_214, F(5)=>ImgReg5IN_213, F(4)=>ImgReg5IN_212, F(3)=>
      ImgReg5IN_211, F(2)=>ImgReg5IN_210, F(1)=>ImgReg5IN_209, F(0)=>
      ImgReg5IN_208);
   loop3_13_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(223), 
      D(14)=>DATA(222), D(13)=>DATA(221), D(12)=>DATA(220), D(11)=>DATA(219), 
      D(10)=>DATA(218), D(9)=>DATA(217), D(8)=>DATA(216), D(7)=>DATA(215), 
      D(6)=>DATA(214), D(5)=>DATA(213), D(4)=>DATA(212), D(3)=>DATA(211), 
      D(2)=>DATA(210), D(1)=>DATA(209), D(0)=>DATA(208), EN=>nx23656, F(15)
      =>ImgReg0IN_223, F(14)=>ImgReg0IN_222, F(13)=>ImgReg0IN_221, F(12)=>
      ImgReg0IN_220, F(11)=>ImgReg0IN_219, F(10)=>ImgReg0IN_218, F(9)=>
      ImgReg0IN_217, F(8)=>ImgReg0IN_216, F(7)=>ImgReg0IN_215, F(6)=>
      ImgReg0IN_214, F(5)=>ImgReg0IN_213, F(4)=>ImgReg0IN_212, F(3)=>
      ImgReg0IN_211, F(2)=>ImgReg0IN_210, F(1)=>ImgReg0IN_209, F(0)=>
      ImgReg0IN_208);
   loop3_13_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(223), 
      D(14)=>DATA(222), D(13)=>DATA(221), D(12)=>DATA(220), D(11)=>DATA(219), 
      D(10)=>DATA(218), D(9)=>DATA(217), D(8)=>DATA(216), D(7)=>DATA(215), 
      D(6)=>DATA(214), D(5)=>DATA(213), D(4)=>DATA(212), D(3)=>DATA(211), 
      D(2)=>DATA(210), D(1)=>DATA(209), D(0)=>DATA(208), EN=>nx23644, F(15)
      =>ImgReg1IN_223, F(14)=>ImgReg1IN_222, F(13)=>ImgReg1IN_221, F(12)=>
      ImgReg1IN_220, F(11)=>ImgReg1IN_219, F(10)=>ImgReg1IN_218, F(9)=>
      ImgReg1IN_217, F(8)=>ImgReg1IN_216, F(7)=>ImgReg1IN_215, F(6)=>
      ImgReg1IN_214, F(5)=>ImgReg1IN_213, F(4)=>ImgReg1IN_212, F(3)=>
      ImgReg1IN_211, F(2)=>ImgReg1IN_210, F(1)=>ImgReg1IN_209, F(0)=>
      ImgReg1IN_208);
   loop3_13_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(223), 
      D(14)=>DATA(222), D(13)=>DATA(221), D(12)=>DATA(220), D(11)=>DATA(219), 
      D(10)=>DATA(218), D(9)=>DATA(217), D(8)=>DATA(216), D(7)=>DATA(215), 
      D(6)=>DATA(214), D(5)=>DATA(213), D(4)=>DATA(212), D(3)=>DATA(211), 
      D(2)=>DATA(210), D(1)=>DATA(209), D(0)=>DATA(208), EN=>nx23632, F(15)
      =>ImgReg2IN_223, F(14)=>ImgReg2IN_222, F(13)=>ImgReg2IN_221, F(12)=>
      ImgReg2IN_220, F(11)=>ImgReg2IN_219, F(10)=>ImgReg2IN_218, F(9)=>
      ImgReg2IN_217, F(8)=>ImgReg2IN_216, F(7)=>ImgReg2IN_215, F(6)=>
      ImgReg2IN_214, F(5)=>ImgReg2IN_213, F(4)=>ImgReg2IN_212, F(3)=>
      ImgReg2IN_211, F(2)=>ImgReg2IN_210, F(1)=>ImgReg2IN_209, F(0)=>
      ImgReg2IN_208);
   loop3_13_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(223), 
      D(14)=>DATA(222), D(13)=>DATA(221), D(12)=>DATA(220), D(11)=>DATA(219), 
      D(10)=>DATA(218), D(9)=>DATA(217), D(8)=>DATA(216), D(7)=>DATA(215), 
      D(6)=>DATA(214), D(5)=>DATA(213), D(4)=>DATA(212), D(3)=>DATA(211), 
      D(2)=>DATA(210), D(1)=>DATA(209), D(0)=>DATA(208), EN=>nx23620, F(15)
      =>ImgReg3IN_223, F(14)=>ImgReg3IN_222, F(13)=>ImgReg3IN_221, F(12)=>
      ImgReg3IN_220, F(11)=>ImgReg3IN_219, F(10)=>ImgReg3IN_218, F(9)=>
      ImgReg3IN_217, F(8)=>ImgReg3IN_216, F(7)=>ImgReg3IN_215, F(6)=>
      ImgReg3IN_214, F(5)=>ImgReg3IN_213, F(4)=>ImgReg3IN_212, F(3)=>
      ImgReg3IN_211, F(2)=>ImgReg3IN_210, F(1)=>ImgReg3IN_209, F(0)=>
      ImgReg3IN_208);
   loop3_13_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(223), 
      D(14)=>DATA(222), D(13)=>DATA(221), D(12)=>DATA(220), D(11)=>DATA(219), 
      D(10)=>DATA(218), D(9)=>DATA(217), D(8)=>DATA(216), D(7)=>DATA(215), 
      D(6)=>DATA(214), D(5)=>DATA(213), D(4)=>DATA(212), D(3)=>DATA(211), 
      D(2)=>DATA(210), D(1)=>DATA(209), D(0)=>DATA(208), EN=>nx23608, F(15)
      =>ImgReg4IN_223, F(14)=>ImgReg4IN_222, F(13)=>ImgReg4IN_221, F(12)=>
      ImgReg4IN_220, F(11)=>ImgReg4IN_219, F(10)=>ImgReg4IN_218, F(9)=>
      ImgReg4IN_217, F(8)=>ImgReg4IN_216, F(7)=>ImgReg4IN_215, F(6)=>
      ImgReg4IN_214, F(5)=>ImgReg4IN_213, F(4)=>ImgReg4IN_212, F(3)=>
      ImgReg4IN_211, F(2)=>ImgReg4IN_210, F(1)=>ImgReg4IN_209, F(0)=>
      ImgReg4IN_208);
   loop3_13_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(223), 
      D(14)=>DATA(222), D(13)=>DATA(221), D(12)=>DATA(220), D(11)=>DATA(219), 
      D(10)=>DATA(218), D(9)=>DATA(217), D(8)=>DATA(216), D(7)=>DATA(215), 
      D(6)=>DATA(214), D(5)=>DATA(213), D(4)=>DATA(212), D(3)=>DATA(211), 
      D(2)=>DATA(210), D(1)=>DATA(209), D(0)=>DATA(208), EN=>nx23596, F(15)
      =>ImgReg5IN_223, F(14)=>ImgReg5IN_222, F(13)=>ImgReg5IN_221, F(12)=>
      ImgReg5IN_220, F(11)=>ImgReg5IN_219, F(10)=>ImgReg5IN_218, F(9)=>
      ImgReg5IN_217, F(8)=>ImgReg5IN_216, F(7)=>ImgReg5IN_215, F(6)=>
      ImgReg5IN_214, F(5)=>ImgReg5IN_213, F(4)=>ImgReg5IN_212, F(3)=>
      ImgReg5IN_211, F(2)=>ImgReg5IN_210, F(1)=>ImgReg5IN_209, F(0)=>
      ImgReg5IN_208);
   loop3_13_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_223_EXMPLR, D(14)=>OutputImg1_222_EXMPLR, D(13)=>
      OutputImg1_221_EXMPLR, D(12)=>OutputImg1_220_EXMPLR, D(11)=>
      OutputImg1_219_EXMPLR, D(10)=>OutputImg1_218_EXMPLR, D(9)=>
      OutputImg1_217_EXMPLR, D(8)=>OutputImg1_216_EXMPLR, D(7)=>
      OutputImg1_215_EXMPLR, D(6)=>OutputImg1_214_EXMPLR, D(5)=>
      OutputImg1_213_EXMPLR, D(4)=>OutputImg1_212_EXMPLR, D(3)=>
      OutputImg1_211_EXMPLR, D(2)=>OutputImg1_210_EXMPLR, D(1)=>
      OutputImg1_209_EXMPLR, D(0)=>OutputImg1_208_EXMPLR, EN=>nx23804, F(15)
      =>ImgReg0IN_223, F(14)=>ImgReg0IN_222, F(13)=>ImgReg0IN_221, F(12)=>
      ImgReg0IN_220, F(11)=>ImgReg0IN_219, F(10)=>ImgReg0IN_218, F(9)=>
      ImgReg0IN_217, F(8)=>ImgReg0IN_216, F(7)=>ImgReg0IN_215, F(6)=>
      ImgReg0IN_214, F(5)=>ImgReg0IN_213, F(4)=>ImgReg0IN_212, F(3)=>
      ImgReg0IN_211, F(2)=>ImgReg0IN_210, F(1)=>ImgReg0IN_209, F(0)=>
      ImgReg0IN_208);
   loop3_13_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_223_EXMPLR, D(14)=>OutputImg2_222_EXMPLR, D(13)=>
      OutputImg2_221_EXMPLR, D(12)=>OutputImg2_220_EXMPLR, D(11)=>
      OutputImg2_219_EXMPLR, D(10)=>OutputImg2_218_EXMPLR, D(9)=>
      OutputImg2_217_EXMPLR, D(8)=>OutputImg2_216_EXMPLR, D(7)=>
      OutputImg2_215_EXMPLR, D(6)=>OutputImg2_214_EXMPLR, D(5)=>
      OutputImg2_213_EXMPLR, D(4)=>OutputImg2_212_EXMPLR, D(3)=>
      OutputImg2_211_EXMPLR, D(2)=>OutputImg2_210_EXMPLR, D(1)=>
      OutputImg2_209_EXMPLR, D(0)=>OutputImg2_208_EXMPLR, EN=>nx23804, F(15)
      =>ImgReg1IN_223, F(14)=>ImgReg1IN_222, F(13)=>ImgReg1IN_221, F(12)=>
      ImgReg1IN_220, F(11)=>ImgReg1IN_219, F(10)=>ImgReg1IN_218, F(9)=>
      ImgReg1IN_217, F(8)=>ImgReg1IN_216, F(7)=>ImgReg1IN_215, F(6)=>
      ImgReg1IN_214, F(5)=>ImgReg1IN_213, F(4)=>ImgReg1IN_212, F(3)=>
      ImgReg1IN_211, F(2)=>ImgReg1IN_210, F(1)=>ImgReg1IN_209, F(0)=>
      ImgReg1IN_208);
   loop3_13_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_223_EXMPLR, D(14)=>OutputImg3_222_EXMPLR, D(13)=>
      OutputImg3_221_EXMPLR, D(12)=>OutputImg3_220_EXMPLR, D(11)=>
      OutputImg3_219_EXMPLR, D(10)=>OutputImg3_218_EXMPLR, D(9)=>
      OutputImg3_217_EXMPLR, D(8)=>OutputImg3_216_EXMPLR, D(7)=>
      OutputImg3_215_EXMPLR, D(6)=>OutputImg3_214_EXMPLR, D(5)=>
      OutputImg3_213_EXMPLR, D(4)=>OutputImg3_212_EXMPLR, D(3)=>
      OutputImg3_211_EXMPLR, D(2)=>OutputImg3_210_EXMPLR, D(1)=>
      OutputImg3_209_EXMPLR, D(0)=>OutputImg3_208_EXMPLR, EN=>nx23804, F(15)
      =>ImgReg2IN_223, F(14)=>ImgReg2IN_222, F(13)=>ImgReg2IN_221, F(12)=>
      ImgReg2IN_220, F(11)=>ImgReg2IN_219, F(10)=>ImgReg2IN_218, F(9)=>
      ImgReg2IN_217, F(8)=>ImgReg2IN_216, F(7)=>ImgReg2IN_215, F(6)=>
      ImgReg2IN_214, F(5)=>ImgReg2IN_213, F(4)=>ImgReg2IN_212, F(3)=>
      ImgReg2IN_211, F(2)=>ImgReg2IN_210, F(1)=>ImgReg2IN_209, F(0)=>
      ImgReg2IN_208);
   loop3_13_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_223_EXMPLR, D(14)=>OutputImg4_222_EXMPLR, D(13)=>
      OutputImg4_221_EXMPLR, D(12)=>OutputImg4_220_EXMPLR, D(11)=>
      OutputImg4_219_EXMPLR, D(10)=>OutputImg4_218_EXMPLR, D(9)=>
      OutputImg4_217_EXMPLR, D(8)=>OutputImg4_216_EXMPLR, D(7)=>
      OutputImg4_215_EXMPLR, D(6)=>OutputImg4_214_EXMPLR, D(5)=>
      OutputImg4_213_EXMPLR, D(4)=>OutputImg4_212_EXMPLR, D(3)=>
      OutputImg4_211_EXMPLR, D(2)=>OutputImg4_210_EXMPLR, D(1)=>
      OutputImg4_209_EXMPLR, D(0)=>OutputImg4_208_EXMPLR, EN=>nx23804, F(15)
      =>ImgReg3IN_223, F(14)=>ImgReg3IN_222, F(13)=>ImgReg3IN_221, F(12)=>
      ImgReg3IN_220, F(11)=>ImgReg3IN_219, F(10)=>ImgReg3IN_218, F(9)=>
      ImgReg3IN_217, F(8)=>ImgReg3IN_216, F(7)=>ImgReg3IN_215, F(6)=>
      ImgReg3IN_214, F(5)=>ImgReg3IN_213, F(4)=>ImgReg3IN_212, F(3)=>
      ImgReg3IN_211, F(2)=>ImgReg3IN_210, F(1)=>ImgReg3IN_209, F(0)=>
      ImgReg3IN_208);
   loop3_13_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_223_EXMPLR, D(14)=>OutputImg5_222_EXMPLR, D(13)=>
      OutputImg5_221_EXMPLR, D(12)=>OutputImg5_220_EXMPLR, D(11)=>
      OutputImg5_219_EXMPLR, D(10)=>OutputImg5_218_EXMPLR, D(9)=>
      OutputImg5_217_EXMPLR, D(8)=>OutputImg5_216_EXMPLR, D(7)=>
      OutputImg5_215_EXMPLR, D(6)=>OutputImg5_214_EXMPLR, D(5)=>
      OutputImg5_213_EXMPLR, D(4)=>OutputImg5_212_EXMPLR, D(3)=>
      OutputImg5_211_EXMPLR, D(2)=>OutputImg5_210_EXMPLR, D(1)=>
      OutputImg5_209_EXMPLR, D(0)=>OutputImg5_208_EXMPLR, EN=>nx23804, F(15)
      =>ImgReg4IN_223, F(14)=>ImgReg4IN_222, F(13)=>ImgReg4IN_221, F(12)=>
      ImgReg4IN_220, F(11)=>ImgReg4IN_219, F(10)=>ImgReg4IN_218, F(9)=>
      ImgReg4IN_217, F(8)=>ImgReg4IN_216, F(7)=>ImgReg4IN_215, F(6)=>
      ImgReg4IN_214, F(5)=>ImgReg4IN_213, F(4)=>ImgReg4IN_212, F(3)=>
      ImgReg4IN_211, F(2)=>ImgReg4IN_210, F(1)=>ImgReg4IN_209, F(0)=>
      ImgReg4IN_208);
   loop3_13_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_223, D(14)=>
      ImgReg0IN_222, D(13)=>ImgReg0IN_221, D(12)=>ImgReg0IN_220, D(11)=>
      ImgReg0IN_219, D(10)=>ImgReg0IN_218, D(9)=>ImgReg0IN_217, D(8)=>
      ImgReg0IN_216, D(7)=>ImgReg0IN_215, D(6)=>ImgReg0IN_214, D(5)=>
      ImgReg0IN_213, D(4)=>ImgReg0IN_212, D(3)=>ImgReg0IN_211, D(2)=>
      ImgReg0IN_210, D(1)=>ImgReg0IN_209, D(0)=>ImgReg0IN_208, CLK=>nx23906, 
      RST=>RST, EN=>nx23720, Q(15)=>OutputImg0_223_EXMPLR, Q(14)=>
      OutputImg0_222_EXMPLR, Q(13)=>OutputImg0_221_EXMPLR, Q(12)=>
      OutputImg0_220_EXMPLR, Q(11)=>OutputImg0_219_EXMPLR, Q(10)=>
      OutputImg0_218_EXMPLR, Q(9)=>OutputImg0_217_EXMPLR, Q(8)=>
      OutputImg0_216_EXMPLR, Q(7)=>OutputImg0_215_EXMPLR, Q(6)=>
      OutputImg0_214_EXMPLR, Q(5)=>OutputImg0_213_EXMPLR, Q(4)=>
      OutputImg0_212_EXMPLR, Q(3)=>OutputImg0_211_EXMPLR, Q(2)=>
      OutputImg0_210_EXMPLR, Q(1)=>OutputImg0_209_EXMPLR, Q(0)=>
      OutputImg0_208_EXMPLR);
   loop3_13_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_223, D(14)=>
      ImgReg1IN_222, D(13)=>ImgReg1IN_221, D(12)=>ImgReg1IN_220, D(11)=>
      ImgReg1IN_219, D(10)=>ImgReg1IN_218, D(9)=>ImgReg1IN_217, D(8)=>
      ImgReg1IN_216, D(7)=>ImgReg1IN_215, D(6)=>ImgReg1IN_214, D(5)=>
      ImgReg1IN_213, D(4)=>ImgReg1IN_212, D(3)=>ImgReg1IN_211, D(2)=>
      ImgReg1IN_210, D(1)=>ImgReg1IN_209, D(0)=>ImgReg1IN_208, CLK=>nx23908, 
      RST=>RST, EN=>nx23730, Q(15)=>OutputImg1_223_EXMPLR, Q(14)=>
      OutputImg1_222_EXMPLR, Q(13)=>OutputImg1_221_EXMPLR, Q(12)=>
      OutputImg1_220_EXMPLR, Q(11)=>OutputImg1_219_EXMPLR, Q(10)=>
      OutputImg1_218_EXMPLR, Q(9)=>OutputImg1_217_EXMPLR, Q(8)=>
      OutputImg1_216_EXMPLR, Q(7)=>OutputImg1_215_EXMPLR, Q(6)=>
      OutputImg1_214_EXMPLR, Q(5)=>OutputImg1_213_EXMPLR, Q(4)=>
      OutputImg1_212_EXMPLR, Q(3)=>OutputImg1_211_EXMPLR, Q(2)=>
      OutputImg1_210_EXMPLR, Q(1)=>OutputImg1_209_EXMPLR, Q(0)=>
      OutputImg1_208_EXMPLR);
   loop3_13_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_223, D(14)=>
      ImgReg2IN_222, D(13)=>ImgReg2IN_221, D(12)=>ImgReg2IN_220, D(11)=>
      ImgReg2IN_219, D(10)=>ImgReg2IN_218, D(9)=>ImgReg2IN_217, D(8)=>
      ImgReg2IN_216, D(7)=>ImgReg2IN_215, D(6)=>ImgReg2IN_214, D(5)=>
      ImgReg2IN_213, D(4)=>ImgReg2IN_212, D(3)=>ImgReg2IN_211, D(2)=>
      ImgReg2IN_210, D(1)=>ImgReg2IN_209, D(0)=>ImgReg2IN_208, CLK=>nx23908, 
      RST=>RST, EN=>nx23740, Q(15)=>OutputImg2_223_EXMPLR, Q(14)=>
      OutputImg2_222_EXMPLR, Q(13)=>OutputImg2_221_EXMPLR, Q(12)=>
      OutputImg2_220_EXMPLR, Q(11)=>OutputImg2_219_EXMPLR, Q(10)=>
      OutputImg2_218_EXMPLR, Q(9)=>OutputImg2_217_EXMPLR, Q(8)=>
      OutputImg2_216_EXMPLR, Q(7)=>OutputImg2_215_EXMPLR, Q(6)=>
      OutputImg2_214_EXMPLR, Q(5)=>OutputImg2_213_EXMPLR, Q(4)=>
      OutputImg2_212_EXMPLR, Q(3)=>OutputImg2_211_EXMPLR, Q(2)=>
      OutputImg2_210_EXMPLR, Q(1)=>OutputImg2_209_EXMPLR, Q(0)=>
      OutputImg2_208_EXMPLR);
   loop3_13_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_223, D(14)=>
      ImgReg3IN_222, D(13)=>ImgReg3IN_221, D(12)=>ImgReg3IN_220, D(11)=>
      ImgReg3IN_219, D(10)=>ImgReg3IN_218, D(9)=>ImgReg3IN_217, D(8)=>
      ImgReg3IN_216, D(7)=>ImgReg3IN_215, D(6)=>ImgReg3IN_214, D(5)=>
      ImgReg3IN_213, D(4)=>ImgReg3IN_212, D(3)=>ImgReg3IN_211, D(2)=>
      ImgReg3IN_210, D(1)=>ImgReg3IN_209, D(0)=>ImgReg3IN_208, CLK=>nx23910, 
      RST=>RST, EN=>nx23750, Q(15)=>OutputImg3_223_EXMPLR, Q(14)=>
      OutputImg3_222_EXMPLR, Q(13)=>OutputImg3_221_EXMPLR, Q(12)=>
      OutputImg3_220_EXMPLR, Q(11)=>OutputImg3_219_EXMPLR, Q(10)=>
      OutputImg3_218_EXMPLR, Q(9)=>OutputImg3_217_EXMPLR, Q(8)=>
      OutputImg3_216_EXMPLR, Q(7)=>OutputImg3_215_EXMPLR, Q(6)=>
      OutputImg3_214_EXMPLR, Q(5)=>OutputImg3_213_EXMPLR, Q(4)=>
      OutputImg3_212_EXMPLR, Q(3)=>OutputImg3_211_EXMPLR, Q(2)=>
      OutputImg3_210_EXMPLR, Q(1)=>OutputImg3_209_EXMPLR, Q(0)=>
      OutputImg3_208_EXMPLR);
   loop3_13_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_223, D(14)=>
      ImgReg4IN_222, D(13)=>ImgReg4IN_221, D(12)=>ImgReg4IN_220, D(11)=>
      ImgReg4IN_219, D(10)=>ImgReg4IN_218, D(9)=>ImgReg4IN_217, D(8)=>
      ImgReg4IN_216, D(7)=>ImgReg4IN_215, D(6)=>ImgReg4IN_214, D(5)=>
      ImgReg4IN_213, D(4)=>ImgReg4IN_212, D(3)=>ImgReg4IN_211, D(2)=>
      ImgReg4IN_210, D(1)=>ImgReg4IN_209, D(0)=>ImgReg4IN_208, CLK=>nx23910, 
      RST=>RST, EN=>nx23760, Q(15)=>OutputImg4_223_EXMPLR, Q(14)=>
      OutputImg4_222_EXMPLR, Q(13)=>OutputImg4_221_EXMPLR, Q(12)=>
      OutputImg4_220_EXMPLR, Q(11)=>OutputImg4_219_EXMPLR, Q(10)=>
      OutputImg4_218_EXMPLR, Q(9)=>OutputImg4_217_EXMPLR, Q(8)=>
      OutputImg4_216_EXMPLR, Q(7)=>OutputImg4_215_EXMPLR, Q(6)=>
      OutputImg4_214_EXMPLR, Q(5)=>OutputImg4_213_EXMPLR, Q(4)=>
      OutputImg4_212_EXMPLR, Q(3)=>OutputImg4_211_EXMPLR, Q(2)=>
      OutputImg4_210_EXMPLR, Q(1)=>OutputImg4_209_EXMPLR, Q(0)=>
      OutputImg4_208_EXMPLR);
   loop3_13_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_223, D(14)=>
      ImgReg5IN_222, D(13)=>ImgReg5IN_221, D(12)=>ImgReg5IN_220, D(11)=>
      ImgReg5IN_219, D(10)=>ImgReg5IN_218, D(9)=>ImgReg5IN_217, D(8)=>
      ImgReg5IN_216, D(7)=>ImgReg5IN_215, D(6)=>ImgReg5IN_214, D(5)=>
      ImgReg5IN_213, D(4)=>ImgReg5IN_212, D(3)=>ImgReg5IN_211, D(2)=>
      ImgReg5IN_210, D(1)=>ImgReg5IN_209, D(0)=>ImgReg5IN_208, CLK=>nx23912, 
      RST=>RST, EN=>nx23770, Q(15)=>OutputImg5_223_EXMPLR, Q(14)=>
      OutputImg5_222_EXMPLR, Q(13)=>OutputImg5_221_EXMPLR, Q(12)=>
      OutputImg5_220_EXMPLR, Q(11)=>OutputImg5_219_EXMPLR, Q(10)=>
      OutputImg5_218_EXMPLR, Q(9)=>OutputImg5_217_EXMPLR, Q(8)=>
      OutputImg5_216_EXMPLR, Q(7)=>OutputImg5_215_EXMPLR, Q(6)=>
      OutputImg5_214_EXMPLR, Q(5)=>OutputImg5_213_EXMPLR, Q(4)=>
      OutputImg5_212_EXMPLR, Q(3)=>OutputImg5_211_EXMPLR, Q(2)=>
      OutputImg5_210_EXMPLR, Q(1)=>OutputImg5_209_EXMPLR, Q(0)=>
      OutputImg5_208_EXMPLR);
   loop3_14_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_255_EXMPLR, D(14)=>OutputImg0_254_EXMPLR, D(13)=>
      OutputImg0_253_EXMPLR, D(12)=>OutputImg0_252_EXMPLR, D(11)=>
      OutputImg0_251_EXMPLR, D(10)=>OutputImg0_250_EXMPLR, D(9)=>
      OutputImg0_249_EXMPLR, D(8)=>OutputImg0_248_EXMPLR, D(7)=>
      OutputImg0_247_EXMPLR, D(6)=>OutputImg0_246_EXMPLR, D(5)=>
      OutputImg0_245_EXMPLR, D(4)=>OutputImg0_244_EXMPLR, D(3)=>
      OutputImg0_243_EXMPLR, D(2)=>OutputImg0_242_EXMPLR, D(1)=>
      OutputImg0_241_EXMPLR, D(0)=>OutputImg0_240_EXMPLR, EN=>nx23690, F(15)
      =>ImgReg0IN_239, F(14)=>ImgReg0IN_238, F(13)=>ImgReg0IN_237, F(12)=>
      ImgReg0IN_236, F(11)=>ImgReg0IN_235, F(10)=>ImgReg0IN_234, F(9)=>
      ImgReg0IN_233, F(8)=>ImgReg0IN_232, F(7)=>ImgReg0IN_231, F(6)=>
      ImgReg0IN_230, F(5)=>ImgReg0IN_229, F(4)=>ImgReg0IN_228, F(3)=>
      ImgReg0IN_227, F(2)=>ImgReg0IN_226, F(1)=>ImgReg0IN_225, F(0)=>
      ImgReg0IN_224);
   loop3_14_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_255_EXMPLR, D(14)=>OutputImg1_254_EXMPLR, D(13)=>
      OutputImg1_253_EXMPLR, D(12)=>OutputImg1_252_EXMPLR, D(11)=>
      OutputImg1_251_EXMPLR, D(10)=>OutputImg1_250_EXMPLR, D(9)=>
      OutputImg1_249_EXMPLR, D(8)=>OutputImg1_248_EXMPLR, D(7)=>
      OutputImg1_247_EXMPLR, D(6)=>OutputImg1_246_EXMPLR, D(5)=>
      OutputImg1_245_EXMPLR, D(4)=>OutputImg1_244_EXMPLR, D(3)=>
      OutputImg1_243_EXMPLR, D(2)=>OutputImg1_242_EXMPLR, D(1)=>
      OutputImg1_241_EXMPLR, D(0)=>OutputImg1_240_EXMPLR, EN=>nx23690, F(15)
      =>ImgReg1IN_239, F(14)=>ImgReg1IN_238, F(13)=>ImgReg1IN_237, F(12)=>
      ImgReg1IN_236, F(11)=>ImgReg1IN_235, F(10)=>ImgReg1IN_234, F(9)=>
      ImgReg1IN_233, F(8)=>ImgReg1IN_232, F(7)=>ImgReg1IN_231, F(6)=>
      ImgReg1IN_230, F(5)=>ImgReg1IN_229, F(4)=>ImgReg1IN_228, F(3)=>
      ImgReg1IN_227, F(2)=>ImgReg1IN_226, F(1)=>ImgReg1IN_225, F(0)=>
      ImgReg1IN_224);
   loop3_14_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_255_EXMPLR, D(14)=>OutputImg2_254_EXMPLR, D(13)=>
      OutputImg2_253_EXMPLR, D(12)=>OutputImg2_252_EXMPLR, D(11)=>
      OutputImg2_251_EXMPLR, D(10)=>OutputImg2_250_EXMPLR, D(9)=>
      OutputImg2_249_EXMPLR, D(8)=>OutputImg2_248_EXMPLR, D(7)=>
      OutputImg2_247_EXMPLR, D(6)=>OutputImg2_246_EXMPLR, D(5)=>
      OutputImg2_245_EXMPLR, D(4)=>OutputImg2_244_EXMPLR, D(3)=>
      OutputImg2_243_EXMPLR, D(2)=>OutputImg2_242_EXMPLR, D(1)=>
      OutputImg2_241_EXMPLR, D(0)=>OutputImg2_240_EXMPLR, EN=>nx23690, F(15)
      =>ImgReg2IN_239, F(14)=>ImgReg2IN_238, F(13)=>ImgReg2IN_237, F(12)=>
      ImgReg2IN_236, F(11)=>ImgReg2IN_235, F(10)=>ImgReg2IN_234, F(9)=>
      ImgReg2IN_233, F(8)=>ImgReg2IN_232, F(7)=>ImgReg2IN_231, F(6)=>
      ImgReg2IN_230, F(5)=>ImgReg2IN_229, F(4)=>ImgReg2IN_228, F(3)=>
      ImgReg2IN_227, F(2)=>ImgReg2IN_226, F(1)=>ImgReg2IN_225, F(0)=>
      ImgReg2IN_224);
   loop3_14_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_255_EXMPLR, D(14)=>OutputImg3_254_EXMPLR, D(13)=>
      OutputImg3_253_EXMPLR, D(12)=>OutputImg3_252_EXMPLR, D(11)=>
      OutputImg3_251_EXMPLR, D(10)=>OutputImg3_250_EXMPLR, D(9)=>
      OutputImg3_249_EXMPLR, D(8)=>OutputImg3_248_EXMPLR, D(7)=>
      OutputImg3_247_EXMPLR, D(6)=>OutputImg3_246_EXMPLR, D(5)=>
      OutputImg3_245_EXMPLR, D(4)=>OutputImg3_244_EXMPLR, D(3)=>
      OutputImg3_243_EXMPLR, D(2)=>OutputImg3_242_EXMPLR, D(1)=>
      OutputImg3_241_EXMPLR, D(0)=>OutputImg3_240_EXMPLR, EN=>nx23690, F(15)
      =>ImgReg3IN_239, F(14)=>ImgReg3IN_238, F(13)=>ImgReg3IN_237, F(12)=>
      ImgReg3IN_236, F(11)=>ImgReg3IN_235, F(10)=>ImgReg3IN_234, F(9)=>
      ImgReg3IN_233, F(8)=>ImgReg3IN_232, F(7)=>ImgReg3IN_231, F(6)=>
      ImgReg3IN_230, F(5)=>ImgReg3IN_229, F(4)=>ImgReg3IN_228, F(3)=>
      ImgReg3IN_227, F(2)=>ImgReg3IN_226, F(1)=>ImgReg3IN_225, F(0)=>
      ImgReg3IN_224);
   loop3_14_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_255_EXMPLR, D(14)=>OutputImg4_254_EXMPLR, D(13)=>
      OutputImg4_253_EXMPLR, D(12)=>OutputImg4_252_EXMPLR, D(11)=>
      OutputImg4_251_EXMPLR, D(10)=>OutputImg4_250_EXMPLR, D(9)=>
      OutputImg4_249_EXMPLR, D(8)=>OutputImg4_248_EXMPLR, D(7)=>
      OutputImg4_247_EXMPLR, D(6)=>OutputImg4_246_EXMPLR, D(5)=>
      OutputImg4_245_EXMPLR, D(4)=>OutputImg4_244_EXMPLR, D(3)=>
      OutputImg4_243_EXMPLR, D(2)=>OutputImg4_242_EXMPLR, D(1)=>
      OutputImg4_241_EXMPLR, D(0)=>OutputImg4_240_EXMPLR, EN=>nx23690, F(15)
      =>ImgReg4IN_239, F(14)=>ImgReg4IN_238, F(13)=>ImgReg4IN_237, F(12)=>
      ImgReg4IN_236, F(11)=>ImgReg4IN_235, F(10)=>ImgReg4IN_234, F(9)=>
      ImgReg4IN_233, F(8)=>ImgReg4IN_232, F(7)=>ImgReg4IN_231, F(6)=>
      ImgReg4IN_230, F(5)=>ImgReg4IN_229, F(4)=>ImgReg4IN_228, F(3)=>
      ImgReg4IN_227, F(2)=>ImgReg4IN_226, F(1)=>ImgReg4IN_225, F(0)=>
      ImgReg4IN_224);
   loop3_14_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_255_EXMPLR, D(14)=>OutputImg5_254_EXMPLR, D(13)=>
      OutputImg5_253_EXMPLR, D(12)=>OutputImg5_252_EXMPLR, D(11)=>
      OutputImg5_251_EXMPLR, D(10)=>OutputImg5_250_EXMPLR, D(9)=>
      OutputImg5_249_EXMPLR, D(8)=>OutputImg5_248_EXMPLR, D(7)=>
      OutputImg5_247_EXMPLR, D(6)=>OutputImg5_246_EXMPLR, D(5)=>
      OutputImg5_245_EXMPLR, D(4)=>OutputImg5_244_EXMPLR, D(3)=>
      OutputImg5_243_EXMPLR, D(2)=>OutputImg5_242_EXMPLR, D(1)=>
      OutputImg5_241_EXMPLR, D(0)=>OutputImg5_240_EXMPLR, EN=>nx23690, F(15)
      =>ImgReg5IN_239, F(14)=>ImgReg5IN_238, F(13)=>ImgReg5IN_237, F(12)=>
      ImgReg5IN_236, F(11)=>ImgReg5IN_235, F(10)=>ImgReg5IN_234, F(9)=>
      ImgReg5IN_233, F(8)=>ImgReg5IN_232, F(7)=>ImgReg5IN_231, F(6)=>
      ImgReg5IN_230, F(5)=>ImgReg5IN_229, F(4)=>ImgReg5IN_228, F(3)=>
      ImgReg5IN_227, F(2)=>ImgReg5IN_226, F(1)=>ImgReg5IN_225, F(0)=>
      ImgReg5IN_224);
   loop3_14_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(239), 
      D(14)=>DATA(238), D(13)=>DATA(237), D(12)=>DATA(236), D(11)=>DATA(235), 
      D(10)=>DATA(234), D(9)=>DATA(233), D(8)=>DATA(232), D(7)=>DATA(231), 
      D(6)=>DATA(230), D(5)=>DATA(229), D(4)=>DATA(228), D(3)=>DATA(227), 
      D(2)=>DATA(226), D(1)=>DATA(225), D(0)=>DATA(224), EN=>nx23658, F(15)
      =>ImgReg0IN_239, F(14)=>ImgReg0IN_238, F(13)=>ImgReg0IN_237, F(12)=>
      ImgReg0IN_236, F(11)=>ImgReg0IN_235, F(10)=>ImgReg0IN_234, F(9)=>
      ImgReg0IN_233, F(8)=>ImgReg0IN_232, F(7)=>ImgReg0IN_231, F(6)=>
      ImgReg0IN_230, F(5)=>ImgReg0IN_229, F(4)=>ImgReg0IN_228, F(3)=>
      ImgReg0IN_227, F(2)=>ImgReg0IN_226, F(1)=>ImgReg0IN_225, F(0)=>
      ImgReg0IN_224);
   loop3_14_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(239), 
      D(14)=>DATA(238), D(13)=>DATA(237), D(12)=>DATA(236), D(11)=>DATA(235), 
      D(10)=>DATA(234), D(9)=>DATA(233), D(8)=>DATA(232), D(7)=>DATA(231), 
      D(6)=>DATA(230), D(5)=>DATA(229), D(4)=>DATA(228), D(3)=>DATA(227), 
      D(2)=>DATA(226), D(1)=>DATA(225), D(0)=>DATA(224), EN=>nx23646, F(15)
      =>ImgReg1IN_239, F(14)=>ImgReg1IN_238, F(13)=>ImgReg1IN_237, F(12)=>
      ImgReg1IN_236, F(11)=>ImgReg1IN_235, F(10)=>ImgReg1IN_234, F(9)=>
      ImgReg1IN_233, F(8)=>ImgReg1IN_232, F(7)=>ImgReg1IN_231, F(6)=>
      ImgReg1IN_230, F(5)=>ImgReg1IN_229, F(4)=>ImgReg1IN_228, F(3)=>
      ImgReg1IN_227, F(2)=>ImgReg1IN_226, F(1)=>ImgReg1IN_225, F(0)=>
      ImgReg1IN_224);
   loop3_14_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(239), 
      D(14)=>DATA(238), D(13)=>DATA(237), D(12)=>DATA(236), D(11)=>DATA(235), 
      D(10)=>DATA(234), D(9)=>DATA(233), D(8)=>DATA(232), D(7)=>DATA(231), 
      D(6)=>DATA(230), D(5)=>DATA(229), D(4)=>DATA(228), D(3)=>DATA(227), 
      D(2)=>DATA(226), D(1)=>DATA(225), D(0)=>DATA(224), EN=>nx23634, F(15)
      =>ImgReg2IN_239, F(14)=>ImgReg2IN_238, F(13)=>ImgReg2IN_237, F(12)=>
      ImgReg2IN_236, F(11)=>ImgReg2IN_235, F(10)=>ImgReg2IN_234, F(9)=>
      ImgReg2IN_233, F(8)=>ImgReg2IN_232, F(7)=>ImgReg2IN_231, F(6)=>
      ImgReg2IN_230, F(5)=>ImgReg2IN_229, F(4)=>ImgReg2IN_228, F(3)=>
      ImgReg2IN_227, F(2)=>ImgReg2IN_226, F(1)=>ImgReg2IN_225, F(0)=>
      ImgReg2IN_224);
   loop3_14_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(239), 
      D(14)=>DATA(238), D(13)=>DATA(237), D(12)=>DATA(236), D(11)=>DATA(235), 
      D(10)=>DATA(234), D(9)=>DATA(233), D(8)=>DATA(232), D(7)=>DATA(231), 
      D(6)=>DATA(230), D(5)=>DATA(229), D(4)=>DATA(228), D(3)=>DATA(227), 
      D(2)=>DATA(226), D(1)=>DATA(225), D(0)=>DATA(224), EN=>nx23622, F(15)
      =>ImgReg3IN_239, F(14)=>ImgReg3IN_238, F(13)=>ImgReg3IN_237, F(12)=>
      ImgReg3IN_236, F(11)=>ImgReg3IN_235, F(10)=>ImgReg3IN_234, F(9)=>
      ImgReg3IN_233, F(8)=>ImgReg3IN_232, F(7)=>ImgReg3IN_231, F(6)=>
      ImgReg3IN_230, F(5)=>ImgReg3IN_229, F(4)=>ImgReg3IN_228, F(3)=>
      ImgReg3IN_227, F(2)=>ImgReg3IN_226, F(1)=>ImgReg3IN_225, F(0)=>
      ImgReg3IN_224);
   loop3_14_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(239), 
      D(14)=>DATA(238), D(13)=>DATA(237), D(12)=>DATA(236), D(11)=>DATA(235), 
      D(10)=>DATA(234), D(9)=>DATA(233), D(8)=>DATA(232), D(7)=>DATA(231), 
      D(6)=>DATA(230), D(5)=>DATA(229), D(4)=>DATA(228), D(3)=>DATA(227), 
      D(2)=>DATA(226), D(1)=>DATA(225), D(0)=>DATA(224), EN=>nx23610, F(15)
      =>ImgReg4IN_239, F(14)=>ImgReg4IN_238, F(13)=>ImgReg4IN_237, F(12)=>
      ImgReg4IN_236, F(11)=>ImgReg4IN_235, F(10)=>ImgReg4IN_234, F(9)=>
      ImgReg4IN_233, F(8)=>ImgReg4IN_232, F(7)=>ImgReg4IN_231, F(6)=>
      ImgReg4IN_230, F(5)=>ImgReg4IN_229, F(4)=>ImgReg4IN_228, F(3)=>
      ImgReg4IN_227, F(2)=>ImgReg4IN_226, F(1)=>ImgReg4IN_225, F(0)=>
      ImgReg4IN_224);
   loop3_14_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(239), 
      D(14)=>DATA(238), D(13)=>DATA(237), D(12)=>DATA(236), D(11)=>DATA(235), 
      D(10)=>DATA(234), D(9)=>DATA(233), D(8)=>DATA(232), D(7)=>DATA(231), 
      D(6)=>DATA(230), D(5)=>DATA(229), D(4)=>DATA(228), D(3)=>DATA(227), 
      D(2)=>DATA(226), D(1)=>DATA(225), D(0)=>DATA(224), EN=>nx23598, F(15)
      =>ImgReg5IN_239, F(14)=>ImgReg5IN_238, F(13)=>ImgReg5IN_237, F(12)=>
      ImgReg5IN_236, F(11)=>ImgReg5IN_235, F(10)=>ImgReg5IN_234, F(9)=>
      ImgReg5IN_233, F(8)=>ImgReg5IN_232, F(7)=>ImgReg5IN_231, F(6)=>
      ImgReg5IN_230, F(5)=>ImgReg5IN_229, F(4)=>ImgReg5IN_228, F(3)=>
      ImgReg5IN_227, F(2)=>ImgReg5IN_226, F(1)=>ImgReg5IN_225, F(0)=>
      ImgReg5IN_224);
   loop3_14_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_239_EXMPLR, D(14)=>OutputImg1_238_EXMPLR, D(13)=>
      OutputImg1_237_EXMPLR, D(12)=>OutputImg1_236_EXMPLR, D(11)=>
      OutputImg1_235_EXMPLR, D(10)=>OutputImg1_234_EXMPLR, D(9)=>
      OutputImg1_233_EXMPLR, D(8)=>OutputImg1_232_EXMPLR, D(7)=>
      OutputImg1_231_EXMPLR, D(6)=>OutputImg1_230_EXMPLR, D(5)=>
      OutputImg1_229_EXMPLR, D(4)=>OutputImg1_228_EXMPLR, D(3)=>
      OutputImg1_227_EXMPLR, D(2)=>OutputImg1_226_EXMPLR, D(1)=>
      OutputImg1_225_EXMPLR, D(0)=>OutputImg1_224_EXMPLR, EN=>nx23806, F(15)
      =>ImgReg0IN_239, F(14)=>ImgReg0IN_238, F(13)=>ImgReg0IN_237, F(12)=>
      ImgReg0IN_236, F(11)=>ImgReg0IN_235, F(10)=>ImgReg0IN_234, F(9)=>
      ImgReg0IN_233, F(8)=>ImgReg0IN_232, F(7)=>ImgReg0IN_231, F(6)=>
      ImgReg0IN_230, F(5)=>ImgReg0IN_229, F(4)=>ImgReg0IN_228, F(3)=>
      ImgReg0IN_227, F(2)=>ImgReg0IN_226, F(1)=>ImgReg0IN_225, F(0)=>
      ImgReg0IN_224);
   loop3_14_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_239_EXMPLR, D(14)=>OutputImg2_238_EXMPLR, D(13)=>
      OutputImg2_237_EXMPLR, D(12)=>OutputImg2_236_EXMPLR, D(11)=>
      OutputImg2_235_EXMPLR, D(10)=>OutputImg2_234_EXMPLR, D(9)=>
      OutputImg2_233_EXMPLR, D(8)=>OutputImg2_232_EXMPLR, D(7)=>
      OutputImg2_231_EXMPLR, D(6)=>OutputImg2_230_EXMPLR, D(5)=>
      OutputImg2_229_EXMPLR, D(4)=>OutputImg2_228_EXMPLR, D(3)=>
      OutputImg2_227_EXMPLR, D(2)=>OutputImg2_226_EXMPLR, D(1)=>
      OutputImg2_225_EXMPLR, D(0)=>OutputImg2_224_EXMPLR, EN=>nx23806, F(15)
      =>ImgReg1IN_239, F(14)=>ImgReg1IN_238, F(13)=>ImgReg1IN_237, F(12)=>
      ImgReg1IN_236, F(11)=>ImgReg1IN_235, F(10)=>ImgReg1IN_234, F(9)=>
      ImgReg1IN_233, F(8)=>ImgReg1IN_232, F(7)=>ImgReg1IN_231, F(6)=>
      ImgReg1IN_230, F(5)=>ImgReg1IN_229, F(4)=>ImgReg1IN_228, F(3)=>
      ImgReg1IN_227, F(2)=>ImgReg1IN_226, F(1)=>ImgReg1IN_225, F(0)=>
      ImgReg1IN_224);
   loop3_14_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_239_EXMPLR, D(14)=>OutputImg3_238_EXMPLR, D(13)=>
      OutputImg3_237_EXMPLR, D(12)=>OutputImg3_236_EXMPLR, D(11)=>
      OutputImg3_235_EXMPLR, D(10)=>OutputImg3_234_EXMPLR, D(9)=>
      OutputImg3_233_EXMPLR, D(8)=>OutputImg3_232_EXMPLR, D(7)=>
      OutputImg3_231_EXMPLR, D(6)=>OutputImg3_230_EXMPLR, D(5)=>
      OutputImg3_229_EXMPLR, D(4)=>OutputImg3_228_EXMPLR, D(3)=>
      OutputImg3_227_EXMPLR, D(2)=>OutputImg3_226_EXMPLR, D(1)=>
      OutputImg3_225_EXMPLR, D(0)=>OutputImg3_224_EXMPLR, EN=>nx23806, F(15)
      =>ImgReg2IN_239, F(14)=>ImgReg2IN_238, F(13)=>ImgReg2IN_237, F(12)=>
      ImgReg2IN_236, F(11)=>ImgReg2IN_235, F(10)=>ImgReg2IN_234, F(9)=>
      ImgReg2IN_233, F(8)=>ImgReg2IN_232, F(7)=>ImgReg2IN_231, F(6)=>
      ImgReg2IN_230, F(5)=>ImgReg2IN_229, F(4)=>ImgReg2IN_228, F(3)=>
      ImgReg2IN_227, F(2)=>ImgReg2IN_226, F(1)=>ImgReg2IN_225, F(0)=>
      ImgReg2IN_224);
   loop3_14_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_239_EXMPLR, D(14)=>OutputImg4_238_EXMPLR, D(13)=>
      OutputImg4_237_EXMPLR, D(12)=>OutputImg4_236_EXMPLR, D(11)=>
      OutputImg4_235_EXMPLR, D(10)=>OutputImg4_234_EXMPLR, D(9)=>
      OutputImg4_233_EXMPLR, D(8)=>OutputImg4_232_EXMPLR, D(7)=>
      OutputImg4_231_EXMPLR, D(6)=>OutputImg4_230_EXMPLR, D(5)=>
      OutputImg4_229_EXMPLR, D(4)=>OutputImg4_228_EXMPLR, D(3)=>
      OutputImg4_227_EXMPLR, D(2)=>OutputImg4_226_EXMPLR, D(1)=>
      OutputImg4_225_EXMPLR, D(0)=>OutputImg4_224_EXMPLR, EN=>nx23806, F(15)
      =>ImgReg3IN_239, F(14)=>ImgReg3IN_238, F(13)=>ImgReg3IN_237, F(12)=>
      ImgReg3IN_236, F(11)=>ImgReg3IN_235, F(10)=>ImgReg3IN_234, F(9)=>
      ImgReg3IN_233, F(8)=>ImgReg3IN_232, F(7)=>ImgReg3IN_231, F(6)=>
      ImgReg3IN_230, F(5)=>ImgReg3IN_229, F(4)=>ImgReg3IN_228, F(3)=>
      ImgReg3IN_227, F(2)=>ImgReg3IN_226, F(1)=>ImgReg3IN_225, F(0)=>
      ImgReg3IN_224);
   loop3_14_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_239_EXMPLR, D(14)=>OutputImg5_238_EXMPLR, D(13)=>
      OutputImg5_237_EXMPLR, D(12)=>OutputImg5_236_EXMPLR, D(11)=>
      OutputImg5_235_EXMPLR, D(10)=>OutputImg5_234_EXMPLR, D(9)=>
      OutputImg5_233_EXMPLR, D(8)=>OutputImg5_232_EXMPLR, D(7)=>
      OutputImg5_231_EXMPLR, D(6)=>OutputImg5_230_EXMPLR, D(5)=>
      OutputImg5_229_EXMPLR, D(4)=>OutputImg5_228_EXMPLR, D(3)=>
      OutputImg5_227_EXMPLR, D(2)=>OutputImg5_226_EXMPLR, D(1)=>
      OutputImg5_225_EXMPLR, D(0)=>OutputImg5_224_EXMPLR, EN=>nx23806, F(15)
      =>ImgReg4IN_239, F(14)=>ImgReg4IN_238, F(13)=>ImgReg4IN_237, F(12)=>
      ImgReg4IN_236, F(11)=>ImgReg4IN_235, F(10)=>ImgReg4IN_234, F(9)=>
      ImgReg4IN_233, F(8)=>ImgReg4IN_232, F(7)=>ImgReg4IN_231, F(6)=>
      ImgReg4IN_230, F(5)=>ImgReg4IN_229, F(4)=>ImgReg4IN_228, F(3)=>
      ImgReg4IN_227, F(2)=>ImgReg4IN_226, F(1)=>ImgReg4IN_225, F(0)=>
      ImgReg4IN_224);
   loop3_14_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_239, D(14)=>
      ImgReg0IN_238, D(13)=>ImgReg0IN_237, D(12)=>ImgReg0IN_236, D(11)=>
      ImgReg0IN_235, D(10)=>ImgReg0IN_234, D(9)=>ImgReg0IN_233, D(8)=>
      ImgReg0IN_232, D(7)=>ImgReg0IN_231, D(6)=>ImgReg0IN_230, D(5)=>
      ImgReg0IN_229, D(4)=>ImgReg0IN_228, D(3)=>ImgReg0IN_227, D(2)=>
      ImgReg0IN_226, D(1)=>ImgReg0IN_225, D(0)=>ImgReg0IN_224, CLK=>nx23912, 
      RST=>RST, EN=>nx23722, Q(15)=>OutputImg0_239_EXMPLR, Q(14)=>
      OutputImg0_238_EXMPLR, Q(13)=>OutputImg0_237_EXMPLR, Q(12)=>
      OutputImg0_236_EXMPLR, Q(11)=>OutputImg0_235_EXMPLR, Q(10)=>
      OutputImg0_234_EXMPLR, Q(9)=>OutputImg0_233_EXMPLR, Q(8)=>
      OutputImg0_232_EXMPLR, Q(7)=>OutputImg0_231_EXMPLR, Q(6)=>
      OutputImg0_230_EXMPLR, Q(5)=>OutputImg0_229_EXMPLR, Q(4)=>
      OutputImg0_228_EXMPLR, Q(3)=>OutputImg0_227_EXMPLR, Q(2)=>
      OutputImg0_226_EXMPLR, Q(1)=>OutputImg0_225_EXMPLR, Q(0)=>
      OutputImg0_224_EXMPLR);
   loop3_14_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_239, D(14)=>
      ImgReg1IN_238, D(13)=>ImgReg1IN_237, D(12)=>ImgReg1IN_236, D(11)=>
      ImgReg1IN_235, D(10)=>ImgReg1IN_234, D(9)=>ImgReg1IN_233, D(8)=>
      ImgReg1IN_232, D(7)=>ImgReg1IN_231, D(6)=>ImgReg1IN_230, D(5)=>
      ImgReg1IN_229, D(4)=>ImgReg1IN_228, D(3)=>ImgReg1IN_227, D(2)=>
      ImgReg1IN_226, D(1)=>ImgReg1IN_225, D(0)=>ImgReg1IN_224, CLK=>nx23914, 
      RST=>RST, EN=>nx23732, Q(15)=>OutputImg1_239_EXMPLR, Q(14)=>
      OutputImg1_238_EXMPLR, Q(13)=>OutputImg1_237_EXMPLR, Q(12)=>
      OutputImg1_236_EXMPLR, Q(11)=>OutputImg1_235_EXMPLR, Q(10)=>
      OutputImg1_234_EXMPLR, Q(9)=>OutputImg1_233_EXMPLR, Q(8)=>
      OutputImg1_232_EXMPLR, Q(7)=>OutputImg1_231_EXMPLR, Q(6)=>
      OutputImg1_230_EXMPLR, Q(5)=>OutputImg1_229_EXMPLR, Q(4)=>
      OutputImg1_228_EXMPLR, Q(3)=>OutputImg1_227_EXMPLR, Q(2)=>
      OutputImg1_226_EXMPLR, Q(1)=>OutputImg1_225_EXMPLR, Q(0)=>
      OutputImg1_224_EXMPLR);
   loop3_14_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_239, D(14)=>
      ImgReg2IN_238, D(13)=>ImgReg2IN_237, D(12)=>ImgReg2IN_236, D(11)=>
      ImgReg2IN_235, D(10)=>ImgReg2IN_234, D(9)=>ImgReg2IN_233, D(8)=>
      ImgReg2IN_232, D(7)=>ImgReg2IN_231, D(6)=>ImgReg2IN_230, D(5)=>
      ImgReg2IN_229, D(4)=>ImgReg2IN_228, D(3)=>ImgReg2IN_227, D(2)=>
      ImgReg2IN_226, D(1)=>ImgReg2IN_225, D(0)=>ImgReg2IN_224, CLK=>nx23914, 
      RST=>RST, EN=>nx23742, Q(15)=>OutputImg2_239_EXMPLR, Q(14)=>
      OutputImg2_238_EXMPLR, Q(13)=>OutputImg2_237_EXMPLR, Q(12)=>
      OutputImg2_236_EXMPLR, Q(11)=>OutputImg2_235_EXMPLR, Q(10)=>
      OutputImg2_234_EXMPLR, Q(9)=>OutputImg2_233_EXMPLR, Q(8)=>
      OutputImg2_232_EXMPLR, Q(7)=>OutputImg2_231_EXMPLR, Q(6)=>
      OutputImg2_230_EXMPLR, Q(5)=>OutputImg2_229_EXMPLR, Q(4)=>
      OutputImg2_228_EXMPLR, Q(3)=>OutputImg2_227_EXMPLR, Q(2)=>
      OutputImg2_226_EXMPLR, Q(1)=>OutputImg2_225_EXMPLR, Q(0)=>
      OutputImg2_224_EXMPLR);
   loop3_14_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_239, D(14)=>
      ImgReg3IN_238, D(13)=>ImgReg3IN_237, D(12)=>ImgReg3IN_236, D(11)=>
      ImgReg3IN_235, D(10)=>ImgReg3IN_234, D(9)=>ImgReg3IN_233, D(8)=>
      ImgReg3IN_232, D(7)=>ImgReg3IN_231, D(6)=>ImgReg3IN_230, D(5)=>
      ImgReg3IN_229, D(4)=>ImgReg3IN_228, D(3)=>ImgReg3IN_227, D(2)=>
      ImgReg3IN_226, D(1)=>ImgReg3IN_225, D(0)=>ImgReg3IN_224, CLK=>nx23916, 
      RST=>RST, EN=>nx23752, Q(15)=>OutputImg3_239_EXMPLR, Q(14)=>
      OutputImg3_238_EXMPLR, Q(13)=>OutputImg3_237_EXMPLR, Q(12)=>
      OutputImg3_236_EXMPLR, Q(11)=>OutputImg3_235_EXMPLR, Q(10)=>
      OutputImg3_234_EXMPLR, Q(9)=>OutputImg3_233_EXMPLR, Q(8)=>
      OutputImg3_232_EXMPLR, Q(7)=>OutputImg3_231_EXMPLR, Q(6)=>
      OutputImg3_230_EXMPLR, Q(5)=>OutputImg3_229_EXMPLR, Q(4)=>
      OutputImg3_228_EXMPLR, Q(3)=>OutputImg3_227_EXMPLR, Q(2)=>
      OutputImg3_226_EXMPLR, Q(1)=>OutputImg3_225_EXMPLR, Q(0)=>
      OutputImg3_224_EXMPLR);
   loop3_14_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_239, D(14)=>
      ImgReg4IN_238, D(13)=>ImgReg4IN_237, D(12)=>ImgReg4IN_236, D(11)=>
      ImgReg4IN_235, D(10)=>ImgReg4IN_234, D(9)=>ImgReg4IN_233, D(8)=>
      ImgReg4IN_232, D(7)=>ImgReg4IN_231, D(6)=>ImgReg4IN_230, D(5)=>
      ImgReg4IN_229, D(4)=>ImgReg4IN_228, D(3)=>ImgReg4IN_227, D(2)=>
      ImgReg4IN_226, D(1)=>ImgReg4IN_225, D(0)=>ImgReg4IN_224, CLK=>nx23916, 
      RST=>RST, EN=>nx23762, Q(15)=>OutputImg4_239_EXMPLR, Q(14)=>
      OutputImg4_238_EXMPLR, Q(13)=>OutputImg4_237_EXMPLR, Q(12)=>
      OutputImg4_236_EXMPLR, Q(11)=>OutputImg4_235_EXMPLR, Q(10)=>
      OutputImg4_234_EXMPLR, Q(9)=>OutputImg4_233_EXMPLR, Q(8)=>
      OutputImg4_232_EXMPLR, Q(7)=>OutputImg4_231_EXMPLR, Q(6)=>
      OutputImg4_230_EXMPLR, Q(5)=>OutputImg4_229_EXMPLR, Q(4)=>
      OutputImg4_228_EXMPLR, Q(3)=>OutputImg4_227_EXMPLR, Q(2)=>
      OutputImg4_226_EXMPLR, Q(1)=>OutputImg4_225_EXMPLR, Q(0)=>
      OutputImg4_224_EXMPLR);
   loop3_14_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_239, D(14)=>
      ImgReg5IN_238, D(13)=>ImgReg5IN_237, D(12)=>ImgReg5IN_236, D(11)=>
      ImgReg5IN_235, D(10)=>ImgReg5IN_234, D(9)=>ImgReg5IN_233, D(8)=>
      ImgReg5IN_232, D(7)=>ImgReg5IN_231, D(6)=>ImgReg5IN_230, D(5)=>
      ImgReg5IN_229, D(4)=>ImgReg5IN_228, D(3)=>ImgReg5IN_227, D(2)=>
      ImgReg5IN_226, D(1)=>ImgReg5IN_225, D(0)=>ImgReg5IN_224, CLK=>nx23918, 
      RST=>RST, EN=>nx23772, Q(15)=>OutputImg5_239_EXMPLR, Q(14)=>
      OutputImg5_238_EXMPLR, Q(13)=>OutputImg5_237_EXMPLR, Q(12)=>
      OutputImg5_236_EXMPLR, Q(11)=>OutputImg5_235_EXMPLR, Q(10)=>
      OutputImg5_234_EXMPLR, Q(9)=>OutputImg5_233_EXMPLR, Q(8)=>
      OutputImg5_232_EXMPLR, Q(7)=>OutputImg5_231_EXMPLR, Q(6)=>
      OutputImg5_230_EXMPLR, Q(5)=>OutputImg5_229_EXMPLR, Q(4)=>
      OutputImg5_228_EXMPLR, Q(3)=>OutputImg5_227_EXMPLR, Q(2)=>
      OutputImg5_226_EXMPLR, Q(1)=>OutputImg5_225_EXMPLR, Q(0)=>
      OutputImg5_224_EXMPLR);
   loop3_15_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_271_EXMPLR, D(14)=>OutputImg0_270_EXMPLR, D(13)=>
      OutputImg0_269_EXMPLR, D(12)=>OutputImg0_268_EXMPLR, D(11)=>
      OutputImg0_267_EXMPLR, D(10)=>OutputImg0_266_EXMPLR, D(9)=>
      OutputImg0_265_EXMPLR, D(8)=>OutputImg0_264_EXMPLR, D(7)=>
      OutputImg0_263_EXMPLR, D(6)=>OutputImg0_262_EXMPLR, D(5)=>
      OutputImg0_261_EXMPLR, D(4)=>OutputImg0_260_EXMPLR, D(3)=>
      OutputImg0_259_EXMPLR, D(2)=>OutputImg0_258_EXMPLR, D(1)=>
      OutputImg0_257_EXMPLR, D(0)=>OutputImg0_256_EXMPLR, EN=>nx23690, F(15)
      =>ImgReg0IN_255, F(14)=>ImgReg0IN_254, F(13)=>ImgReg0IN_253, F(12)=>
      ImgReg0IN_252, F(11)=>ImgReg0IN_251, F(10)=>ImgReg0IN_250, F(9)=>
      ImgReg0IN_249, F(8)=>ImgReg0IN_248, F(7)=>ImgReg0IN_247, F(6)=>
      ImgReg0IN_246, F(5)=>ImgReg0IN_245, F(4)=>ImgReg0IN_244, F(3)=>
      ImgReg0IN_243, F(2)=>ImgReg0IN_242, F(1)=>ImgReg0IN_241, F(0)=>
      ImgReg0IN_240);
   loop3_15_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_271_EXMPLR, D(14)=>OutputImg1_270_EXMPLR, D(13)=>
      OutputImg1_269_EXMPLR, D(12)=>OutputImg1_268_EXMPLR, D(11)=>
      OutputImg1_267_EXMPLR, D(10)=>OutputImg1_266_EXMPLR, D(9)=>
      OutputImg1_265_EXMPLR, D(8)=>OutputImg1_264_EXMPLR, D(7)=>
      OutputImg1_263_EXMPLR, D(6)=>OutputImg1_262_EXMPLR, D(5)=>
      OutputImg1_261_EXMPLR, D(4)=>OutputImg1_260_EXMPLR, D(3)=>
      OutputImg1_259_EXMPLR, D(2)=>OutputImg1_258_EXMPLR, D(1)=>
      OutputImg1_257_EXMPLR, D(0)=>OutputImg1_256_EXMPLR, EN=>nx23692, F(15)
      =>ImgReg1IN_255, F(14)=>ImgReg1IN_254, F(13)=>ImgReg1IN_253, F(12)=>
      ImgReg1IN_252, F(11)=>ImgReg1IN_251, F(10)=>ImgReg1IN_250, F(9)=>
      ImgReg1IN_249, F(8)=>ImgReg1IN_248, F(7)=>ImgReg1IN_247, F(6)=>
      ImgReg1IN_246, F(5)=>ImgReg1IN_245, F(4)=>ImgReg1IN_244, F(3)=>
      ImgReg1IN_243, F(2)=>ImgReg1IN_242, F(1)=>ImgReg1IN_241, F(0)=>
      ImgReg1IN_240);
   loop3_15_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_271_EXMPLR, D(14)=>OutputImg2_270_EXMPLR, D(13)=>
      OutputImg2_269_EXMPLR, D(12)=>OutputImg2_268_EXMPLR, D(11)=>
      OutputImg2_267_EXMPLR, D(10)=>OutputImg2_266_EXMPLR, D(9)=>
      OutputImg2_265_EXMPLR, D(8)=>OutputImg2_264_EXMPLR, D(7)=>
      OutputImg2_263_EXMPLR, D(6)=>OutputImg2_262_EXMPLR, D(5)=>
      OutputImg2_261_EXMPLR, D(4)=>OutputImg2_260_EXMPLR, D(3)=>
      OutputImg2_259_EXMPLR, D(2)=>OutputImg2_258_EXMPLR, D(1)=>
      OutputImg2_257_EXMPLR, D(0)=>OutputImg2_256_EXMPLR, EN=>nx23692, F(15)
      =>ImgReg2IN_255, F(14)=>ImgReg2IN_254, F(13)=>ImgReg2IN_253, F(12)=>
      ImgReg2IN_252, F(11)=>ImgReg2IN_251, F(10)=>ImgReg2IN_250, F(9)=>
      ImgReg2IN_249, F(8)=>ImgReg2IN_248, F(7)=>ImgReg2IN_247, F(6)=>
      ImgReg2IN_246, F(5)=>ImgReg2IN_245, F(4)=>ImgReg2IN_244, F(3)=>
      ImgReg2IN_243, F(2)=>ImgReg2IN_242, F(1)=>ImgReg2IN_241, F(0)=>
      ImgReg2IN_240);
   loop3_15_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_271_EXMPLR, D(14)=>OutputImg3_270_EXMPLR, D(13)=>
      OutputImg3_269_EXMPLR, D(12)=>OutputImg3_268_EXMPLR, D(11)=>
      OutputImg3_267_EXMPLR, D(10)=>OutputImg3_266_EXMPLR, D(9)=>
      OutputImg3_265_EXMPLR, D(8)=>OutputImg3_264_EXMPLR, D(7)=>
      OutputImg3_263_EXMPLR, D(6)=>OutputImg3_262_EXMPLR, D(5)=>
      OutputImg3_261_EXMPLR, D(4)=>OutputImg3_260_EXMPLR, D(3)=>
      OutputImg3_259_EXMPLR, D(2)=>OutputImg3_258_EXMPLR, D(1)=>
      OutputImg3_257_EXMPLR, D(0)=>OutputImg3_256_EXMPLR, EN=>nx23692, F(15)
      =>ImgReg3IN_255, F(14)=>ImgReg3IN_254, F(13)=>ImgReg3IN_253, F(12)=>
      ImgReg3IN_252, F(11)=>ImgReg3IN_251, F(10)=>ImgReg3IN_250, F(9)=>
      ImgReg3IN_249, F(8)=>ImgReg3IN_248, F(7)=>ImgReg3IN_247, F(6)=>
      ImgReg3IN_246, F(5)=>ImgReg3IN_245, F(4)=>ImgReg3IN_244, F(3)=>
      ImgReg3IN_243, F(2)=>ImgReg3IN_242, F(1)=>ImgReg3IN_241, F(0)=>
      ImgReg3IN_240);
   loop3_15_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_271_EXMPLR, D(14)=>OutputImg4_270_EXMPLR, D(13)=>
      OutputImg4_269_EXMPLR, D(12)=>OutputImg4_268_EXMPLR, D(11)=>
      OutputImg4_267_EXMPLR, D(10)=>OutputImg4_266_EXMPLR, D(9)=>
      OutputImg4_265_EXMPLR, D(8)=>OutputImg4_264_EXMPLR, D(7)=>
      OutputImg4_263_EXMPLR, D(6)=>OutputImg4_262_EXMPLR, D(5)=>
      OutputImg4_261_EXMPLR, D(4)=>OutputImg4_260_EXMPLR, D(3)=>
      OutputImg4_259_EXMPLR, D(2)=>OutputImg4_258_EXMPLR, D(1)=>
      OutputImg4_257_EXMPLR, D(0)=>OutputImg4_256_EXMPLR, EN=>nx23692, F(15)
      =>ImgReg4IN_255, F(14)=>ImgReg4IN_254, F(13)=>ImgReg4IN_253, F(12)=>
      ImgReg4IN_252, F(11)=>ImgReg4IN_251, F(10)=>ImgReg4IN_250, F(9)=>
      ImgReg4IN_249, F(8)=>ImgReg4IN_248, F(7)=>ImgReg4IN_247, F(6)=>
      ImgReg4IN_246, F(5)=>ImgReg4IN_245, F(4)=>ImgReg4IN_244, F(3)=>
      ImgReg4IN_243, F(2)=>ImgReg4IN_242, F(1)=>ImgReg4IN_241, F(0)=>
      ImgReg4IN_240);
   loop3_15_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_271_EXMPLR, D(14)=>OutputImg5_270_EXMPLR, D(13)=>
      OutputImg5_269_EXMPLR, D(12)=>OutputImg5_268_EXMPLR, D(11)=>
      OutputImg5_267_EXMPLR, D(10)=>OutputImg5_266_EXMPLR, D(9)=>
      OutputImg5_265_EXMPLR, D(8)=>OutputImg5_264_EXMPLR, D(7)=>
      OutputImg5_263_EXMPLR, D(6)=>OutputImg5_262_EXMPLR, D(5)=>
      OutputImg5_261_EXMPLR, D(4)=>OutputImg5_260_EXMPLR, D(3)=>
      OutputImg5_259_EXMPLR, D(2)=>OutputImg5_258_EXMPLR, D(1)=>
      OutputImg5_257_EXMPLR, D(0)=>OutputImg5_256_EXMPLR, EN=>nx23692, F(15)
      =>ImgReg5IN_255, F(14)=>ImgReg5IN_254, F(13)=>ImgReg5IN_253, F(12)=>
      ImgReg5IN_252, F(11)=>ImgReg5IN_251, F(10)=>ImgReg5IN_250, F(9)=>
      ImgReg5IN_249, F(8)=>ImgReg5IN_248, F(7)=>ImgReg5IN_247, F(6)=>
      ImgReg5IN_246, F(5)=>ImgReg5IN_245, F(4)=>ImgReg5IN_244, F(3)=>
      ImgReg5IN_243, F(2)=>ImgReg5IN_242, F(1)=>ImgReg5IN_241, F(0)=>
      ImgReg5IN_240);
   loop3_15_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(255), 
      D(14)=>DATA(254), D(13)=>DATA(253), D(12)=>DATA(252), D(11)=>DATA(251), 
      D(10)=>DATA(250), D(9)=>DATA(249), D(8)=>DATA(248), D(7)=>DATA(247), 
      D(6)=>DATA(246), D(5)=>DATA(245), D(4)=>DATA(244), D(3)=>DATA(243), 
      D(2)=>DATA(242), D(1)=>DATA(241), D(0)=>DATA(240), EN=>nx23658, F(15)
      =>ImgReg0IN_255, F(14)=>ImgReg0IN_254, F(13)=>ImgReg0IN_253, F(12)=>
      ImgReg0IN_252, F(11)=>ImgReg0IN_251, F(10)=>ImgReg0IN_250, F(9)=>
      ImgReg0IN_249, F(8)=>ImgReg0IN_248, F(7)=>ImgReg0IN_247, F(6)=>
      ImgReg0IN_246, F(5)=>ImgReg0IN_245, F(4)=>ImgReg0IN_244, F(3)=>
      ImgReg0IN_243, F(2)=>ImgReg0IN_242, F(1)=>ImgReg0IN_241, F(0)=>
      ImgReg0IN_240);
   loop3_15_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(255), 
      D(14)=>DATA(254), D(13)=>DATA(253), D(12)=>DATA(252), D(11)=>DATA(251), 
      D(10)=>DATA(250), D(9)=>DATA(249), D(8)=>DATA(248), D(7)=>DATA(247), 
      D(6)=>DATA(246), D(5)=>DATA(245), D(4)=>DATA(244), D(3)=>DATA(243), 
      D(2)=>DATA(242), D(1)=>DATA(241), D(0)=>DATA(240), EN=>nx23646, F(15)
      =>ImgReg1IN_255, F(14)=>ImgReg1IN_254, F(13)=>ImgReg1IN_253, F(12)=>
      ImgReg1IN_252, F(11)=>ImgReg1IN_251, F(10)=>ImgReg1IN_250, F(9)=>
      ImgReg1IN_249, F(8)=>ImgReg1IN_248, F(7)=>ImgReg1IN_247, F(6)=>
      ImgReg1IN_246, F(5)=>ImgReg1IN_245, F(4)=>ImgReg1IN_244, F(3)=>
      ImgReg1IN_243, F(2)=>ImgReg1IN_242, F(1)=>ImgReg1IN_241, F(0)=>
      ImgReg1IN_240);
   loop3_15_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(255), 
      D(14)=>DATA(254), D(13)=>DATA(253), D(12)=>DATA(252), D(11)=>DATA(251), 
      D(10)=>DATA(250), D(9)=>DATA(249), D(8)=>DATA(248), D(7)=>DATA(247), 
      D(6)=>DATA(246), D(5)=>DATA(245), D(4)=>DATA(244), D(3)=>DATA(243), 
      D(2)=>DATA(242), D(1)=>DATA(241), D(0)=>DATA(240), EN=>nx23634, F(15)
      =>ImgReg2IN_255, F(14)=>ImgReg2IN_254, F(13)=>ImgReg2IN_253, F(12)=>
      ImgReg2IN_252, F(11)=>ImgReg2IN_251, F(10)=>ImgReg2IN_250, F(9)=>
      ImgReg2IN_249, F(8)=>ImgReg2IN_248, F(7)=>ImgReg2IN_247, F(6)=>
      ImgReg2IN_246, F(5)=>ImgReg2IN_245, F(4)=>ImgReg2IN_244, F(3)=>
      ImgReg2IN_243, F(2)=>ImgReg2IN_242, F(1)=>ImgReg2IN_241, F(0)=>
      ImgReg2IN_240);
   loop3_15_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(255), 
      D(14)=>DATA(254), D(13)=>DATA(253), D(12)=>DATA(252), D(11)=>DATA(251), 
      D(10)=>DATA(250), D(9)=>DATA(249), D(8)=>DATA(248), D(7)=>DATA(247), 
      D(6)=>DATA(246), D(5)=>DATA(245), D(4)=>DATA(244), D(3)=>DATA(243), 
      D(2)=>DATA(242), D(1)=>DATA(241), D(0)=>DATA(240), EN=>nx23622, F(15)
      =>ImgReg3IN_255, F(14)=>ImgReg3IN_254, F(13)=>ImgReg3IN_253, F(12)=>
      ImgReg3IN_252, F(11)=>ImgReg3IN_251, F(10)=>ImgReg3IN_250, F(9)=>
      ImgReg3IN_249, F(8)=>ImgReg3IN_248, F(7)=>ImgReg3IN_247, F(6)=>
      ImgReg3IN_246, F(5)=>ImgReg3IN_245, F(4)=>ImgReg3IN_244, F(3)=>
      ImgReg3IN_243, F(2)=>ImgReg3IN_242, F(1)=>ImgReg3IN_241, F(0)=>
      ImgReg3IN_240);
   loop3_15_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(255), 
      D(14)=>DATA(254), D(13)=>DATA(253), D(12)=>DATA(252), D(11)=>DATA(251), 
      D(10)=>DATA(250), D(9)=>DATA(249), D(8)=>DATA(248), D(7)=>DATA(247), 
      D(6)=>DATA(246), D(5)=>DATA(245), D(4)=>DATA(244), D(3)=>DATA(243), 
      D(2)=>DATA(242), D(1)=>DATA(241), D(0)=>DATA(240), EN=>nx23610, F(15)
      =>ImgReg4IN_255, F(14)=>ImgReg4IN_254, F(13)=>ImgReg4IN_253, F(12)=>
      ImgReg4IN_252, F(11)=>ImgReg4IN_251, F(10)=>ImgReg4IN_250, F(9)=>
      ImgReg4IN_249, F(8)=>ImgReg4IN_248, F(7)=>ImgReg4IN_247, F(6)=>
      ImgReg4IN_246, F(5)=>ImgReg4IN_245, F(4)=>ImgReg4IN_244, F(3)=>
      ImgReg4IN_243, F(2)=>ImgReg4IN_242, F(1)=>ImgReg4IN_241, F(0)=>
      ImgReg4IN_240);
   loop3_15_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(255), 
      D(14)=>DATA(254), D(13)=>DATA(253), D(12)=>DATA(252), D(11)=>DATA(251), 
      D(10)=>DATA(250), D(9)=>DATA(249), D(8)=>DATA(248), D(7)=>DATA(247), 
      D(6)=>DATA(246), D(5)=>DATA(245), D(4)=>DATA(244), D(3)=>DATA(243), 
      D(2)=>DATA(242), D(1)=>DATA(241), D(0)=>DATA(240), EN=>nx23598, F(15)
      =>ImgReg5IN_255, F(14)=>ImgReg5IN_254, F(13)=>ImgReg5IN_253, F(12)=>
      ImgReg5IN_252, F(11)=>ImgReg5IN_251, F(10)=>ImgReg5IN_250, F(9)=>
      ImgReg5IN_249, F(8)=>ImgReg5IN_248, F(7)=>ImgReg5IN_247, F(6)=>
      ImgReg5IN_246, F(5)=>ImgReg5IN_245, F(4)=>ImgReg5IN_244, F(3)=>
      ImgReg5IN_243, F(2)=>ImgReg5IN_242, F(1)=>ImgReg5IN_241, F(0)=>
      ImgReg5IN_240);
   loop3_15_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_255_EXMPLR, D(14)=>OutputImg1_254_EXMPLR, D(13)=>
      OutputImg1_253_EXMPLR, D(12)=>OutputImg1_252_EXMPLR, D(11)=>
      OutputImg1_251_EXMPLR, D(10)=>OutputImg1_250_EXMPLR, D(9)=>
      OutputImg1_249_EXMPLR, D(8)=>OutputImg1_248_EXMPLR, D(7)=>
      OutputImg1_247_EXMPLR, D(6)=>OutputImg1_246_EXMPLR, D(5)=>
      OutputImg1_245_EXMPLR, D(4)=>OutputImg1_244_EXMPLR, D(3)=>
      OutputImg1_243_EXMPLR, D(2)=>OutputImg1_242_EXMPLR, D(1)=>
      OutputImg1_241_EXMPLR, D(0)=>OutputImg1_240_EXMPLR, EN=>nx23806, F(15)
      =>ImgReg0IN_255, F(14)=>ImgReg0IN_254, F(13)=>ImgReg0IN_253, F(12)=>
      ImgReg0IN_252, F(11)=>ImgReg0IN_251, F(10)=>ImgReg0IN_250, F(9)=>
      ImgReg0IN_249, F(8)=>ImgReg0IN_248, F(7)=>ImgReg0IN_247, F(6)=>
      ImgReg0IN_246, F(5)=>ImgReg0IN_245, F(4)=>ImgReg0IN_244, F(3)=>
      ImgReg0IN_243, F(2)=>ImgReg0IN_242, F(1)=>ImgReg0IN_241, F(0)=>
      ImgReg0IN_240);
   loop3_15_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_255_EXMPLR, D(14)=>OutputImg2_254_EXMPLR, D(13)=>
      OutputImg2_253_EXMPLR, D(12)=>OutputImg2_252_EXMPLR, D(11)=>
      OutputImg2_251_EXMPLR, D(10)=>OutputImg2_250_EXMPLR, D(9)=>
      OutputImg2_249_EXMPLR, D(8)=>OutputImg2_248_EXMPLR, D(7)=>
      OutputImg2_247_EXMPLR, D(6)=>OutputImg2_246_EXMPLR, D(5)=>
      OutputImg2_245_EXMPLR, D(4)=>OutputImg2_244_EXMPLR, D(3)=>
      OutputImg2_243_EXMPLR, D(2)=>OutputImg2_242_EXMPLR, D(1)=>
      OutputImg2_241_EXMPLR, D(0)=>OutputImg2_240_EXMPLR, EN=>nx23806, F(15)
      =>ImgReg1IN_255, F(14)=>ImgReg1IN_254, F(13)=>ImgReg1IN_253, F(12)=>
      ImgReg1IN_252, F(11)=>ImgReg1IN_251, F(10)=>ImgReg1IN_250, F(9)=>
      ImgReg1IN_249, F(8)=>ImgReg1IN_248, F(7)=>ImgReg1IN_247, F(6)=>
      ImgReg1IN_246, F(5)=>ImgReg1IN_245, F(4)=>ImgReg1IN_244, F(3)=>
      ImgReg1IN_243, F(2)=>ImgReg1IN_242, F(1)=>ImgReg1IN_241, F(0)=>
      ImgReg1IN_240);
   loop3_15_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_255_EXMPLR, D(14)=>OutputImg3_254_EXMPLR, D(13)=>
      OutputImg3_253_EXMPLR, D(12)=>OutputImg3_252_EXMPLR, D(11)=>
      OutputImg3_251_EXMPLR, D(10)=>OutputImg3_250_EXMPLR, D(9)=>
      OutputImg3_249_EXMPLR, D(8)=>OutputImg3_248_EXMPLR, D(7)=>
      OutputImg3_247_EXMPLR, D(6)=>OutputImg3_246_EXMPLR, D(5)=>
      OutputImg3_245_EXMPLR, D(4)=>OutputImg3_244_EXMPLR, D(3)=>
      OutputImg3_243_EXMPLR, D(2)=>OutputImg3_242_EXMPLR, D(1)=>
      OutputImg3_241_EXMPLR, D(0)=>OutputImg3_240_EXMPLR, EN=>nx23808, F(15)
      =>ImgReg2IN_255, F(14)=>ImgReg2IN_254, F(13)=>ImgReg2IN_253, F(12)=>
      ImgReg2IN_252, F(11)=>ImgReg2IN_251, F(10)=>ImgReg2IN_250, F(9)=>
      ImgReg2IN_249, F(8)=>ImgReg2IN_248, F(7)=>ImgReg2IN_247, F(6)=>
      ImgReg2IN_246, F(5)=>ImgReg2IN_245, F(4)=>ImgReg2IN_244, F(3)=>
      ImgReg2IN_243, F(2)=>ImgReg2IN_242, F(1)=>ImgReg2IN_241, F(0)=>
      ImgReg2IN_240);
   loop3_15_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_255_EXMPLR, D(14)=>OutputImg4_254_EXMPLR, D(13)=>
      OutputImg4_253_EXMPLR, D(12)=>OutputImg4_252_EXMPLR, D(11)=>
      OutputImg4_251_EXMPLR, D(10)=>OutputImg4_250_EXMPLR, D(9)=>
      OutputImg4_249_EXMPLR, D(8)=>OutputImg4_248_EXMPLR, D(7)=>
      OutputImg4_247_EXMPLR, D(6)=>OutputImg4_246_EXMPLR, D(5)=>
      OutputImg4_245_EXMPLR, D(4)=>OutputImg4_244_EXMPLR, D(3)=>
      OutputImg4_243_EXMPLR, D(2)=>OutputImg4_242_EXMPLR, D(1)=>
      OutputImg4_241_EXMPLR, D(0)=>OutputImg4_240_EXMPLR, EN=>nx23808, F(15)
      =>ImgReg3IN_255, F(14)=>ImgReg3IN_254, F(13)=>ImgReg3IN_253, F(12)=>
      ImgReg3IN_252, F(11)=>ImgReg3IN_251, F(10)=>ImgReg3IN_250, F(9)=>
      ImgReg3IN_249, F(8)=>ImgReg3IN_248, F(7)=>ImgReg3IN_247, F(6)=>
      ImgReg3IN_246, F(5)=>ImgReg3IN_245, F(4)=>ImgReg3IN_244, F(3)=>
      ImgReg3IN_243, F(2)=>ImgReg3IN_242, F(1)=>ImgReg3IN_241, F(0)=>
      ImgReg3IN_240);
   loop3_15_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_255_EXMPLR, D(14)=>OutputImg5_254_EXMPLR, D(13)=>
      OutputImg5_253_EXMPLR, D(12)=>OutputImg5_252_EXMPLR, D(11)=>
      OutputImg5_251_EXMPLR, D(10)=>OutputImg5_250_EXMPLR, D(9)=>
      OutputImg5_249_EXMPLR, D(8)=>OutputImg5_248_EXMPLR, D(7)=>
      OutputImg5_247_EXMPLR, D(6)=>OutputImg5_246_EXMPLR, D(5)=>
      OutputImg5_245_EXMPLR, D(4)=>OutputImg5_244_EXMPLR, D(3)=>
      OutputImg5_243_EXMPLR, D(2)=>OutputImg5_242_EXMPLR, D(1)=>
      OutputImg5_241_EXMPLR, D(0)=>OutputImg5_240_EXMPLR, EN=>nx23808, F(15)
      =>ImgReg4IN_255, F(14)=>ImgReg4IN_254, F(13)=>ImgReg4IN_253, F(12)=>
      ImgReg4IN_252, F(11)=>ImgReg4IN_251, F(10)=>ImgReg4IN_250, F(9)=>
      ImgReg4IN_249, F(8)=>ImgReg4IN_248, F(7)=>ImgReg4IN_247, F(6)=>
      ImgReg4IN_246, F(5)=>ImgReg4IN_245, F(4)=>ImgReg4IN_244, F(3)=>
      ImgReg4IN_243, F(2)=>ImgReg4IN_242, F(1)=>ImgReg4IN_241, F(0)=>
      ImgReg4IN_240);
   loop3_15_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_255, D(14)=>
      ImgReg0IN_254, D(13)=>ImgReg0IN_253, D(12)=>ImgReg0IN_252, D(11)=>
      ImgReg0IN_251, D(10)=>ImgReg0IN_250, D(9)=>ImgReg0IN_249, D(8)=>
      ImgReg0IN_248, D(7)=>ImgReg0IN_247, D(6)=>ImgReg0IN_246, D(5)=>
      ImgReg0IN_245, D(4)=>ImgReg0IN_244, D(3)=>ImgReg0IN_243, D(2)=>
      ImgReg0IN_242, D(1)=>ImgReg0IN_241, D(0)=>ImgReg0IN_240, CLK=>nx23918, 
      RST=>RST, EN=>nx23722, Q(15)=>OutputImg0_255_EXMPLR, Q(14)=>
      OutputImg0_254_EXMPLR, Q(13)=>OutputImg0_253_EXMPLR, Q(12)=>
      OutputImg0_252_EXMPLR, Q(11)=>OutputImg0_251_EXMPLR, Q(10)=>
      OutputImg0_250_EXMPLR, Q(9)=>OutputImg0_249_EXMPLR, Q(8)=>
      OutputImg0_248_EXMPLR, Q(7)=>OutputImg0_247_EXMPLR, Q(6)=>
      OutputImg0_246_EXMPLR, Q(5)=>OutputImg0_245_EXMPLR, Q(4)=>
      OutputImg0_244_EXMPLR, Q(3)=>OutputImg0_243_EXMPLR, Q(2)=>
      OutputImg0_242_EXMPLR, Q(1)=>OutputImg0_241_EXMPLR, Q(0)=>
      OutputImg0_240_EXMPLR);
   loop3_15_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_255, D(14)=>
      ImgReg1IN_254, D(13)=>ImgReg1IN_253, D(12)=>ImgReg1IN_252, D(11)=>
      ImgReg1IN_251, D(10)=>ImgReg1IN_250, D(9)=>ImgReg1IN_249, D(8)=>
      ImgReg1IN_248, D(7)=>ImgReg1IN_247, D(6)=>ImgReg1IN_246, D(5)=>
      ImgReg1IN_245, D(4)=>ImgReg1IN_244, D(3)=>ImgReg1IN_243, D(2)=>
      ImgReg1IN_242, D(1)=>ImgReg1IN_241, D(0)=>ImgReg1IN_240, CLK=>nx23920, 
      RST=>RST, EN=>nx23732, Q(15)=>OutputImg1_255_EXMPLR, Q(14)=>
      OutputImg1_254_EXMPLR, Q(13)=>OutputImg1_253_EXMPLR, Q(12)=>
      OutputImg1_252_EXMPLR, Q(11)=>OutputImg1_251_EXMPLR, Q(10)=>
      OutputImg1_250_EXMPLR, Q(9)=>OutputImg1_249_EXMPLR, Q(8)=>
      OutputImg1_248_EXMPLR, Q(7)=>OutputImg1_247_EXMPLR, Q(6)=>
      OutputImg1_246_EXMPLR, Q(5)=>OutputImg1_245_EXMPLR, Q(4)=>
      OutputImg1_244_EXMPLR, Q(3)=>OutputImg1_243_EXMPLR, Q(2)=>
      OutputImg1_242_EXMPLR, Q(1)=>OutputImg1_241_EXMPLR, Q(0)=>
      OutputImg1_240_EXMPLR);
   loop3_15_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_255, D(14)=>
      ImgReg2IN_254, D(13)=>ImgReg2IN_253, D(12)=>ImgReg2IN_252, D(11)=>
      ImgReg2IN_251, D(10)=>ImgReg2IN_250, D(9)=>ImgReg2IN_249, D(8)=>
      ImgReg2IN_248, D(7)=>ImgReg2IN_247, D(6)=>ImgReg2IN_246, D(5)=>
      ImgReg2IN_245, D(4)=>ImgReg2IN_244, D(3)=>ImgReg2IN_243, D(2)=>
      ImgReg2IN_242, D(1)=>ImgReg2IN_241, D(0)=>ImgReg2IN_240, CLK=>nx23920, 
      RST=>RST, EN=>nx23742, Q(15)=>OutputImg2_255_EXMPLR, Q(14)=>
      OutputImg2_254_EXMPLR, Q(13)=>OutputImg2_253_EXMPLR, Q(12)=>
      OutputImg2_252_EXMPLR, Q(11)=>OutputImg2_251_EXMPLR, Q(10)=>
      OutputImg2_250_EXMPLR, Q(9)=>OutputImg2_249_EXMPLR, Q(8)=>
      OutputImg2_248_EXMPLR, Q(7)=>OutputImg2_247_EXMPLR, Q(6)=>
      OutputImg2_246_EXMPLR, Q(5)=>OutputImg2_245_EXMPLR, Q(4)=>
      OutputImg2_244_EXMPLR, Q(3)=>OutputImg2_243_EXMPLR, Q(2)=>
      OutputImg2_242_EXMPLR, Q(1)=>OutputImg2_241_EXMPLR, Q(0)=>
      OutputImg2_240_EXMPLR);
   loop3_15_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_255, D(14)=>
      ImgReg3IN_254, D(13)=>ImgReg3IN_253, D(12)=>ImgReg3IN_252, D(11)=>
      ImgReg3IN_251, D(10)=>ImgReg3IN_250, D(9)=>ImgReg3IN_249, D(8)=>
      ImgReg3IN_248, D(7)=>ImgReg3IN_247, D(6)=>ImgReg3IN_246, D(5)=>
      ImgReg3IN_245, D(4)=>ImgReg3IN_244, D(3)=>ImgReg3IN_243, D(2)=>
      ImgReg3IN_242, D(1)=>ImgReg3IN_241, D(0)=>ImgReg3IN_240, CLK=>nx23922, 
      RST=>RST, EN=>nx23752, Q(15)=>OutputImg3_255_EXMPLR, Q(14)=>
      OutputImg3_254_EXMPLR, Q(13)=>OutputImg3_253_EXMPLR, Q(12)=>
      OutputImg3_252_EXMPLR, Q(11)=>OutputImg3_251_EXMPLR, Q(10)=>
      OutputImg3_250_EXMPLR, Q(9)=>OutputImg3_249_EXMPLR, Q(8)=>
      OutputImg3_248_EXMPLR, Q(7)=>OutputImg3_247_EXMPLR, Q(6)=>
      OutputImg3_246_EXMPLR, Q(5)=>OutputImg3_245_EXMPLR, Q(4)=>
      OutputImg3_244_EXMPLR, Q(3)=>OutputImg3_243_EXMPLR, Q(2)=>
      OutputImg3_242_EXMPLR, Q(1)=>OutputImg3_241_EXMPLR, Q(0)=>
      OutputImg3_240_EXMPLR);
   loop3_15_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_255, D(14)=>
      ImgReg4IN_254, D(13)=>ImgReg4IN_253, D(12)=>ImgReg4IN_252, D(11)=>
      ImgReg4IN_251, D(10)=>ImgReg4IN_250, D(9)=>ImgReg4IN_249, D(8)=>
      ImgReg4IN_248, D(7)=>ImgReg4IN_247, D(6)=>ImgReg4IN_246, D(5)=>
      ImgReg4IN_245, D(4)=>ImgReg4IN_244, D(3)=>ImgReg4IN_243, D(2)=>
      ImgReg4IN_242, D(1)=>ImgReg4IN_241, D(0)=>ImgReg4IN_240, CLK=>nx23922, 
      RST=>RST, EN=>nx23762, Q(15)=>OutputImg4_255_EXMPLR, Q(14)=>
      OutputImg4_254_EXMPLR, Q(13)=>OutputImg4_253_EXMPLR, Q(12)=>
      OutputImg4_252_EXMPLR, Q(11)=>OutputImg4_251_EXMPLR, Q(10)=>
      OutputImg4_250_EXMPLR, Q(9)=>OutputImg4_249_EXMPLR, Q(8)=>
      OutputImg4_248_EXMPLR, Q(7)=>OutputImg4_247_EXMPLR, Q(6)=>
      OutputImg4_246_EXMPLR, Q(5)=>OutputImg4_245_EXMPLR, Q(4)=>
      OutputImg4_244_EXMPLR, Q(3)=>OutputImg4_243_EXMPLR, Q(2)=>
      OutputImg4_242_EXMPLR, Q(1)=>OutputImg4_241_EXMPLR, Q(0)=>
      OutputImg4_240_EXMPLR);
   loop3_15_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_255, D(14)=>
      ImgReg5IN_254, D(13)=>ImgReg5IN_253, D(12)=>ImgReg5IN_252, D(11)=>
      ImgReg5IN_251, D(10)=>ImgReg5IN_250, D(9)=>ImgReg5IN_249, D(8)=>
      ImgReg5IN_248, D(7)=>ImgReg5IN_247, D(6)=>ImgReg5IN_246, D(5)=>
      ImgReg5IN_245, D(4)=>ImgReg5IN_244, D(3)=>ImgReg5IN_243, D(2)=>
      ImgReg5IN_242, D(1)=>ImgReg5IN_241, D(0)=>ImgReg5IN_240, CLK=>nx23924, 
      RST=>RST, EN=>nx23772, Q(15)=>OutputImg5_255_EXMPLR, Q(14)=>
      OutputImg5_254_EXMPLR, Q(13)=>OutputImg5_253_EXMPLR, Q(12)=>
      OutputImg5_252_EXMPLR, Q(11)=>OutputImg5_251_EXMPLR, Q(10)=>
      OutputImg5_250_EXMPLR, Q(9)=>OutputImg5_249_EXMPLR, Q(8)=>
      OutputImg5_248_EXMPLR, Q(7)=>OutputImg5_247_EXMPLR, Q(6)=>
      OutputImg5_246_EXMPLR, Q(5)=>OutputImg5_245_EXMPLR, Q(4)=>
      OutputImg5_244_EXMPLR, Q(3)=>OutputImg5_243_EXMPLR, Q(2)=>
      OutputImg5_242_EXMPLR, Q(1)=>OutputImg5_241_EXMPLR, Q(0)=>
      OutputImg5_240_EXMPLR);
   loop3_16_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_287_EXMPLR, D(14)=>OutputImg0_286_EXMPLR, D(13)=>
      OutputImg0_285_EXMPLR, D(12)=>OutputImg0_284_EXMPLR, D(11)=>
      OutputImg0_283_EXMPLR, D(10)=>OutputImg0_282_EXMPLR, D(9)=>
      OutputImg0_281_EXMPLR, D(8)=>OutputImg0_280_EXMPLR, D(7)=>
      OutputImg0_279_EXMPLR, D(6)=>OutputImg0_278_EXMPLR, D(5)=>
      OutputImg0_277_EXMPLR, D(4)=>OutputImg0_276_EXMPLR, D(3)=>
      OutputImg0_275_EXMPLR, D(2)=>OutputImg0_274_EXMPLR, D(1)=>
      OutputImg0_273_EXMPLR, D(0)=>OutputImg0_272_EXMPLR, EN=>nx23692, F(15)
      =>ImgReg0IN_271, F(14)=>ImgReg0IN_270, F(13)=>ImgReg0IN_269, F(12)=>
      ImgReg0IN_268, F(11)=>ImgReg0IN_267, F(10)=>ImgReg0IN_266, F(9)=>
      ImgReg0IN_265, F(8)=>ImgReg0IN_264, F(7)=>ImgReg0IN_263, F(6)=>
      ImgReg0IN_262, F(5)=>ImgReg0IN_261, F(4)=>ImgReg0IN_260, F(3)=>
      ImgReg0IN_259, F(2)=>ImgReg0IN_258, F(1)=>ImgReg0IN_257, F(0)=>
      ImgReg0IN_256);
   loop3_16_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_287_EXMPLR, D(14)=>OutputImg1_286_EXMPLR, D(13)=>
      OutputImg1_285_EXMPLR, D(12)=>OutputImg1_284_EXMPLR, D(11)=>
      OutputImg1_283_EXMPLR, D(10)=>OutputImg1_282_EXMPLR, D(9)=>
      OutputImg1_281_EXMPLR, D(8)=>OutputImg1_280_EXMPLR, D(7)=>
      OutputImg1_279_EXMPLR, D(6)=>OutputImg1_278_EXMPLR, D(5)=>
      OutputImg1_277_EXMPLR, D(4)=>OutputImg1_276_EXMPLR, D(3)=>
      OutputImg1_275_EXMPLR, D(2)=>OutputImg1_274_EXMPLR, D(1)=>
      OutputImg1_273_EXMPLR, D(0)=>OutputImg1_272_EXMPLR, EN=>nx23692, F(15)
      =>ImgReg1IN_271, F(14)=>ImgReg1IN_270, F(13)=>ImgReg1IN_269, F(12)=>
      ImgReg1IN_268, F(11)=>ImgReg1IN_267, F(10)=>ImgReg1IN_266, F(9)=>
      ImgReg1IN_265, F(8)=>ImgReg1IN_264, F(7)=>ImgReg1IN_263, F(6)=>
      ImgReg1IN_262, F(5)=>ImgReg1IN_261, F(4)=>ImgReg1IN_260, F(3)=>
      ImgReg1IN_259, F(2)=>ImgReg1IN_258, F(1)=>ImgReg1IN_257, F(0)=>
      ImgReg1IN_256);
   loop3_16_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_287_EXMPLR, D(14)=>OutputImg2_286_EXMPLR, D(13)=>
      OutputImg2_285_EXMPLR, D(12)=>OutputImg2_284_EXMPLR, D(11)=>
      OutputImg2_283_EXMPLR, D(10)=>OutputImg2_282_EXMPLR, D(9)=>
      OutputImg2_281_EXMPLR, D(8)=>OutputImg2_280_EXMPLR, D(7)=>
      OutputImg2_279_EXMPLR, D(6)=>OutputImg2_278_EXMPLR, D(5)=>
      OutputImg2_277_EXMPLR, D(4)=>OutputImg2_276_EXMPLR, D(3)=>
      OutputImg2_275_EXMPLR, D(2)=>OutputImg2_274_EXMPLR, D(1)=>
      OutputImg2_273_EXMPLR, D(0)=>OutputImg2_272_EXMPLR, EN=>nx23694, F(15)
      =>ImgReg2IN_271, F(14)=>ImgReg2IN_270, F(13)=>ImgReg2IN_269, F(12)=>
      ImgReg2IN_268, F(11)=>ImgReg2IN_267, F(10)=>ImgReg2IN_266, F(9)=>
      ImgReg2IN_265, F(8)=>ImgReg2IN_264, F(7)=>ImgReg2IN_263, F(6)=>
      ImgReg2IN_262, F(5)=>ImgReg2IN_261, F(4)=>ImgReg2IN_260, F(3)=>
      ImgReg2IN_259, F(2)=>ImgReg2IN_258, F(1)=>ImgReg2IN_257, F(0)=>
      ImgReg2IN_256);
   loop3_16_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_287_EXMPLR, D(14)=>OutputImg3_286_EXMPLR, D(13)=>
      OutputImg3_285_EXMPLR, D(12)=>OutputImg3_284_EXMPLR, D(11)=>
      OutputImg3_283_EXMPLR, D(10)=>OutputImg3_282_EXMPLR, D(9)=>
      OutputImg3_281_EXMPLR, D(8)=>OutputImg3_280_EXMPLR, D(7)=>
      OutputImg3_279_EXMPLR, D(6)=>OutputImg3_278_EXMPLR, D(5)=>
      OutputImg3_277_EXMPLR, D(4)=>OutputImg3_276_EXMPLR, D(3)=>
      OutputImg3_275_EXMPLR, D(2)=>OutputImg3_274_EXMPLR, D(1)=>
      OutputImg3_273_EXMPLR, D(0)=>OutputImg3_272_EXMPLR, EN=>nx23694, F(15)
      =>ImgReg3IN_271, F(14)=>ImgReg3IN_270, F(13)=>ImgReg3IN_269, F(12)=>
      ImgReg3IN_268, F(11)=>ImgReg3IN_267, F(10)=>ImgReg3IN_266, F(9)=>
      ImgReg3IN_265, F(8)=>ImgReg3IN_264, F(7)=>ImgReg3IN_263, F(6)=>
      ImgReg3IN_262, F(5)=>ImgReg3IN_261, F(4)=>ImgReg3IN_260, F(3)=>
      ImgReg3IN_259, F(2)=>ImgReg3IN_258, F(1)=>ImgReg3IN_257, F(0)=>
      ImgReg3IN_256);
   loop3_16_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_287_EXMPLR, D(14)=>OutputImg4_286_EXMPLR, D(13)=>
      OutputImg4_285_EXMPLR, D(12)=>OutputImg4_284_EXMPLR, D(11)=>
      OutputImg4_283_EXMPLR, D(10)=>OutputImg4_282_EXMPLR, D(9)=>
      OutputImg4_281_EXMPLR, D(8)=>OutputImg4_280_EXMPLR, D(7)=>
      OutputImg4_279_EXMPLR, D(6)=>OutputImg4_278_EXMPLR, D(5)=>
      OutputImg4_277_EXMPLR, D(4)=>OutputImg4_276_EXMPLR, D(3)=>
      OutputImg4_275_EXMPLR, D(2)=>OutputImg4_274_EXMPLR, D(1)=>
      OutputImg4_273_EXMPLR, D(0)=>OutputImg4_272_EXMPLR, EN=>nx23694, F(15)
      =>ImgReg4IN_271, F(14)=>ImgReg4IN_270, F(13)=>ImgReg4IN_269, F(12)=>
      ImgReg4IN_268, F(11)=>ImgReg4IN_267, F(10)=>ImgReg4IN_266, F(9)=>
      ImgReg4IN_265, F(8)=>ImgReg4IN_264, F(7)=>ImgReg4IN_263, F(6)=>
      ImgReg4IN_262, F(5)=>ImgReg4IN_261, F(4)=>ImgReg4IN_260, F(3)=>
      ImgReg4IN_259, F(2)=>ImgReg4IN_258, F(1)=>ImgReg4IN_257, F(0)=>
      ImgReg4IN_256);
   loop3_16_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_287_EXMPLR, D(14)=>OutputImg5_286_EXMPLR, D(13)=>
      OutputImg5_285_EXMPLR, D(12)=>OutputImg5_284_EXMPLR, D(11)=>
      OutputImg5_283_EXMPLR, D(10)=>OutputImg5_282_EXMPLR, D(9)=>
      OutputImg5_281_EXMPLR, D(8)=>OutputImg5_280_EXMPLR, D(7)=>
      OutputImg5_279_EXMPLR, D(6)=>OutputImg5_278_EXMPLR, D(5)=>
      OutputImg5_277_EXMPLR, D(4)=>OutputImg5_276_EXMPLR, D(3)=>
      OutputImg5_275_EXMPLR, D(2)=>OutputImg5_274_EXMPLR, D(1)=>
      OutputImg5_273_EXMPLR, D(0)=>OutputImg5_272_EXMPLR, EN=>nx23694, F(15)
      =>ImgReg5IN_271, F(14)=>ImgReg5IN_270, F(13)=>ImgReg5IN_269, F(12)=>
      ImgReg5IN_268, F(11)=>ImgReg5IN_267, F(10)=>ImgReg5IN_266, F(9)=>
      ImgReg5IN_265, F(8)=>ImgReg5IN_264, F(7)=>ImgReg5IN_263, F(6)=>
      ImgReg5IN_262, F(5)=>ImgReg5IN_261, F(4)=>ImgReg5IN_260, F(3)=>
      ImgReg5IN_259, F(2)=>ImgReg5IN_258, F(1)=>ImgReg5IN_257, F(0)=>
      ImgReg5IN_256);
   loop3_16_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(271), 
      D(14)=>DATA(270), D(13)=>DATA(269), D(12)=>DATA(268), D(11)=>DATA(267), 
      D(10)=>DATA(266), D(9)=>DATA(265), D(8)=>DATA(264), D(7)=>DATA(263), 
      D(6)=>DATA(262), D(5)=>DATA(261), D(4)=>DATA(260), D(3)=>DATA(259), 
      D(2)=>DATA(258), D(1)=>DATA(257), D(0)=>DATA(256), EN=>nx23658, F(15)
      =>ImgReg0IN_271, F(14)=>ImgReg0IN_270, F(13)=>ImgReg0IN_269, F(12)=>
      ImgReg0IN_268, F(11)=>ImgReg0IN_267, F(10)=>ImgReg0IN_266, F(9)=>
      ImgReg0IN_265, F(8)=>ImgReg0IN_264, F(7)=>ImgReg0IN_263, F(6)=>
      ImgReg0IN_262, F(5)=>ImgReg0IN_261, F(4)=>ImgReg0IN_260, F(3)=>
      ImgReg0IN_259, F(2)=>ImgReg0IN_258, F(1)=>ImgReg0IN_257, F(0)=>
      ImgReg0IN_256);
   loop3_16_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(271), 
      D(14)=>DATA(270), D(13)=>DATA(269), D(12)=>DATA(268), D(11)=>DATA(267), 
      D(10)=>DATA(266), D(9)=>DATA(265), D(8)=>DATA(264), D(7)=>DATA(263), 
      D(6)=>DATA(262), D(5)=>DATA(261), D(4)=>DATA(260), D(3)=>DATA(259), 
      D(2)=>DATA(258), D(1)=>DATA(257), D(0)=>DATA(256), EN=>nx23646, F(15)
      =>ImgReg1IN_271, F(14)=>ImgReg1IN_270, F(13)=>ImgReg1IN_269, F(12)=>
      ImgReg1IN_268, F(11)=>ImgReg1IN_267, F(10)=>ImgReg1IN_266, F(9)=>
      ImgReg1IN_265, F(8)=>ImgReg1IN_264, F(7)=>ImgReg1IN_263, F(6)=>
      ImgReg1IN_262, F(5)=>ImgReg1IN_261, F(4)=>ImgReg1IN_260, F(3)=>
      ImgReg1IN_259, F(2)=>ImgReg1IN_258, F(1)=>ImgReg1IN_257, F(0)=>
      ImgReg1IN_256);
   loop3_16_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(271), 
      D(14)=>DATA(270), D(13)=>DATA(269), D(12)=>DATA(268), D(11)=>DATA(267), 
      D(10)=>DATA(266), D(9)=>DATA(265), D(8)=>DATA(264), D(7)=>DATA(263), 
      D(6)=>DATA(262), D(5)=>DATA(261), D(4)=>DATA(260), D(3)=>DATA(259), 
      D(2)=>DATA(258), D(1)=>DATA(257), D(0)=>DATA(256), EN=>nx23634, F(15)
      =>ImgReg2IN_271, F(14)=>ImgReg2IN_270, F(13)=>ImgReg2IN_269, F(12)=>
      ImgReg2IN_268, F(11)=>ImgReg2IN_267, F(10)=>ImgReg2IN_266, F(9)=>
      ImgReg2IN_265, F(8)=>ImgReg2IN_264, F(7)=>ImgReg2IN_263, F(6)=>
      ImgReg2IN_262, F(5)=>ImgReg2IN_261, F(4)=>ImgReg2IN_260, F(3)=>
      ImgReg2IN_259, F(2)=>ImgReg2IN_258, F(1)=>ImgReg2IN_257, F(0)=>
      ImgReg2IN_256);
   loop3_16_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(271), 
      D(14)=>DATA(270), D(13)=>DATA(269), D(12)=>DATA(268), D(11)=>DATA(267), 
      D(10)=>DATA(266), D(9)=>DATA(265), D(8)=>DATA(264), D(7)=>DATA(263), 
      D(6)=>DATA(262), D(5)=>DATA(261), D(4)=>DATA(260), D(3)=>DATA(259), 
      D(2)=>DATA(258), D(1)=>DATA(257), D(0)=>DATA(256), EN=>nx23622, F(15)
      =>ImgReg3IN_271, F(14)=>ImgReg3IN_270, F(13)=>ImgReg3IN_269, F(12)=>
      ImgReg3IN_268, F(11)=>ImgReg3IN_267, F(10)=>ImgReg3IN_266, F(9)=>
      ImgReg3IN_265, F(8)=>ImgReg3IN_264, F(7)=>ImgReg3IN_263, F(6)=>
      ImgReg3IN_262, F(5)=>ImgReg3IN_261, F(4)=>ImgReg3IN_260, F(3)=>
      ImgReg3IN_259, F(2)=>ImgReg3IN_258, F(1)=>ImgReg3IN_257, F(0)=>
      ImgReg3IN_256);
   loop3_16_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(271), 
      D(14)=>DATA(270), D(13)=>DATA(269), D(12)=>DATA(268), D(11)=>DATA(267), 
      D(10)=>DATA(266), D(9)=>DATA(265), D(8)=>DATA(264), D(7)=>DATA(263), 
      D(6)=>DATA(262), D(5)=>DATA(261), D(4)=>DATA(260), D(3)=>DATA(259), 
      D(2)=>DATA(258), D(1)=>DATA(257), D(0)=>DATA(256), EN=>nx23610, F(15)
      =>ImgReg4IN_271, F(14)=>ImgReg4IN_270, F(13)=>ImgReg4IN_269, F(12)=>
      ImgReg4IN_268, F(11)=>ImgReg4IN_267, F(10)=>ImgReg4IN_266, F(9)=>
      ImgReg4IN_265, F(8)=>ImgReg4IN_264, F(7)=>ImgReg4IN_263, F(6)=>
      ImgReg4IN_262, F(5)=>ImgReg4IN_261, F(4)=>ImgReg4IN_260, F(3)=>
      ImgReg4IN_259, F(2)=>ImgReg4IN_258, F(1)=>ImgReg4IN_257, F(0)=>
      ImgReg4IN_256);
   loop3_16_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(271), 
      D(14)=>DATA(270), D(13)=>DATA(269), D(12)=>DATA(268), D(11)=>DATA(267), 
      D(10)=>DATA(266), D(9)=>DATA(265), D(8)=>DATA(264), D(7)=>DATA(263), 
      D(6)=>DATA(262), D(5)=>DATA(261), D(4)=>DATA(260), D(3)=>DATA(259), 
      D(2)=>DATA(258), D(1)=>DATA(257), D(0)=>DATA(256), EN=>nx23598, F(15)
      =>ImgReg5IN_271, F(14)=>ImgReg5IN_270, F(13)=>ImgReg5IN_269, F(12)=>
      ImgReg5IN_268, F(11)=>ImgReg5IN_267, F(10)=>ImgReg5IN_266, F(9)=>
      ImgReg5IN_265, F(8)=>ImgReg5IN_264, F(7)=>ImgReg5IN_263, F(6)=>
      ImgReg5IN_262, F(5)=>ImgReg5IN_261, F(4)=>ImgReg5IN_260, F(3)=>
      ImgReg5IN_259, F(2)=>ImgReg5IN_258, F(1)=>ImgReg5IN_257, F(0)=>
      ImgReg5IN_256);
   loop3_16_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_271_EXMPLR, D(14)=>OutputImg1_270_EXMPLR, D(13)=>
      OutputImg1_269_EXMPLR, D(12)=>OutputImg1_268_EXMPLR, D(11)=>
      OutputImg1_267_EXMPLR, D(10)=>OutputImg1_266_EXMPLR, D(9)=>
      OutputImg1_265_EXMPLR, D(8)=>OutputImg1_264_EXMPLR, D(7)=>
      OutputImg1_263_EXMPLR, D(6)=>OutputImg1_262_EXMPLR, D(5)=>
      OutputImg1_261_EXMPLR, D(4)=>OutputImg1_260_EXMPLR, D(3)=>
      OutputImg1_259_EXMPLR, D(2)=>OutputImg1_258_EXMPLR, D(1)=>
      OutputImg1_257_EXMPLR, D(0)=>OutputImg1_256_EXMPLR, EN=>nx23808, F(15)
      =>ImgReg0IN_271, F(14)=>ImgReg0IN_270, F(13)=>ImgReg0IN_269, F(12)=>
      ImgReg0IN_268, F(11)=>ImgReg0IN_267, F(10)=>ImgReg0IN_266, F(9)=>
      ImgReg0IN_265, F(8)=>ImgReg0IN_264, F(7)=>ImgReg0IN_263, F(6)=>
      ImgReg0IN_262, F(5)=>ImgReg0IN_261, F(4)=>ImgReg0IN_260, F(3)=>
      ImgReg0IN_259, F(2)=>ImgReg0IN_258, F(1)=>ImgReg0IN_257, F(0)=>
      ImgReg0IN_256);
   loop3_16_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_271_EXMPLR, D(14)=>OutputImg2_270_EXMPLR, D(13)=>
      OutputImg2_269_EXMPLR, D(12)=>OutputImg2_268_EXMPLR, D(11)=>
      OutputImg2_267_EXMPLR, D(10)=>OutputImg2_266_EXMPLR, D(9)=>
      OutputImg2_265_EXMPLR, D(8)=>OutputImg2_264_EXMPLR, D(7)=>
      OutputImg2_263_EXMPLR, D(6)=>OutputImg2_262_EXMPLR, D(5)=>
      OutputImg2_261_EXMPLR, D(4)=>OutputImg2_260_EXMPLR, D(3)=>
      OutputImg2_259_EXMPLR, D(2)=>OutputImg2_258_EXMPLR, D(1)=>
      OutputImg2_257_EXMPLR, D(0)=>OutputImg2_256_EXMPLR, EN=>nx23808, F(15)
      =>ImgReg1IN_271, F(14)=>ImgReg1IN_270, F(13)=>ImgReg1IN_269, F(12)=>
      ImgReg1IN_268, F(11)=>ImgReg1IN_267, F(10)=>ImgReg1IN_266, F(9)=>
      ImgReg1IN_265, F(8)=>ImgReg1IN_264, F(7)=>ImgReg1IN_263, F(6)=>
      ImgReg1IN_262, F(5)=>ImgReg1IN_261, F(4)=>ImgReg1IN_260, F(3)=>
      ImgReg1IN_259, F(2)=>ImgReg1IN_258, F(1)=>ImgReg1IN_257, F(0)=>
      ImgReg1IN_256);
   loop3_16_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_271_EXMPLR, D(14)=>OutputImg3_270_EXMPLR, D(13)=>
      OutputImg3_269_EXMPLR, D(12)=>OutputImg3_268_EXMPLR, D(11)=>
      OutputImg3_267_EXMPLR, D(10)=>OutputImg3_266_EXMPLR, D(9)=>
      OutputImg3_265_EXMPLR, D(8)=>OutputImg3_264_EXMPLR, D(7)=>
      OutputImg3_263_EXMPLR, D(6)=>OutputImg3_262_EXMPLR, D(5)=>
      OutputImg3_261_EXMPLR, D(4)=>OutputImg3_260_EXMPLR, D(3)=>
      OutputImg3_259_EXMPLR, D(2)=>OutputImg3_258_EXMPLR, D(1)=>
      OutputImg3_257_EXMPLR, D(0)=>OutputImg3_256_EXMPLR, EN=>nx23808, F(15)
      =>ImgReg2IN_271, F(14)=>ImgReg2IN_270, F(13)=>ImgReg2IN_269, F(12)=>
      ImgReg2IN_268, F(11)=>ImgReg2IN_267, F(10)=>ImgReg2IN_266, F(9)=>
      ImgReg2IN_265, F(8)=>ImgReg2IN_264, F(7)=>ImgReg2IN_263, F(6)=>
      ImgReg2IN_262, F(5)=>ImgReg2IN_261, F(4)=>ImgReg2IN_260, F(3)=>
      ImgReg2IN_259, F(2)=>ImgReg2IN_258, F(1)=>ImgReg2IN_257, F(0)=>
      ImgReg2IN_256);
   loop3_16_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_271_EXMPLR, D(14)=>OutputImg4_270_EXMPLR, D(13)=>
      OutputImg4_269_EXMPLR, D(12)=>OutputImg4_268_EXMPLR, D(11)=>
      OutputImg4_267_EXMPLR, D(10)=>OutputImg4_266_EXMPLR, D(9)=>
      OutputImg4_265_EXMPLR, D(8)=>OutputImg4_264_EXMPLR, D(7)=>
      OutputImg4_263_EXMPLR, D(6)=>OutputImg4_262_EXMPLR, D(5)=>
      OutputImg4_261_EXMPLR, D(4)=>OutputImg4_260_EXMPLR, D(3)=>
      OutputImg4_259_EXMPLR, D(2)=>OutputImg4_258_EXMPLR, D(1)=>
      OutputImg4_257_EXMPLR, D(0)=>OutputImg4_256_EXMPLR, EN=>nx23808, F(15)
      =>ImgReg3IN_271, F(14)=>ImgReg3IN_270, F(13)=>ImgReg3IN_269, F(12)=>
      ImgReg3IN_268, F(11)=>ImgReg3IN_267, F(10)=>ImgReg3IN_266, F(9)=>
      ImgReg3IN_265, F(8)=>ImgReg3IN_264, F(7)=>ImgReg3IN_263, F(6)=>
      ImgReg3IN_262, F(5)=>ImgReg3IN_261, F(4)=>ImgReg3IN_260, F(3)=>
      ImgReg3IN_259, F(2)=>ImgReg3IN_258, F(1)=>ImgReg3IN_257, F(0)=>
      ImgReg3IN_256);
   loop3_16_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_271_EXMPLR, D(14)=>OutputImg5_270_EXMPLR, D(13)=>
      OutputImg5_269_EXMPLR, D(12)=>OutputImg5_268_EXMPLR, D(11)=>
      OutputImg5_267_EXMPLR, D(10)=>OutputImg5_266_EXMPLR, D(9)=>
      OutputImg5_265_EXMPLR, D(8)=>OutputImg5_264_EXMPLR, D(7)=>
      OutputImg5_263_EXMPLR, D(6)=>OutputImg5_262_EXMPLR, D(5)=>
      OutputImg5_261_EXMPLR, D(4)=>OutputImg5_260_EXMPLR, D(3)=>
      OutputImg5_259_EXMPLR, D(2)=>OutputImg5_258_EXMPLR, D(1)=>
      OutputImg5_257_EXMPLR, D(0)=>OutputImg5_256_EXMPLR, EN=>nx23810, F(15)
      =>ImgReg4IN_271, F(14)=>ImgReg4IN_270, F(13)=>ImgReg4IN_269, F(12)=>
      ImgReg4IN_268, F(11)=>ImgReg4IN_267, F(10)=>ImgReg4IN_266, F(9)=>
      ImgReg4IN_265, F(8)=>ImgReg4IN_264, F(7)=>ImgReg4IN_263, F(6)=>
      ImgReg4IN_262, F(5)=>ImgReg4IN_261, F(4)=>ImgReg4IN_260, F(3)=>
      ImgReg4IN_259, F(2)=>ImgReg4IN_258, F(1)=>ImgReg4IN_257, F(0)=>
      ImgReg4IN_256);
   loop3_16_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_271, D(14)=>
      ImgReg0IN_270, D(13)=>ImgReg0IN_269, D(12)=>ImgReg0IN_268, D(11)=>
      ImgReg0IN_267, D(10)=>ImgReg0IN_266, D(9)=>ImgReg0IN_265, D(8)=>
      ImgReg0IN_264, D(7)=>ImgReg0IN_263, D(6)=>ImgReg0IN_262, D(5)=>
      ImgReg0IN_261, D(4)=>ImgReg0IN_260, D(3)=>ImgReg0IN_259, D(2)=>
      ImgReg0IN_258, D(1)=>ImgReg0IN_257, D(0)=>ImgReg0IN_256, CLK=>nx23924, 
      RST=>RST, EN=>nx23722, Q(15)=>OutputImg0_271_EXMPLR, Q(14)=>
      OutputImg0_270_EXMPLR, Q(13)=>OutputImg0_269_EXMPLR, Q(12)=>
      OutputImg0_268_EXMPLR, Q(11)=>OutputImg0_267_EXMPLR, Q(10)=>
      OutputImg0_266_EXMPLR, Q(9)=>OutputImg0_265_EXMPLR, Q(8)=>
      OutputImg0_264_EXMPLR, Q(7)=>OutputImg0_263_EXMPLR, Q(6)=>
      OutputImg0_262_EXMPLR, Q(5)=>OutputImg0_261_EXMPLR, Q(4)=>
      OutputImg0_260_EXMPLR, Q(3)=>OutputImg0_259_EXMPLR, Q(2)=>
      OutputImg0_258_EXMPLR, Q(1)=>OutputImg0_257_EXMPLR, Q(0)=>
      OutputImg0_256_EXMPLR);
   loop3_16_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_271, D(14)=>
      ImgReg1IN_270, D(13)=>ImgReg1IN_269, D(12)=>ImgReg1IN_268, D(11)=>
      ImgReg1IN_267, D(10)=>ImgReg1IN_266, D(9)=>ImgReg1IN_265, D(8)=>
      ImgReg1IN_264, D(7)=>ImgReg1IN_263, D(6)=>ImgReg1IN_262, D(5)=>
      ImgReg1IN_261, D(4)=>ImgReg1IN_260, D(3)=>ImgReg1IN_259, D(2)=>
      ImgReg1IN_258, D(1)=>ImgReg1IN_257, D(0)=>ImgReg1IN_256, CLK=>nx23926, 
      RST=>RST, EN=>nx23732, Q(15)=>OutputImg1_271_EXMPLR, Q(14)=>
      OutputImg1_270_EXMPLR, Q(13)=>OutputImg1_269_EXMPLR, Q(12)=>
      OutputImg1_268_EXMPLR, Q(11)=>OutputImg1_267_EXMPLR, Q(10)=>
      OutputImg1_266_EXMPLR, Q(9)=>OutputImg1_265_EXMPLR, Q(8)=>
      OutputImg1_264_EXMPLR, Q(7)=>OutputImg1_263_EXMPLR, Q(6)=>
      OutputImg1_262_EXMPLR, Q(5)=>OutputImg1_261_EXMPLR, Q(4)=>
      OutputImg1_260_EXMPLR, Q(3)=>OutputImg1_259_EXMPLR, Q(2)=>
      OutputImg1_258_EXMPLR, Q(1)=>OutputImg1_257_EXMPLR, Q(0)=>
      OutputImg1_256_EXMPLR);
   loop3_16_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_271, D(14)=>
      ImgReg2IN_270, D(13)=>ImgReg2IN_269, D(12)=>ImgReg2IN_268, D(11)=>
      ImgReg2IN_267, D(10)=>ImgReg2IN_266, D(9)=>ImgReg2IN_265, D(8)=>
      ImgReg2IN_264, D(7)=>ImgReg2IN_263, D(6)=>ImgReg2IN_262, D(5)=>
      ImgReg2IN_261, D(4)=>ImgReg2IN_260, D(3)=>ImgReg2IN_259, D(2)=>
      ImgReg2IN_258, D(1)=>ImgReg2IN_257, D(0)=>ImgReg2IN_256, CLK=>nx23926, 
      RST=>RST, EN=>nx23742, Q(15)=>OutputImg2_271_EXMPLR, Q(14)=>
      OutputImg2_270_EXMPLR, Q(13)=>OutputImg2_269_EXMPLR, Q(12)=>
      OutputImg2_268_EXMPLR, Q(11)=>OutputImg2_267_EXMPLR, Q(10)=>
      OutputImg2_266_EXMPLR, Q(9)=>OutputImg2_265_EXMPLR, Q(8)=>
      OutputImg2_264_EXMPLR, Q(7)=>OutputImg2_263_EXMPLR, Q(6)=>
      OutputImg2_262_EXMPLR, Q(5)=>OutputImg2_261_EXMPLR, Q(4)=>
      OutputImg2_260_EXMPLR, Q(3)=>OutputImg2_259_EXMPLR, Q(2)=>
      OutputImg2_258_EXMPLR, Q(1)=>OutputImg2_257_EXMPLR, Q(0)=>
      OutputImg2_256_EXMPLR);
   loop3_16_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_271, D(14)=>
      ImgReg3IN_270, D(13)=>ImgReg3IN_269, D(12)=>ImgReg3IN_268, D(11)=>
      ImgReg3IN_267, D(10)=>ImgReg3IN_266, D(9)=>ImgReg3IN_265, D(8)=>
      ImgReg3IN_264, D(7)=>ImgReg3IN_263, D(6)=>ImgReg3IN_262, D(5)=>
      ImgReg3IN_261, D(4)=>ImgReg3IN_260, D(3)=>ImgReg3IN_259, D(2)=>
      ImgReg3IN_258, D(1)=>ImgReg3IN_257, D(0)=>ImgReg3IN_256, CLK=>nx23928, 
      RST=>RST, EN=>nx23752, Q(15)=>OutputImg3_271_EXMPLR, Q(14)=>
      OutputImg3_270_EXMPLR, Q(13)=>OutputImg3_269_EXMPLR, Q(12)=>
      OutputImg3_268_EXMPLR, Q(11)=>OutputImg3_267_EXMPLR, Q(10)=>
      OutputImg3_266_EXMPLR, Q(9)=>OutputImg3_265_EXMPLR, Q(8)=>
      OutputImg3_264_EXMPLR, Q(7)=>OutputImg3_263_EXMPLR, Q(6)=>
      OutputImg3_262_EXMPLR, Q(5)=>OutputImg3_261_EXMPLR, Q(4)=>
      OutputImg3_260_EXMPLR, Q(3)=>OutputImg3_259_EXMPLR, Q(2)=>
      OutputImg3_258_EXMPLR, Q(1)=>OutputImg3_257_EXMPLR, Q(0)=>
      OutputImg3_256_EXMPLR);
   loop3_16_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_271, D(14)=>
      ImgReg4IN_270, D(13)=>ImgReg4IN_269, D(12)=>ImgReg4IN_268, D(11)=>
      ImgReg4IN_267, D(10)=>ImgReg4IN_266, D(9)=>ImgReg4IN_265, D(8)=>
      ImgReg4IN_264, D(7)=>ImgReg4IN_263, D(6)=>ImgReg4IN_262, D(5)=>
      ImgReg4IN_261, D(4)=>ImgReg4IN_260, D(3)=>ImgReg4IN_259, D(2)=>
      ImgReg4IN_258, D(1)=>ImgReg4IN_257, D(0)=>ImgReg4IN_256, CLK=>nx23928, 
      RST=>RST, EN=>nx23762, Q(15)=>OutputImg4_271_EXMPLR, Q(14)=>
      OutputImg4_270_EXMPLR, Q(13)=>OutputImg4_269_EXMPLR, Q(12)=>
      OutputImg4_268_EXMPLR, Q(11)=>OutputImg4_267_EXMPLR, Q(10)=>
      OutputImg4_266_EXMPLR, Q(9)=>OutputImg4_265_EXMPLR, Q(8)=>
      OutputImg4_264_EXMPLR, Q(7)=>OutputImg4_263_EXMPLR, Q(6)=>
      OutputImg4_262_EXMPLR, Q(5)=>OutputImg4_261_EXMPLR, Q(4)=>
      OutputImg4_260_EXMPLR, Q(3)=>OutputImg4_259_EXMPLR, Q(2)=>
      OutputImg4_258_EXMPLR, Q(1)=>OutputImg4_257_EXMPLR, Q(0)=>
      OutputImg4_256_EXMPLR);
   loop3_16_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_271, D(14)=>
      ImgReg5IN_270, D(13)=>ImgReg5IN_269, D(12)=>ImgReg5IN_268, D(11)=>
      ImgReg5IN_267, D(10)=>ImgReg5IN_266, D(9)=>ImgReg5IN_265, D(8)=>
      ImgReg5IN_264, D(7)=>ImgReg5IN_263, D(6)=>ImgReg5IN_262, D(5)=>
      ImgReg5IN_261, D(4)=>ImgReg5IN_260, D(3)=>ImgReg5IN_259, D(2)=>
      ImgReg5IN_258, D(1)=>ImgReg5IN_257, D(0)=>ImgReg5IN_256, CLK=>nx23930, 
      RST=>RST, EN=>nx23772, Q(15)=>OutputImg5_271_EXMPLR, Q(14)=>
      OutputImg5_270_EXMPLR, Q(13)=>OutputImg5_269_EXMPLR, Q(12)=>
      OutputImg5_268_EXMPLR, Q(11)=>OutputImg5_267_EXMPLR, Q(10)=>
      OutputImg5_266_EXMPLR, Q(9)=>OutputImg5_265_EXMPLR, Q(8)=>
      OutputImg5_264_EXMPLR, Q(7)=>OutputImg5_263_EXMPLR, Q(6)=>
      OutputImg5_262_EXMPLR, Q(5)=>OutputImg5_261_EXMPLR, Q(4)=>
      OutputImg5_260_EXMPLR, Q(3)=>OutputImg5_259_EXMPLR, Q(2)=>
      OutputImg5_258_EXMPLR, Q(1)=>OutputImg5_257_EXMPLR, Q(0)=>
      OutputImg5_256_EXMPLR);
   loop3_17_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_303_EXMPLR, D(14)=>OutputImg0_302_EXMPLR, D(13)=>
      OutputImg0_301_EXMPLR, D(12)=>OutputImg0_300_EXMPLR, D(11)=>
      OutputImg0_299_EXMPLR, D(10)=>OutputImg0_298_EXMPLR, D(9)=>
      OutputImg0_297_EXMPLR, D(8)=>OutputImg0_296_EXMPLR, D(7)=>
      OutputImg0_295_EXMPLR, D(6)=>OutputImg0_294_EXMPLR, D(5)=>
      OutputImg0_293_EXMPLR, D(4)=>OutputImg0_292_EXMPLR, D(3)=>
      OutputImg0_291_EXMPLR, D(2)=>OutputImg0_290_EXMPLR, D(1)=>
      OutputImg0_289_EXMPLR, D(0)=>OutputImg0_288_EXMPLR, EN=>nx23694, F(15)
      =>ImgReg0IN_287, F(14)=>ImgReg0IN_286, F(13)=>ImgReg0IN_285, F(12)=>
      ImgReg0IN_284, F(11)=>ImgReg0IN_283, F(10)=>ImgReg0IN_282, F(9)=>
      ImgReg0IN_281, F(8)=>ImgReg0IN_280, F(7)=>ImgReg0IN_279, F(6)=>
      ImgReg0IN_278, F(5)=>ImgReg0IN_277, F(4)=>ImgReg0IN_276, F(3)=>
      ImgReg0IN_275, F(2)=>ImgReg0IN_274, F(1)=>ImgReg0IN_273, F(0)=>
      ImgReg0IN_272);
   loop3_17_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_303_EXMPLR, D(14)=>OutputImg1_302_EXMPLR, D(13)=>
      OutputImg1_301_EXMPLR, D(12)=>OutputImg1_300_EXMPLR, D(11)=>
      OutputImg1_299_EXMPLR, D(10)=>OutputImg1_298_EXMPLR, D(9)=>
      OutputImg1_297_EXMPLR, D(8)=>OutputImg1_296_EXMPLR, D(7)=>
      OutputImg1_295_EXMPLR, D(6)=>OutputImg1_294_EXMPLR, D(5)=>
      OutputImg1_293_EXMPLR, D(4)=>OutputImg1_292_EXMPLR, D(3)=>
      OutputImg1_291_EXMPLR, D(2)=>OutputImg1_290_EXMPLR, D(1)=>
      OutputImg1_289_EXMPLR, D(0)=>OutputImg1_288_EXMPLR, EN=>nx23694, F(15)
      =>ImgReg1IN_287, F(14)=>ImgReg1IN_286, F(13)=>ImgReg1IN_285, F(12)=>
      ImgReg1IN_284, F(11)=>ImgReg1IN_283, F(10)=>ImgReg1IN_282, F(9)=>
      ImgReg1IN_281, F(8)=>ImgReg1IN_280, F(7)=>ImgReg1IN_279, F(6)=>
      ImgReg1IN_278, F(5)=>ImgReg1IN_277, F(4)=>ImgReg1IN_276, F(3)=>
      ImgReg1IN_275, F(2)=>ImgReg1IN_274, F(1)=>ImgReg1IN_273, F(0)=>
      ImgReg1IN_272);
   loop3_17_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_303_EXMPLR, D(14)=>OutputImg2_302_EXMPLR, D(13)=>
      OutputImg2_301_EXMPLR, D(12)=>OutputImg2_300_EXMPLR, D(11)=>
      OutputImg2_299_EXMPLR, D(10)=>OutputImg2_298_EXMPLR, D(9)=>
      OutputImg2_297_EXMPLR, D(8)=>OutputImg2_296_EXMPLR, D(7)=>
      OutputImg2_295_EXMPLR, D(6)=>OutputImg2_294_EXMPLR, D(5)=>
      OutputImg2_293_EXMPLR, D(4)=>OutputImg2_292_EXMPLR, D(3)=>
      OutputImg2_291_EXMPLR, D(2)=>OutputImg2_290_EXMPLR, D(1)=>
      OutputImg2_289_EXMPLR, D(0)=>OutputImg2_288_EXMPLR, EN=>nx23694, F(15)
      =>ImgReg2IN_287, F(14)=>ImgReg2IN_286, F(13)=>ImgReg2IN_285, F(12)=>
      ImgReg2IN_284, F(11)=>ImgReg2IN_283, F(10)=>ImgReg2IN_282, F(9)=>
      ImgReg2IN_281, F(8)=>ImgReg2IN_280, F(7)=>ImgReg2IN_279, F(6)=>
      ImgReg2IN_278, F(5)=>ImgReg2IN_277, F(4)=>ImgReg2IN_276, F(3)=>
      ImgReg2IN_275, F(2)=>ImgReg2IN_274, F(1)=>ImgReg2IN_273, F(0)=>
      ImgReg2IN_272);
   loop3_17_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_303_EXMPLR, D(14)=>OutputImg3_302_EXMPLR, D(13)=>
      OutputImg3_301_EXMPLR, D(12)=>OutputImg3_300_EXMPLR, D(11)=>
      OutputImg3_299_EXMPLR, D(10)=>OutputImg3_298_EXMPLR, D(9)=>
      OutputImg3_297_EXMPLR, D(8)=>OutputImg3_296_EXMPLR, D(7)=>
      OutputImg3_295_EXMPLR, D(6)=>OutputImg3_294_EXMPLR, D(5)=>
      OutputImg3_293_EXMPLR, D(4)=>OutputImg3_292_EXMPLR, D(3)=>
      OutputImg3_291_EXMPLR, D(2)=>OutputImg3_290_EXMPLR, D(1)=>
      OutputImg3_289_EXMPLR, D(0)=>OutputImg3_288_EXMPLR, EN=>nx23696, F(15)
      =>ImgReg3IN_287, F(14)=>ImgReg3IN_286, F(13)=>ImgReg3IN_285, F(12)=>
      ImgReg3IN_284, F(11)=>ImgReg3IN_283, F(10)=>ImgReg3IN_282, F(9)=>
      ImgReg3IN_281, F(8)=>ImgReg3IN_280, F(7)=>ImgReg3IN_279, F(6)=>
      ImgReg3IN_278, F(5)=>ImgReg3IN_277, F(4)=>ImgReg3IN_276, F(3)=>
      ImgReg3IN_275, F(2)=>ImgReg3IN_274, F(1)=>ImgReg3IN_273, F(0)=>
      ImgReg3IN_272);
   loop3_17_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_303_EXMPLR, D(14)=>OutputImg4_302_EXMPLR, D(13)=>
      OutputImg4_301_EXMPLR, D(12)=>OutputImg4_300_EXMPLR, D(11)=>
      OutputImg4_299_EXMPLR, D(10)=>OutputImg4_298_EXMPLR, D(9)=>
      OutputImg4_297_EXMPLR, D(8)=>OutputImg4_296_EXMPLR, D(7)=>
      OutputImg4_295_EXMPLR, D(6)=>OutputImg4_294_EXMPLR, D(5)=>
      OutputImg4_293_EXMPLR, D(4)=>OutputImg4_292_EXMPLR, D(3)=>
      OutputImg4_291_EXMPLR, D(2)=>OutputImg4_290_EXMPLR, D(1)=>
      OutputImg4_289_EXMPLR, D(0)=>OutputImg4_288_EXMPLR, EN=>nx23696, F(15)
      =>ImgReg4IN_287, F(14)=>ImgReg4IN_286, F(13)=>ImgReg4IN_285, F(12)=>
      ImgReg4IN_284, F(11)=>ImgReg4IN_283, F(10)=>ImgReg4IN_282, F(9)=>
      ImgReg4IN_281, F(8)=>ImgReg4IN_280, F(7)=>ImgReg4IN_279, F(6)=>
      ImgReg4IN_278, F(5)=>ImgReg4IN_277, F(4)=>ImgReg4IN_276, F(3)=>
      ImgReg4IN_275, F(2)=>ImgReg4IN_274, F(1)=>ImgReg4IN_273, F(0)=>
      ImgReg4IN_272);
   loop3_17_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_303_EXMPLR, D(14)=>OutputImg5_302_EXMPLR, D(13)=>
      OutputImg5_301_EXMPLR, D(12)=>OutputImg5_300_EXMPLR, D(11)=>
      OutputImg5_299_EXMPLR, D(10)=>OutputImg5_298_EXMPLR, D(9)=>
      OutputImg5_297_EXMPLR, D(8)=>OutputImg5_296_EXMPLR, D(7)=>
      OutputImg5_295_EXMPLR, D(6)=>OutputImg5_294_EXMPLR, D(5)=>
      OutputImg5_293_EXMPLR, D(4)=>OutputImg5_292_EXMPLR, D(3)=>
      OutputImg5_291_EXMPLR, D(2)=>OutputImg5_290_EXMPLR, D(1)=>
      OutputImg5_289_EXMPLR, D(0)=>OutputImg5_288_EXMPLR, EN=>nx23696, F(15)
      =>ImgReg5IN_287, F(14)=>ImgReg5IN_286, F(13)=>ImgReg5IN_285, F(12)=>
      ImgReg5IN_284, F(11)=>ImgReg5IN_283, F(10)=>ImgReg5IN_282, F(9)=>
      ImgReg5IN_281, F(8)=>ImgReg5IN_280, F(7)=>ImgReg5IN_279, F(6)=>
      ImgReg5IN_278, F(5)=>ImgReg5IN_277, F(4)=>ImgReg5IN_276, F(3)=>
      ImgReg5IN_275, F(2)=>ImgReg5IN_274, F(1)=>ImgReg5IN_273, F(0)=>
      ImgReg5IN_272);
   loop3_17_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(287), 
      D(14)=>DATA(286), D(13)=>DATA(285), D(12)=>DATA(284), D(11)=>DATA(283), 
      D(10)=>DATA(282), D(9)=>DATA(281), D(8)=>DATA(280), D(7)=>DATA(279), 
      D(6)=>DATA(278), D(5)=>DATA(277), D(4)=>DATA(276), D(3)=>DATA(275), 
      D(2)=>DATA(274), D(1)=>DATA(273), D(0)=>DATA(272), EN=>nx23658, F(15)
      =>ImgReg0IN_287, F(14)=>ImgReg0IN_286, F(13)=>ImgReg0IN_285, F(12)=>
      ImgReg0IN_284, F(11)=>ImgReg0IN_283, F(10)=>ImgReg0IN_282, F(9)=>
      ImgReg0IN_281, F(8)=>ImgReg0IN_280, F(7)=>ImgReg0IN_279, F(6)=>
      ImgReg0IN_278, F(5)=>ImgReg0IN_277, F(4)=>ImgReg0IN_276, F(3)=>
      ImgReg0IN_275, F(2)=>ImgReg0IN_274, F(1)=>ImgReg0IN_273, F(0)=>
      ImgReg0IN_272);
   loop3_17_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(287), 
      D(14)=>DATA(286), D(13)=>DATA(285), D(12)=>DATA(284), D(11)=>DATA(283), 
      D(10)=>DATA(282), D(9)=>DATA(281), D(8)=>DATA(280), D(7)=>DATA(279), 
      D(6)=>DATA(278), D(5)=>DATA(277), D(4)=>DATA(276), D(3)=>DATA(275), 
      D(2)=>DATA(274), D(1)=>DATA(273), D(0)=>DATA(272), EN=>nx23646, F(15)
      =>ImgReg1IN_287, F(14)=>ImgReg1IN_286, F(13)=>ImgReg1IN_285, F(12)=>
      ImgReg1IN_284, F(11)=>ImgReg1IN_283, F(10)=>ImgReg1IN_282, F(9)=>
      ImgReg1IN_281, F(8)=>ImgReg1IN_280, F(7)=>ImgReg1IN_279, F(6)=>
      ImgReg1IN_278, F(5)=>ImgReg1IN_277, F(4)=>ImgReg1IN_276, F(3)=>
      ImgReg1IN_275, F(2)=>ImgReg1IN_274, F(1)=>ImgReg1IN_273, F(0)=>
      ImgReg1IN_272);
   loop3_17_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(287), 
      D(14)=>DATA(286), D(13)=>DATA(285), D(12)=>DATA(284), D(11)=>DATA(283), 
      D(10)=>DATA(282), D(9)=>DATA(281), D(8)=>DATA(280), D(7)=>DATA(279), 
      D(6)=>DATA(278), D(5)=>DATA(277), D(4)=>DATA(276), D(3)=>DATA(275), 
      D(2)=>DATA(274), D(1)=>DATA(273), D(0)=>DATA(272), EN=>nx23634, F(15)
      =>ImgReg2IN_287, F(14)=>ImgReg2IN_286, F(13)=>ImgReg2IN_285, F(12)=>
      ImgReg2IN_284, F(11)=>ImgReg2IN_283, F(10)=>ImgReg2IN_282, F(9)=>
      ImgReg2IN_281, F(8)=>ImgReg2IN_280, F(7)=>ImgReg2IN_279, F(6)=>
      ImgReg2IN_278, F(5)=>ImgReg2IN_277, F(4)=>ImgReg2IN_276, F(3)=>
      ImgReg2IN_275, F(2)=>ImgReg2IN_274, F(1)=>ImgReg2IN_273, F(0)=>
      ImgReg2IN_272);
   loop3_17_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(287), 
      D(14)=>DATA(286), D(13)=>DATA(285), D(12)=>DATA(284), D(11)=>DATA(283), 
      D(10)=>DATA(282), D(9)=>DATA(281), D(8)=>DATA(280), D(7)=>DATA(279), 
      D(6)=>DATA(278), D(5)=>DATA(277), D(4)=>DATA(276), D(3)=>DATA(275), 
      D(2)=>DATA(274), D(1)=>DATA(273), D(0)=>DATA(272), EN=>nx23622, F(15)
      =>ImgReg3IN_287, F(14)=>ImgReg3IN_286, F(13)=>ImgReg3IN_285, F(12)=>
      ImgReg3IN_284, F(11)=>ImgReg3IN_283, F(10)=>ImgReg3IN_282, F(9)=>
      ImgReg3IN_281, F(8)=>ImgReg3IN_280, F(7)=>ImgReg3IN_279, F(6)=>
      ImgReg3IN_278, F(5)=>ImgReg3IN_277, F(4)=>ImgReg3IN_276, F(3)=>
      ImgReg3IN_275, F(2)=>ImgReg3IN_274, F(1)=>ImgReg3IN_273, F(0)=>
      ImgReg3IN_272);
   loop3_17_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(287), 
      D(14)=>DATA(286), D(13)=>DATA(285), D(12)=>DATA(284), D(11)=>DATA(283), 
      D(10)=>DATA(282), D(9)=>DATA(281), D(8)=>DATA(280), D(7)=>DATA(279), 
      D(6)=>DATA(278), D(5)=>DATA(277), D(4)=>DATA(276), D(3)=>DATA(275), 
      D(2)=>DATA(274), D(1)=>DATA(273), D(0)=>DATA(272), EN=>nx23610, F(15)
      =>ImgReg4IN_287, F(14)=>ImgReg4IN_286, F(13)=>ImgReg4IN_285, F(12)=>
      ImgReg4IN_284, F(11)=>ImgReg4IN_283, F(10)=>ImgReg4IN_282, F(9)=>
      ImgReg4IN_281, F(8)=>ImgReg4IN_280, F(7)=>ImgReg4IN_279, F(6)=>
      ImgReg4IN_278, F(5)=>ImgReg4IN_277, F(4)=>ImgReg4IN_276, F(3)=>
      ImgReg4IN_275, F(2)=>ImgReg4IN_274, F(1)=>ImgReg4IN_273, F(0)=>
      ImgReg4IN_272);
   loop3_17_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(287), 
      D(14)=>DATA(286), D(13)=>DATA(285), D(12)=>DATA(284), D(11)=>DATA(283), 
      D(10)=>DATA(282), D(9)=>DATA(281), D(8)=>DATA(280), D(7)=>DATA(279), 
      D(6)=>DATA(278), D(5)=>DATA(277), D(4)=>DATA(276), D(3)=>DATA(275), 
      D(2)=>DATA(274), D(1)=>DATA(273), D(0)=>DATA(272), EN=>nx23598, F(15)
      =>ImgReg5IN_287, F(14)=>ImgReg5IN_286, F(13)=>ImgReg5IN_285, F(12)=>
      ImgReg5IN_284, F(11)=>ImgReg5IN_283, F(10)=>ImgReg5IN_282, F(9)=>
      ImgReg5IN_281, F(8)=>ImgReg5IN_280, F(7)=>ImgReg5IN_279, F(6)=>
      ImgReg5IN_278, F(5)=>ImgReg5IN_277, F(4)=>ImgReg5IN_276, F(3)=>
      ImgReg5IN_275, F(2)=>ImgReg5IN_274, F(1)=>ImgReg5IN_273, F(0)=>
      ImgReg5IN_272);
   loop3_17_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_287_EXMPLR, D(14)=>OutputImg1_286_EXMPLR, D(13)=>
      OutputImg1_285_EXMPLR, D(12)=>OutputImg1_284_EXMPLR, D(11)=>
      OutputImg1_283_EXMPLR, D(10)=>OutputImg1_282_EXMPLR, D(9)=>
      OutputImg1_281_EXMPLR, D(8)=>OutputImg1_280_EXMPLR, D(7)=>
      OutputImg1_279_EXMPLR, D(6)=>OutputImg1_278_EXMPLR, D(5)=>
      OutputImg1_277_EXMPLR, D(4)=>OutputImg1_276_EXMPLR, D(3)=>
      OutputImg1_275_EXMPLR, D(2)=>OutputImg1_274_EXMPLR, D(1)=>
      OutputImg1_273_EXMPLR, D(0)=>OutputImg1_272_EXMPLR, EN=>nx23810, F(15)
      =>ImgReg0IN_287, F(14)=>ImgReg0IN_286, F(13)=>ImgReg0IN_285, F(12)=>
      ImgReg0IN_284, F(11)=>ImgReg0IN_283, F(10)=>ImgReg0IN_282, F(9)=>
      ImgReg0IN_281, F(8)=>ImgReg0IN_280, F(7)=>ImgReg0IN_279, F(6)=>
      ImgReg0IN_278, F(5)=>ImgReg0IN_277, F(4)=>ImgReg0IN_276, F(3)=>
      ImgReg0IN_275, F(2)=>ImgReg0IN_274, F(1)=>ImgReg0IN_273, F(0)=>
      ImgReg0IN_272);
   loop3_17_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_287_EXMPLR, D(14)=>OutputImg2_286_EXMPLR, D(13)=>
      OutputImg2_285_EXMPLR, D(12)=>OutputImg2_284_EXMPLR, D(11)=>
      OutputImg2_283_EXMPLR, D(10)=>OutputImg2_282_EXMPLR, D(9)=>
      OutputImg2_281_EXMPLR, D(8)=>OutputImg2_280_EXMPLR, D(7)=>
      OutputImg2_279_EXMPLR, D(6)=>OutputImg2_278_EXMPLR, D(5)=>
      OutputImg2_277_EXMPLR, D(4)=>OutputImg2_276_EXMPLR, D(3)=>
      OutputImg2_275_EXMPLR, D(2)=>OutputImg2_274_EXMPLR, D(1)=>
      OutputImg2_273_EXMPLR, D(0)=>OutputImg2_272_EXMPLR, EN=>nx23810, F(15)
      =>ImgReg1IN_287, F(14)=>ImgReg1IN_286, F(13)=>ImgReg1IN_285, F(12)=>
      ImgReg1IN_284, F(11)=>ImgReg1IN_283, F(10)=>ImgReg1IN_282, F(9)=>
      ImgReg1IN_281, F(8)=>ImgReg1IN_280, F(7)=>ImgReg1IN_279, F(6)=>
      ImgReg1IN_278, F(5)=>ImgReg1IN_277, F(4)=>ImgReg1IN_276, F(3)=>
      ImgReg1IN_275, F(2)=>ImgReg1IN_274, F(1)=>ImgReg1IN_273, F(0)=>
      ImgReg1IN_272);
   loop3_17_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_287_EXMPLR, D(14)=>OutputImg3_286_EXMPLR, D(13)=>
      OutputImg3_285_EXMPLR, D(12)=>OutputImg3_284_EXMPLR, D(11)=>
      OutputImg3_283_EXMPLR, D(10)=>OutputImg3_282_EXMPLR, D(9)=>
      OutputImg3_281_EXMPLR, D(8)=>OutputImg3_280_EXMPLR, D(7)=>
      OutputImg3_279_EXMPLR, D(6)=>OutputImg3_278_EXMPLR, D(5)=>
      OutputImg3_277_EXMPLR, D(4)=>OutputImg3_276_EXMPLR, D(3)=>
      OutputImg3_275_EXMPLR, D(2)=>OutputImg3_274_EXMPLR, D(1)=>
      OutputImg3_273_EXMPLR, D(0)=>OutputImg3_272_EXMPLR, EN=>nx23810, F(15)
      =>ImgReg2IN_287, F(14)=>ImgReg2IN_286, F(13)=>ImgReg2IN_285, F(12)=>
      ImgReg2IN_284, F(11)=>ImgReg2IN_283, F(10)=>ImgReg2IN_282, F(9)=>
      ImgReg2IN_281, F(8)=>ImgReg2IN_280, F(7)=>ImgReg2IN_279, F(6)=>
      ImgReg2IN_278, F(5)=>ImgReg2IN_277, F(4)=>ImgReg2IN_276, F(3)=>
      ImgReg2IN_275, F(2)=>ImgReg2IN_274, F(1)=>ImgReg2IN_273, F(0)=>
      ImgReg2IN_272);
   loop3_17_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_287_EXMPLR, D(14)=>OutputImg4_286_EXMPLR, D(13)=>
      OutputImg4_285_EXMPLR, D(12)=>OutputImg4_284_EXMPLR, D(11)=>
      OutputImg4_283_EXMPLR, D(10)=>OutputImg4_282_EXMPLR, D(9)=>
      OutputImg4_281_EXMPLR, D(8)=>OutputImg4_280_EXMPLR, D(7)=>
      OutputImg4_279_EXMPLR, D(6)=>OutputImg4_278_EXMPLR, D(5)=>
      OutputImg4_277_EXMPLR, D(4)=>OutputImg4_276_EXMPLR, D(3)=>
      OutputImg4_275_EXMPLR, D(2)=>OutputImg4_274_EXMPLR, D(1)=>
      OutputImg4_273_EXMPLR, D(0)=>OutputImg4_272_EXMPLR, EN=>nx23810, F(15)
      =>ImgReg3IN_287, F(14)=>ImgReg3IN_286, F(13)=>ImgReg3IN_285, F(12)=>
      ImgReg3IN_284, F(11)=>ImgReg3IN_283, F(10)=>ImgReg3IN_282, F(9)=>
      ImgReg3IN_281, F(8)=>ImgReg3IN_280, F(7)=>ImgReg3IN_279, F(6)=>
      ImgReg3IN_278, F(5)=>ImgReg3IN_277, F(4)=>ImgReg3IN_276, F(3)=>
      ImgReg3IN_275, F(2)=>ImgReg3IN_274, F(1)=>ImgReg3IN_273, F(0)=>
      ImgReg3IN_272);
   loop3_17_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_287_EXMPLR, D(14)=>OutputImg5_286_EXMPLR, D(13)=>
      OutputImg5_285_EXMPLR, D(12)=>OutputImg5_284_EXMPLR, D(11)=>
      OutputImg5_283_EXMPLR, D(10)=>OutputImg5_282_EXMPLR, D(9)=>
      OutputImg5_281_EXMPLR, D(8)=>OutputImg5_280_EXMPLR, D(7)=>
      OutputImg5_279_EXMPLR, D(6)=>OutputImg5_278_EXMPLR, D(5)=>
      OutputImg5_277_EXMPLR, D(4)=>OutputImg5_276_EXMPLR, D(3)=>
      OutputImg5_275_EXMPLR, D(2)=>OutputImg5_274_EXMPLR, D(1)=>
      OutputImg5_273_EXMPLR, D(0)=>OutputImg5_272_EXMPLR, EN=>nx23810, F(15)
      =>ImgReg4IN_287, F(14)=>ImgReg4IN_286, F(13)=>ImgReg4IN_285, F(12)=>
      ImgReg4IN_284, F(11)=>ImgReg4IN_283, F(10)=>ImgReg4IN_282, F(9)=>
      ImgReg4IN_281, F(8)=>ImgReg4IN_280, F(7)=>ImgReg4IN_279, F(6)=>
      ImgReg4IN_278, F(5)=>ImgReg4IN_277, F(4)=>ImgReg4IN_276, F(3)=>
      ImgReg4IN_275, F(2)=>ImgReg4IN_274, F(1)=>ImgReg4IN_273, F(0)=>
      ImgReg4IN_272);
   loop3_17_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_287, D(14)=>
      ImgReg0IN_286, D(13)=>ImgReg0IN_285, D(12)=>ImgReg0IN_284, D(11)=>
      ImgReg0IN_283, D(10)=>ImgReg0IN_282, D(9)=>ImgReg0IN_281, D(8)=>
      ImgReg0IN_280, D(7)=>ImgReg0IN_279, D(6)=>ImgReg0IN_278, D(5)=>
      ImgReg0IN_277, D(4)=>ImgReg0IN_276, D(3)=>ImgReg0IN_275, D(2)=>
      ImgReg0IN_274, D(1)=>ImgReg0IN_273, D(0)=>ImgReg0IN_272, CLK=>nx23930, 
      RST=>RST, EN=>nx23722, Q(15)=>OutputImg0_287_EXMPLR, Q(14)=>
      OutputImg0_286_EXMPLR, Q(13)=>OutputImg0_285_EXMPLR, Q(12)=>
      OutputImg0_284_EXMPLR, Q(11)=>OutputImg0_283_EXMPLR, Q(10)=>
      OutputImg0_282_EXMPLR, Q(9)=>OutputImg0_281_EXMPLR, Q(8)=>
      OutputImg0_280_EXMPLR, Q(7)=>OutputImg0_279_EXMPLR, Q(6)=>
      OutputImg0_278_EXMPLR, Q(5)=>OutputImg0_277_EXMPLR, Q(4)=>
      OutputImg0_276_EXMPLR, Q(3)=>OutputImg0_275_EXMPLR, Q(2)=>
      OutputImg0_274_EXMPLR, Q(1)=>OutputImg0_273_EXMPLR, Q(0)=>
      OutputImg0_272_EXMPLR);
   loop3_17_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_287, D(14)=>
      ImgReg1IN_286, D(13)=>ImgReg1IN_285, D(12)=>ImgReg1IN_284, D(11)=>
      ImgReg1IN_283, D(10)=>ImgReg1IN_282, D(9)=>ImgReg1IN_281, D(8)=>
      ImgReg1IN_280, D(7)=>ImgReg1IN_279, D(6)=>ImgReg1IN_278, D(5)=>
      ImgReg1IN_277, D(4)=>ImgReg1IN_276, D(3)=>ImgReg1IN_275, D(2)=>
      ImgReg1IN_274, D(1)=>ImgReg1IN_273, D(0)=>ImgReg1IN_272, CLK=>nx23932, 
      RST=>RST, EN=>nx23732, Q(15)=>OutputImg1_287_EXMPLR, Q(14)=>
      OutputImg1_286_EXMPLR, Q(13)=>OutputImg1_285_EXMPLR, Q(12)=>
      OutputImg1_284_EXMPLR, Q(11)=>OutputImg1_283_EXMPLR, Q(10)=>
      OutputImg1_282_EXMPLR, Q(9)=>OutputImg1_281_EXMPLR, Q(8)=>
      OutputImg1_280_EXMPLR, Q(7)=>OutputImg1_279_EXMPLR, Q(6)=>
      OutputImg1_278_EXMPLR, Q(5)=>OutputImg1_277_EXMPLR, Q(4)=>
      OutputImg1_276_EXMPLR, Q(3)=>OutputImg1_275_EXMPLR, Q(2)=>
      OutputImg1_274_EXMPLR, Q(1)=>OutputImg1_273_EXMPLR, Q(0)=>
      OutputImg1_272_EXMPLR);
   loop3_17_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_287, D(14)=>
      ImgReg2IN_286, D(13)=>ImgReg2IN_285, D(12)=>ImgReg2IN_284, D(11)=>
      ImgReg2IN_283, D(10)=>ImgReg2IN_282, D(9)=>ImgReg2IN_281, D(8)=>
      ImgReg2IN_280, D(7)=>ImgReg2IN_279, D(6)=>ImgReg2IN_278, D(5)=>
      ImgReg2IN_277, D(4)=>ImgReg2IN_276, D(3)=>ImgReg2IN_275, D(2)=>
      ImgReg2IN_274, D(1)=>ImgReg2IN_273, D(0)=>ImgReg2IN_272, CLK=>nx23932, 
      RST=>RST, EN=>nx23742, Q(15)=>OutputImg2_287_EXMPLR, Q(14)=>
      OutputImg2_286_EXMPLR, Q(13)=>OutputImg2_285_EXMPLR, Q(12)=>
      OutputImg2_284_EXMPLR, Q(11)=>OutputImg2_283_EXMPLR, Q(10)=>
      OutputImg2_282_EXMPLR, Q(9)=>OutputImg2_281_EXMPLR, Q(8)=>
      OutputImg2_280_EXMPLR, Q(7)=>OutputImg2_279_EXMPLR, Q(6)=>
      OutputImg2_278_EXMPLR, Q(5)=>OutputImg2_277_EXMPLR, Q(4)=>
      OutputImg2_276_EXMPLR, Q(3)=>OutputImg2_275_EXMPLR, Q(2)=>
      OutputImg2_274_EXMPLR, Q(1)=>OutputImg2_273_EXMPLR, Q(0)=>
      OutputImg2_272_EXMPLR);
   loop3_17_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_287, D(14)=>
      ImgReg3IN_286, D(13)=>ImgReg3IN_285, D(12)=>ImgReg3IN_284, D(11)=>
      ImgReg3IN_283, D(10)=>ImgReg3IN_282, D(9)=>ImgReg3IN_281, D(8)=>
      ImgReg3IN_280, D(7)=>ImgReg3IN_279, D(6)=>ImgReg3IN_278, D(5)=>
      ImgReg3IN_277, D(4)=>ImgReg3IN_276, D(3)=>ImgReg3IN_275, D(2)=>
      ImgReg3IN_274, D(1)=>ImgReg3IN_273, D(0)=>ImgReg3IN_272, CLK=>nx23934, 
      RST=>RST, EN=>nx23752, Q(15)=>OutputImg3_287_EXMPLR, Q(14)=>
      OutputImg3_286_EXMPLR, Q(13)=>OutputImg3_285_EXMPLR, Q(12)=>
      OutputImg3_284_EXMPLR, Q(11)=>OutputImg3_283_EXMPLR, Q(10)=>
      OutputImg3_282_EXMPLR, Q(9)=>OutputImg3_281_EXMPLR, Q(8)=>
      OutputImg3_280_EXMPLR, Q(7)=>OutputImg3_279_EXMPLR, Q(6)=>
      OutputImg3_278_EXMPLR, Q(5)=>OutputImg3_277_EXMPLR, Q(4)=>
      OutputImg3_276_EXMPLR, Q(3)=>OutputImg3_275_EXMPLR, Q(2)=>
      OutputImg3_274_EXMPLR, Q(1)=>OutputImg3_273_EXMPLR, Q(0)=>
      OutputImg3_272_EXMPLR);
   loop3_17_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_287, D(14)=>
      ImgReg4IN_286, D(13)=>ImgReg4IN_285, D(12)=>ImgReg4IN_284, D(11)=>
      ImgReg4IN_283, D(10)=>ImgReg4IN_282, D(9)=>ImgReg4IN_281, D(8)=>
      ImgReg4IN_280, D(7)=>ImgReg4IN_279, D(6)=>ImgReg4IN_278, D(5)=>
      ImgReg4IN_277, D(4)=>ImgReg4IN_276, D(3)=>ImgReg4IN_275, D(2)=>
      ImgReg4IN_274, D(1)=>ImgReg4IN_273, D(0)=>ImgReg4IN_272, CLK=>nx23934, 
      RST=>RST, EN=>nx23762, Q(15)=>OutputImg4_287_EXMPLR, Q(14)=>
      OutputImg4_286_EXMPLR, Q(13)=>OutputImg4_285_EXMPLR, Q(12)=>
      OutputImg4_284_EXMPLR, Q(11)=>OutputImg4_283_EXMPLR, Q(10)=>
      OutputImg4_282_EXMPLR, Q(9)=>OutputImg4_281_EXMPLR, Q(8)=>
      OutputImg4_280_EXMPLR, Q(7)=>OutputImg4_279_EXMPLR, Q(6)=>
      OutputImg4_278_EXMPLR, Q(5)=>OutputImg4_277_EXMPLR, Q(4)=>
      OutputImg4_276_EXMPLR, Q(3)=>OutputImg4_275_EXMPLR, Q(2)=>
      OutputImg4_274_EXMPLR, Q(1)=>OutputImg4_273_EXMPLR, Q(0)=>
      OutputImg4_272_EXMPLR);
   loop3_17_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_287, D(14)=>
      ImgReg5IN_286, D(13)=>ImgReg5IN_285, D(12)=>ImgReg5IN_284, D(11)=>
      ImgReg5IN_283, D(10)=>ImgReg5IN_282, D(9)=>ImgReg5IN_281, D(8)=>
      ImgReg5IN_280, D(7)=>ImgReg5IN_279, D(6)=>ImgReg5IN_278, D(5)=>
      ImgReg5IN_277, D(4)=>ImgReg5IN_276, D(3)=>ImgReg5IN_275, D(2)=>
      ImgReg5IN_274, D(1)=>ImgReg5IN_273, D(0)=>ImgReg5IN_272, CLK=>nx23936, 
      RST=>RST, EN=>nx23772, Q(15)=>OutputImg5_287_EXMPLR, Q(14)=>
      OutputImg5_286_EXMPLR, Q(13)=>OutputImg5_285_EXMPLR, Q(12)=>
      OutputImg5_284_EXMPLR, Q(11)=>OutputImg5_283_EXMPLR, Q(10)=>
      OutputImg5_282_EXMPLR, Q(9)=>OutputImg5_281_EXMPLR, Q(8)=>
      OutputImg5_280_EXMPLR, Q(7)=>OutputImg5_279_EXMPLR, Q(6)=>
      OutputImg5_278_EXMPLR, Q(5)=>OutputImg5_277_EXMPLR, Q(4)=>
      OutputImg5_276_EXMPLR, Q(3)=>OutputImg5_275_EXMPLR, Q(2)=>
      OutputImg5_274_EXMPLR, Q(1)=>OutputImg5_273_EXMPLR, Q(0)=>
      OutputImg5_272_EXMPLR);
   loop3_18_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_319_EXMPLR, D(14)=>OutputImg0_318_EXMPLR, D(13)=>
      OutputImg0_317_EXMPLR, D(12)=>OutputImg0_316_EXMPLR, D(11)=>
      OutputImg0_315_EXMPLR, D(10)=>OutputImg0_314_EXMPLR, D(9)=>
      OutputImg0_313_EXMPLR, D(8)=>OutputImg0_312_EXMPLR, D(7)=>
      OutputImg0_311_EXMPLR, D(6)=>OutputImg0_310_EXMPLR, D(5)=>
      OutputImg0_309_EXMPLR, D(4)=>OutputImg0_308_EXMPLR, D(3)=>
      OutputImg0_307_EXMPLR, D(2)=>OutputImg0_306_EXMPLR, D(1)=>
      OutputImg0_305_EXMPLR, D(0)=>OutputImg0_304_EXMPLR, EN=>nx23696, F(15)
      =>ImgReg0IN_303, F(14)=>ImgReg0IN_302, F(13)=>ImgReg0IN_301, F(12)=>
      ImgReg0IN_300, F(11)=>ImgReg0IN_299, F(10)=>ImgReg0IN_298, F(9)=>
      ImgReg0IN_297, F(8)=>ImgReg0IN_296, F(7)=>ImgReg0IN_295, F(6)=>
      ImgReg0IN_294, F(5)=>ImgReg0IN_293, F(4)=>ImgReg0IN_292, F(3)=>
      ImgReg0IN_291, F(2)=>ImgReg0IN_290, F(1)=>ImgReg0IN_289, F(0)=>
      ImgReg0IN_288);
   loop3_18_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_319_EXMPLR, D(14)=>OutputImg1_318_EXMPLR, D(13)=>
      OutputImg1_317_EXMPLR, D(12)=>OutputImg1_316_EXMPLR, D(11)=>
      OutputImg1_315_EXMPLR, D(10)=>OutputImg1_314_EXMPLR, D(9)=>
      OutputImg1_313_EXMPLR, D(8)=>OutputImg1_312_EXMPLR, D(7)=>
      OutputImg1_311_EXMPLR, D(6)=>OutputImg1_310_EXMPLR, D(5)=>
      OutputImg1_309_EXMPLR, D(4)=>OutputImg1_308_EXMPLR, D(3)=>
      OutputImg1_307_EXMPLR, D(2)=>OutputImg1_306_EXMPLR, D(1)=>
      OutputImg1_305_EXMPLR, D(0)=>OutputImg1_304_EXMPLR, EN=>nx23696, F(15)
      =>ImgReg1IN_303, F(14)=>ImgReg1IN_302, F(13)=>ImgReg1IN_301, F(12)=>
      ImgReg1IN_300, F(11)=>ImgReg1IN_299, F(10)=>ImgReg1IN_298, F(9)=>
      ImgReg1IN_297, F(8)=>ImgReg1IN_296, F(7)=>ImgReg1IN_295, F(6)=>
      ImgReg1IN_294, F(5)=>ImgReg1IN_293, F(4)=>ImgReg1IN_292, F(3)=>
      ImgReg1IN_291, F(2)=>ImgReg1IN_290, F(1)=>ImgReg1IN_289, F(0)=>
      ImgReg1IN_288);
   loop3_18_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_319_EXMPLR, D(14)=>OutputImg2_318_EXMPLR, D(13)=>
      OutputImg2_317_EXMPLR, D(12)=>OutputImg2_316_EXMPLR, D(11)=>
      OutputImg2_315_EXMPLR, D(10)=>OutputImg2_314_EXMPLR, D(9)=>
      OutputImg2_313_EXMPLR, D(8)=>OutputImg2_312_EXMPLR, D(7)=>
      OutputImg2_311_EXMPLR, D(6)=>OutputImg2_310_EXMPLR, D(5)=>
      OutputImg2_309_EXMPLR, D(4)=>OutputImg2_308_EXMPLR, D(3)=>
      OutputImg2_307_EXMPLR, D(2)=>OutputImg2_306_EXMPLR, D(1)=>
      OutputImg2_305_EXMPLR, D(0)=>OutputImg2_304_EXMPLR, EN=>nx23696, F(15)
      =>ImgReg2IN_303, F(14)=>ImgReg2IN_302, F(13)=>ImgReg2IN_301, F(12)=>
      ImgReg2IN_300, F(11)=>ImgReg2IN_299, F(10)=>ImgReg2IN_298, F(9)=>
      ImgReg2IN_297, F(8)=>ImgReg2IN_296, F(7)=>ImgReg2IN_295, F(6)=>
      ImgReg2IN_294, F(5)=>ImgReg2IN_293, F(4)=>ImgReg2IN_292, F(3)=>
      ImgReg2IN_291, F(2)=>ImgReg2IN_290, F(1)=>ImgReg2IN_289, F(0)=>
      ImgReg2IN_288);
   loop3_18_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_319_EXMPLR, D(14)=>OutputImg3_318_EXMPLR, D(13)=>
      OutputImg3_317_EXMPLR, D(12)=>OutputImg3_316_EXMPLR, D(11)=>
      OutputImg3_315_EXMPLR, D(10)=>OutputImg3_314_EXMPLR, D(9)=>
      OutputImg3_313_EXMPLR, D(8)=>OutputImg3_312_EXMPLR, D(7)=>
      OutputImg3_311_EXMPLR, D(6)=>OutputImg3_310_EXMPLR, D(5)=>
      OutputImg3_309_EXMPLR, D(4)=>OutputImg3_308_EXMPLR, D(3)=>
      OutputImg3_307_EXMPLR, D(2)=>OutputImg3_306_EXMPLR, D(1)=>
      OutputImg3_305_EXMPLR, D(0)=>OutputImg3_304_EXMPLR, EN=>nx23696, F(15)
      =>ImgReg3IN_303, F(14)=>ImgReg3IN_302, F(13)=>ImgReg3IN_301, F(12)=>
      ImgReg3IN_300, F(11)=>ImgReg3IN_299, F(10)=>ImgReg3IN_298, F(9)=>
      ImgReg3IN_297, F(8)=>ImgReg3IN_296, F(7)=>ImgReg3IN_295, F(6)=>
      ImgReg3IN_294, F(5)=>ImgReg3IN_293, F(4)=>ImgReg3IN_292, F(3)=>
      ImgReg3IN_291, F(2)=>ImgReg3IN_290, F(1)=>ImgReg3IN_289, F(0)=>
      ImgReg3IN_288);
   loop3_18_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_319_EXMPLR, D(14)=>OutputImg4_318_EXMPLR, D(13)=>
      OutputImg4_317_EXMPLR, D(12)=>OutputImg4_316_EXMPLR, D(11)=>
      OutputImg4_315_EXMPLR, D(10)=>OutputImg4_314_EXMPLR, D(9)=>
      OutputImg4_313_EXMPLR, D(8)=>OutputImg4_312_EXMPLR, D(7)=>
      OutputImg4_311_EXMPLR, D(6)=>OutputImg4_310_EXMPLR, D(5)=>
      OutputImg4_309_EXMPLR, D(4)=>OutputImg4_308_EXMPLR, D(3)=>
      OutputImg4_307_EXMPLR, D(2)=>OutputImg4_306_EXMPLR, D(1)=>
      OutputImg4_305_EXMPLR, D(0)=>OutputImg4_304_EXMPLR, EN=>nx23698, F(15)
      =>ImgReg4IN_303, F(14)=>ImgReg4IN_302, F(13)=>ImgReg4IN_301, F(12)=>
      ImgReg4IN_300, F(11)=>ImgReg4IN_299, F(10)=>ImgReg4IN_298, F(9)=>
      ImgReg4IN_297, F(8)=>ImgReg4IN_296, F(7)=>ImgReg4IN_295, F(6)=>
      ImgReg4IN_294, F(5)=>ImgReg4IN_293, F(4)=>ImgReg4IN_292, F(3)=>
      ImgReg4IN_291, F(2)=>ImgReg4IN_290, F(1)=>ImgReg4IN_289, F(0)=>
      ImgReg4IN_288);
   loop3_18_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_319_EXMPLR, D(14)=>OutputImg5_318_EXMPLR, D(13)=>
      OutputImg5_317_EXMPLR, D(12)=>OutputImg5_316_EXMPLR, D(11)=>
      OutputImg5_315_EXMPLR, D(10)=>OutputImg5_314_EXMPLR, D(9)=>
      OutputImg5_313_EXMPLR, D(8)=>OutputImg5_312_EXMPLR, D(7)=>
      OutputImg5_311_EXMPLR, D(6)=>OutputImg5_310_EXMPLR, D(5)=>
      OutputImg5_309_EXMPLR, D(4)=>OutputImg5_308_EXMPLR, D(3)=>
      OutputImg5_307_EXMPLR, D(2)=>OutputImg5_306_EXMPLR, D(1)=>
      OutputImg5_305_EXMPLR, D(0)=>OutputImg5_304_EXMPLR, EN=>nx23698, F(15)
      =>ImgReg5IN_303, F(14)=>ImgReg5IN_302, F(13)=>ImgReg5IN_301, F(12)=>
      ImgReg5IN_300, F(11)=>ImgReg5IN_299, F(10)=>ImgReg5IN_298, F(9)=>
      ImgReg5IN_297, F(8)=>ImgReg5IN_296, F(7)=>ImgReg5IN_295, F(6)=>
      ImgReg5IN_294, F(5)=>ImgReg5IN_293, F(4)=>ImgReg5IN_292, F(3)=>
      ImgReg5IN_291, F(2)=>ImgReg5IN_290, F(1)=>ImgReg5IN_289, F(0)=>
      ImgReg5IN_288);
   loop3_18_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(303), 
      D(14)=>DATA(302), D(13)=>DATA(301), D(12)=>DATA(300), D(11)=>DATA(299), 
      D(10)=>DATA(298), D(9)=>DATA(297), D(8)=>DATA(296), D(7)=>DATA(295), 
      D(6)=>DATA(294), D(5)=>DATA(293), D(4)=>DATA(292), D(3)=>DATA(291), 
      D(2)=>DATA(290), D(1)=>DATA(289), D(0)=>DATA(288), EN=>nx23658, F(15)
      =>ImgReg0IN_303, F(14)=>ImgReg0IN_302, F(13)=>ImgReg0IN_301, F(12)=>
      ImgReg0IN_300, F(11)=>ImgReg0IN_299, F(10)=>ImgReg0IN_298, F(9)=>
      ImgReg0IN_297, F(8)=>ImgReg0IN_296, F(7)=>ImgReg0IN_295, F(6)=>
      ImgReg0IN_294, F(5)=>ImgReg0IN_293, F(4)=>ImgReg0IN_292, F(3)=>
      ImgReg0IN_291, F(2)=>ImgReg0IN_290, F(1)=>ImgReg0IN_289, F(0)=>
      ImgReg0IN_288);
   loop3_18_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(303), 
      D(14)=>DATA(302), D(13)=>DATA(301), D(12)=>DATA(300), D(11)=>DATA(299), 
      D(10)=>DATA(298), D(9)=>DATA(297), D(8)=>DATA(296), D(7)=>DATA(295), 
      D(6)=>DATA(294), D(5)=>DATA(293), D(4)=>DATA(292), D(3)=>DATA(291), 
      D(2)=>DATA(290), D(1)=>DATA(289), D(0)=>DATA(288), EN=>nx23646, F(15)
      =>ImgReg1IN_303, F(14)=>ImgReg1IN_302, F(13)=>ImgReg1IN_301, F(12)=>
      ImgReg1IN_300, F(11)=>ImgReg1IN_299, F(10)=>ImgReg1IN_298, F(9)=>
      ImgReg1IN_297, F(8)=>ImgReg1IN_296, F(7)=>ImgReg1IN_295, F(6)=>
      ImgReg1IN_294, F(5)=>ImgReg1IN_293, F(4)=>ImgReg1IN_292, F(3)=>
      ImgReg1IN_291, F(2)=>ImgReg1IN_290, F(1)=>ImgReg1IN_289, F(0)=>
      ImgReg1IN_288);
   loop3_18_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(303), 
      D(14)=>DATA(302), D(13)=>DATA(301), D(12)=>DATA(300), D(11)=>DATA(299), 
      D(10)=>DATA(298), D(9)=>DATA(297), D(8)=>DATA(296), D(7)=>DATA(295), 
      D(6)=>DATA(294), D(5)=>DATA(293), D(4)=>DATA(292), D(3)=>DATA(291), 
      D(2)=>DATA(290), D(1)=>DATA(289), D(0)=>DATA(288), EN=>nx23634, F(15)
      =>ImgReg2IN_303, F(14)=>ImgReg2IN_302, F(13)=>ImgReg2IN_301, F(12)=>
      ImgReg2IN_300, F(11)=>ImgReg2IN_299, F(10)=>ImgReg2IN_298, F(9)=>
      ImgReg2IN_297, F(8)=>ImgReg2IN_296, F(7)=>ImgReg2IN_295, F(6)=>
      ImgReg2IN_294, F(5)=>ImgReg2IN_293, F(4)=>ImgReg2IN_292, F(3)=>
      ImgReg2IN_291, F(2)=>ImgReg2IN_290, F(1)=>ImgReg2IN_289, F(0)=>
      ImgReg2IN_288);
   loop3_18_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(303), 
      D(14)=>DATA(302), D(13)=>DATA(301), D(12)=>DATA(300), D(11)=>DATA(299), 
      D(10)=>DATA(298), D(9)=>DATA(297), D(8)=>DATA(296), D(7)=>DATA(295), 
      D(6)=>DATA(294), D(5)=>DATA(293), D(4)=>DATA(292), D(3)=>DATA(291), 
      D(2)=>DATA(290), D(1)=>DATA(289), D(0)=>DATA(288), EN=>nx23622, F(15)
      =>ImgReg3IN_303, F(14)=>ImgReg3IN_302, F(13)=>ImgReg3IN_301, F(12)=>
      ImgReg3IN_300, F(11)=>ImgReg3IN_299, F(10)=>ImgReg3IN_298, F(9)=>
      ImgReg3IN_297, F(8)=>ImgReg3IN_296, F(7)=>ImgReg3IN_295, F(6)=>
      ImgReg3IN_294, F(5)=>ImgReg3IN_293, F(4)=>ImgReg3IN_292, F(3)=>
      ImgReg3IN_291, F(2)=>ImgReg3IN_290, F(1)=>ImgReg3IN_289, F(0)=>
      ImgReg3IN_288);
   loop3_18_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(303), 
      D(14)=>DATA(302), D(13)=>DATA(301), D(12)=>DATA(300), D(11)=>DATA(299), 
      D(10)=>DATA(298), D(9)=>DATA(297), D(8)=>DATA(296), D(7)=>DATA(295), 
      D(6)=>DATA(294), D(5)=>DATA(293), D(4)=>DATA(292), D(3)=>DATA(291), 
      D(2)=>DATA(290), D(1)=>DATA(289), D(0)=>DATA(288), EN=>nx23610, F(15)
      =>ImgReg4IN_303, F(14)=>ImgReg4IN_302, F(13)=>ImgReg4IN_301, F(12)=>
      ImgReg4IN_300, F(11)=>ImgReg4IN_299, F(10)=>ImgReg4IN_298, F(9)=>
      ImgReg4IN_297, F(8)=>ImgReg4IN_296, F(7)=>ImgReg4IN_295, F(6)=>
      ImgReg4IN_294, F(5)=>ImgReg4IN_293, F(4)=>ImgReg4IN_292, F(3)=>
      ImgReg4IN_291, F(2)=>ImgReg4IN_290, F(1)=>ImgReg4IN_289, F(0)=>
      ImgReg4IN_288);
   loop3_18_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(303), 
      D(14)=>DATA(302), D(13)=>DATA(301), D(12)=>DATA(300), D(11)=>DATA(299), 
      D(10)=>DATA(298), D(9)=>DATA(297), D(8)=>DATA(296), D(7)=>DATA(295), 
      D(6)=>DATA(294), D(5)=>DATA(293), D(4)=>DATA(292), D(3)=>DATA(291), 
      D(2)=>DATA(290), D(1)=>DATA(289), D(0)=>DATA(288), EN=>nx23598, F(15)
      =>ImgReg5IN_303, F(14)=>ImgReg5IN_302, F(13)=>ImgReg5IN_301, F(12)=>
      ImgReg5IN_300, F(11)=>ImgReg5IN_299, F(10)=>ImgReg5IN_298, F(9)=>
      ImgReg5IN_297, F(8)=>ImgReg5IN_296, F(7)=>ImgReg5IN_295, F(6)=>
      ImgReg5IN_294, F(5)=>ImgReg5IN_293, F(4)=>ImgReg5IN_292, F(3)=>
      ImgReg5IN_291, F(2)=>ImgReg5IN_290, F(1)=>ImgReg5IN_289, F(0)=>
      ImgReg5IN_288);
   loop3_18_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_303_EXMPLR, D(14)=>OutputImg1_302_EXMPLR, D(13)=>
      OutputImg1_301_EXMPLR, D(12)=>OutputImg1_300_EXMPLR, D(11)=>
      OutputImg1_299_EXMPLR, D(10)=>OutputImg1_298_EXMPLR, D(9)=>
      OutputImg1_297_EXMPLR, D(8)=>OutputImg1_296_EXMPLR, D(7)=>
      OutputImg1_295_EXMPLR, D(6)=>OutputImg1_294_EXMPLR, D(5)=>
      OutputImg1_293_EXMPLR, D(4)=>OutputImg1_292_EXMPLR, D(3)=>
      OutputImg1_291_EXMPLR, D(2)=>OutputImg1_290_EXMPLR, D(1)=>
      OutputImg1_289_EXMPLR, D(0)=>OutputImg1_288_EXMPLR, EN=>nx23810, F(15)
      =>ImgReg0IN_303, F(14)=>ImgReg0IN_302, F(13)=>ImgReg0IN_301, F(12)=>
      ImgReg0IN_300, F(11)=>ImgReg0IN_299, F(10)=>ImgReg0IN_298, F(9)=>
      ImgReg0IN_297, F(8)=>ImgReg0IN_296, F(7)=>ImgReg0IN_295, F(6)=>
      ImgReg0IN_294, F(5)=>ImgReg0IN_293, F(4)=>ImgReg0IN_292, F(3)=>
      ImgReg0IN_291, F(2)=>ImgReg0IN_290, F(1)=>ImgReg0IN_289, F(0)=>
      ImgReg0IN_288);
   loop3_18_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_303_EXMPLR, D(14)=>OutputImg2_302_EXMPLR, D(13)=>
      OutputImg2_301_EXMPLR, D(12)=>OutputImg2_300_EXMPLR, D(11)=>
      OutputImg2_299_EXMPLR, D(10)=>OutputImg2_298_EXMPLR, D(9)=>
      OutputImg2_297_EXMPLR, D(8)=>OutputImg2_296_EXMPLR, D(7)=>
      OutputImg2_295_EXMPLR, D(6)=>OutputImg2_294_EXMPLR, D(5)=>
      OutputImg2_293_EXMPLR, D(4)=>OutputImg2_292_EXMPLR, D(3)=>
      OutputImg2_291_EXMPLR, D(2)=>OutputImg2_290_EXMPLR, D(1)=>
      OutputImg2_289_EXMPLR, D(0)=>OutputImg2_288_EXMPLR, EN=>nx23812, F(15)
      =>ImgReg1IN_303, F(14)=>ImgReg1IN_302, F(13)=>ImgReg1IN_301, F(12)=>
      ImgReg1IN_300, F(11)=>ImgReg1IN_299, F(10)=>ImgReg1IN_298, F(9)=>
      ImgReg1IN_297, F(8)=>ImgReg1IN_296, F(7)=>ImgReg1IN_295, F(6)=>
      ImgReg1IN_294, F(5)=>ImgReg1IN_293, F(4)=>ImgReg1IN_292, F(3)=>
      ImgReg1IN_291, F(2)=>ImgReg1IN_290, F(1)=>ImgReg1IN_289, F(0)=>
      ImgReg1IN_288);
   loop3_18_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_303_EXMPLR, D(14)=>OutputImg3_302_EXMPLR, D(13)=>
      OutputImg3_301_EXMPLR, D(12)=>OutputImg3_300_EXMPLR, D(11)=>
      OutputImg3_299_EXMPLR, D(10)=>OutputImg3_298_EXMPLR, D(9)=>
      OutputImg3_297_EXMPLR, D(8)=>OutputImg3_296_EXMPLR, D(7)=>
      OutputImg3_295_EXMPLR, D(6)=>OutputImg3_294_EXMPLR, D(5)=>
      OutputImg3_293_EXMPLR, D(4)=>OutputImg3_292_EXMPLR, D(3)=>
      OutputImg3_291_EXMPLR, D(2)=>OutputImg3_290_EXMPLR, D(1)=>
      OutputImg3_289_EXMPLR, D(0)=>OutputImg3_288_EXMPLR, EN=>nx23812, F(15)
      =>ImgReg2IN_303, F(14)=>ImgReg2IN_302, F(13)=>ImgReg2IN_301, F(12)=>
      ImgReg2IN_300, F(11)=>ImgReg2IN_299, F(10)=>ImgReg2IN_298, F(9)=>
      ImgReg2IN_297, F(8)=>ImgReg2IN_296, F(7)=>ImgReg2IN_295, F(6)=>
      ImgReg2IN_294, F(5)=>ImgReg2IN_293, F(4)=>ImgReg2IN_292, F(3)=>
      ImgReg2IN_291, F(2)=>ImgReg2IN_290, F(1)=>ImgReg2IN_289, F(0)=>
      ImgReg2IN_288);
   loop3_18_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_303_EXMPLR, D(14)=>OutputImg4_302_EXMPLR, D(13)=>
      OutputImg4_301_EXMPLR, D(12)=>OutputImg4_300_EXMPLR, D(11)=>
      OutputImg4_299_EXMPLR, D(10)=>OutputImg4_298_EXMPLR, D(9)=>
      OutputImg4_297_EXMPLR, D(8)=>OutputImg4_296_EXMPLR, D(7)=>
      OutputImg4_295_EXMPLR, D(6)=>OutputImg4_294_EXMPLR, D(5)=>
      OutputImg4_293_EXMPLR, D(4)=>OutputImg4_292_EXMPLR, D(3)=>
      OutputImg4_291_EXMPLR, D(2)=>OutputImg4_290_EXMPLR, D(1)=>
      OutputImg4_289_EXMPLR, D(0)=>OutputImg4_288_EXMPLR, EN=>nx23812, F(15)
      =>ImgReg3IN_303, F(14)=>ImgReg3IN_302, F(13)=>ImgReg3IN_301, F(12)=>
      ImgReg3IN_300, F(11)=>ImgReg3IN_299, F(10)=>ImgReg3IN_298, F(9)=>
      ImgReg3IN_297, F(8)=>ImgReg3IN_296, F(7)=>ImgReg3IN_295, F(6)=>
      ImgReg3IN_294, F(5)=>ImgReg3IN_293, F(4)=>ImgReg3IN_292, F(3)=>
      ImgReg3IN_291, F(2)=>ImgReg3IN_290, F(1)=>ImgReg3IN_289, F(0)=>
      ImgReg3IN_288);
   loop3_18_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_303_EXMPLR, D(14)=>OutputImg5_302_EXMPLR, D(13)=>
      OutputImg5_301_EXMPLR, D(12)=>OutputImg5_300_EXMPLR, D(11)=>
      OutputImg5_299_EXMPLR, D(10)=>OutputImg5_298_EXMPLR, D(9)=>
      OutputImg5_297_EXMPLR, D(8)=>OutputImg5_296_EXMPLR, D(7)=>
      OutputImg5_295_EXMPLR, D(6)=>OutputImg5_294_EXMPLR, D(5)=>
      OutputImg5_293_EXMPLR, D(4)=>OutputImg5_292_EXMPLR, D(3)=>
      OutputImg5_291_EXMPLR, D(2)=>OutputImg5_290_EXMPLR, D(1)=>
      OutputImg5_289_EXMPLR, D(0)=>OutputImg5_288_EXMPLR, EN=>nx23812, F(15)
      =>ImgReg4IN_303, F(14)=>ImgReg4IN_302, F(13)=>ImgReg4IN_301, F(12)=>
      ImgReg4IN_300, F(11)=>ImgReg4IN_299, F(10)=>ImgReg4IN_298, F(9)=>
      ImgReg4IN_297, F(8)=>ImgReg4IN_296, F(7)=>ImgReg4IN_295, F(6)=>
      ImgReg4IN_294, F(5)=>ImgReg4IN_293, F(4)=>ImgReg4IN_292, F(3)=>
      ImgReg4IN_291, F(2)=>ImgReg4IN_290, F(1)=>ImgReg4IN_289, F(0)=>
      ImgReg4IN_288);
   loop3_18_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_303, D(14)=>
      ImgReg0IN_302, D(13)=>ImgReg0IN_301, D(12)=>ImgReg0IN_300, D(11)=>
      ImgReg0IN_299, D(10)=>ImgReg0IN_298, D(9)=>ImgReg0IN_297, D(8)=>
      ImgReg0IN_296, D(7)=>ImgReg0IN_295, D(6)=>ImgReg0IN_294, D(5)=>
      ImgReg0IN_293, D(4)=>ImgReg0IN_292, D(3)=>ImgReg0IN_291, D(2)=>
      ImgReg0IN_290, D(1)=>ImgReg0IN_289, D(0)=>ImgReg0IN_288, CLK=>nx23936, 
      RST=>RST, EN=>nx23722, Q(15)=>OutputImg0_303_EXMPLR, Q(14)=>
      OutputImg0_302_EXMPLR, Q(13)=>OutputImg0_301_EXMPLR, Q(12)=>
      OutputImg0_300_EXMPLR, Q(11)=>OutputImg0_299_EXMPLR, Q(10)=>
      OutputImg0_298_EXMPLR, Q(9)=>OutputImg0_297_EXMPLR, Q(8)=>
      OutputImg0_296_EXMPLR, Q(7)=>OutputImg0_295_EXMPLR, Q(6)=>
      OutputImg0_294_EXMPLR, Q(5)=>OutputImg0_293_EXMPLR, Q(4)=>
      OutputImg0_292_EXMPLR, Q(3)=>OutputImg0_291_EXMPLR, Q(2)=>
      OutputImg0_290_EXMPLR, Q(1)=>OutputImg0_289_EXMPLR, Q(0)=>
      OutputImg0_288_EXMPLR);
   loop3_18_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_303, D(14)=>
      ImgReg1IN_302, D(13)=>ImgReg1IN_301, D(12)=>ImgReg1IN_300, D(11)=>
      ImgReg1IN_299, D(10)=>ImgReg1IN_298, D(9)=>ImgReg1IN_297, D(8)=>
      ImgReg1IN_296, D(7)=>ImgReg1IN_295, D(6)=>ImgReg1IN_294, D(5)=>
      ImgReg1IN_293, D(4)=>ImgReg1IN_292, D(3)=>ImgReg1IN_291, D(2)=>
      ImgReg1IN_290, D(1)=>ImgReg1IN_289, D(0)=>ImgReg1IN_288, CLK=>nx23938, 
      RST=>RST, EN=>nx23732, Q(15)=>OutputImg1_303_EXMPLR, Q(14)=>
      OutputImg1_302_EXMPLR, Q(13)=>OutputImg1_301_EXMPLR, Q(12)=>
      OutputImg1_300_EXMPLR, Q(11)=>OutputImg1_299_EXMPLR, Q(10)=>
      OutputImg1_298_EXMPLR, Q(9)=>OutputImg1_297_EXMPLR, Q(8)=>
      OutputImg1_296_EXMPLR, Q(7)=>OutputImg1_295_EXMPLR, Q(6)=>
      OutputImg1_294_EXMPLR, Q(5)=>OutputImg1_293_EXMPLR, Q(4)=>
      OutputImg1_292_EXMPLR, Q(3)=>OutputImg1_291_EXMPLR, Q(2)=>
      OutputImg1_290_EXMPLR, Q(1)=>OutputImg1_289_EXMPLR, Q(0)=>
      OutputImg1_288_EXMPLR);
   loop3_18_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_303, D(14)=>
      ImgReg2IN_302, D(13)=>ImgReg2IN_301, D(12)=>ImgReg2IN_300, D(11)=>
      ImgReg2IN_299, D(10)=>ImgReg2IN_298, D(9)=>ImgReg2IN_297, D(8)=>
      ImgReg2IN_296, D(7)=>ImgReg2IN_295, D(6)=>ImgReg2IN_294, D(5)=>
      ImgReg2IN_293, D(4)=>ImgReg2IN_292, D(3)=>ImgReg2IN_291, D(2)=>
      ImgReg2IN_290, D(1)=>ImgReg2IN_289, D(0)=>ImgReg2IN_288, CLK=>nx23938, 
      RST=>RST, EN=>nx23742, Q(15)=>OutputImg2_303_EXMPLR, Q(14)=>
      OutputImg2_302_EXMPLR, Q(13)=>OutputImg2_301_EXMPLR, Q(12)=>
      OutputImg2_300_EXMPLR, Q(11)=>OutputImg2_299_EXMPLR, Q(10)=>
      OutputImg2_298_EXMPLR, Q(9)=>OutputImg2_297_EXMPLR, Q(8)=>
      OutputImg2_296_EXMPLR, Q(7)=>OutputImg2_295_EXMPLR, Q(6)=>
      OutputImg2_294_EXMPLR, Q(5)=>OutputImg2_293_EXMPLR, Q(4)=>
      OutputImg2_292_EXMPLR, Q(3)=>OutputImg2_291_EXMPLR, Q(2)=>
      OutputImg2_290_EXMPLR, Q(1)=>OutputImg2_289_EXMPLR, Q(0)=>
      OutputImg2_288_EXMPLR);
   loop3_18_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_303, D(14)=>
      ImgReg3IN_302, D(13)=>ImgReg3IN_301, D(12)=>ImgReg3IN_300, D(11)=>
      ImgReg3IN_299, D(10)=>ImgReg3IN_298, D(9)=>ImgReg3IN_297, D(8)=>
      ImgReg3IN_296, D(7)=>ImgReg3IN_295, D(6)=>ImgReg3IN_294, D(5)=>
      ImgReg3IN_293, D(4)=>ImgReg3IN_292, D(3)=>ImgReg3IN_291, D(2)=>
      ImgReg3IN_290, D(1)=>ImgReg3IN_289, D(0)=>ImgReg3IN_288, CLK=>nx23940, 
      RST=>RST, EN=>nx23752, Q(15)=>OutputImg3_303_EXMPLR, Q(14)=>
      OutputImg3_302_EXMPLR, Q(13)=>OutputImg3_301_EXMPLR, Q(12)=>
      OutputImg3_300_EXMPLR, Q(11)=>OutputImg3_299_EXMPLR, Q(10)=>
      OutputImg3_298_EXMPLR, Q(9)=>OutputImg3_297_EXMPLR, Q(8)=>
      OutputImg3_296_EXMPLR, Q(7)=>OutputImg3_295_EXMPLR, Q(6)=>
      OutputImg3_294_EXMPLR, Q(5)=>OutputImg3_293_EXMPLR, Q(4)=>
      OutputImg3_292_EXMPLR, Q(3)=>OutputImg3_291_EXMPLR, Q(2)=>
      OutputImg3_290_EXMPLR, Q(1)=>OutputImg3_289_EXMPLR, Q(0)=>
      OutputImg3_288_EXMPLR);
   loop3_18_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_303, D(14)=>
      ImgReg4IN_302, D(13)=>ImgReg4IN_301, D(12)=>ImgReg4IN_300, D(11)=>
      ImgReg4IN_299, D(10)=>ImgReg4IN_298, D(9)=>ImgReg4IN_297, D(8)=>
      ImgReg4IN_296, D(7)=>ImgReg4IN_295, D(6)=>ImgReg4IN_294, D(5)=>
      ImgReg4IN_293, D(4)=>ImgReg4IN_292, D(3)=>ImgReg4IN_291, D(2)=>
      ImgReg4IN_290, D(1)=>ImgReg4IN_289, D(0)=>ImgReg4IN_288, CLK=>nx23940, 
      RST=>RST, EN=>nx23762, Q(15)=>OutputImg4_303_EXMPLR, Q(14)=>
      OutputImg4_302_EXMPLR, Q(13)=>OutputImg4_301_EXMPLR, Q(12)=>
      OutputImg4_300_EXMPLR, Q(11)=>OutputImg4_299_EXMPLR, Q(10)=>
      OutputImg4_298_EXMPLR, Q(9)=>OutputImg4_297_EXMPLR, Q(8)=>
      OutputImg4_296_EXMPLR, Q(7)=>OutputImg4_295_EXMPLR, Q(6)=>
      OutputImg4_294_EXMPLR, Q(5)=>OutputImg4_293_EXMPLR, Q(4)=>
      OutputImg4_292_EXMPLR, Q(3)=>OutputImg4_291_EXMPLR, Q(2)=>
      OutputImg4_290_EXMPLR, Q(1)=>OutputImg4_289_EXMPLR, Q(0)=>
      OutputImg4_288_EXMPLR);
   loop3_18_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_303, D(14)=>
      ImgReg5IN_302, D(13)=>ImgReg5IN_301, D(12)=>ImgReg5IN_300, D(11)=>
      ImgReg5IN_299, D(10)=>ImgReg5IN_298, D(9)=>ImgReg5IN_297, D(8)=>
      ImgReg5IN_296, D(7)=>ImgReg5IN_295, D(6)=>ImgReg5IN_294, D(5)=>
      ImgReg5IN_293, D(4)=>ImgReg5IN_292, D(3)=>ImgReg5IN_291, D(2)=>
      ImgReg5IN_290, D(1)=>ImgReg5IN_289, D(0)=>ImgReg5IN_288, CLK=>nx23942, 
      RST=>RST, EN=>nx23772, Q(15)=>OutputImg5_303_EXMPLR, Q(14)=>
      OutputImg5_302_EXMPLR, Q(13)=>OutputImg5_301_EXMPLR, Q(12)=>
      OutputImg5_300_EXMPLR, Q(11)=>OutputImg5_299_EXMPLR, Q(10)=>
      OutputImg5_298_EXMPLR, Q(9)=>OutputImg5_297_EXMPLR, Q(8)=>
      OutputImg5_296_EXMPLR, Q(7)=>OutputImg5_295_EXMPLR, Q(6)=>
      OutputImg5_294_EXMPLR, Q(5)=>OutputImg5_293_EXMPLR, Q(4)=>
      OutputImg5_292_EXMPLR, Q(3)=>OutputImg5_291_EXMPLR, Q(2)=>
      OutputImg5_290_EXMPLR, Q(1)=>OutputImg5_289_EXMPLR, Q(0)=>
      OutputImg5_288_EXMPLR);
   loop3_19_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_335_EXMPLR, D(14)=>OutputImg0_334_EXMPLR, D(13)=>
      OutputImg0_333_EXMPLR, D(12)=>OutputImg0_332_EXMPLR, D(11)=>
      OutputImg0_331_EXMPLR, D(10)=>OutputImg0_330_EXMPLR, D(9)=>
      OutputImg0_329_EXMPLR, D(8)=>OutputImg0_328_EXMPLR, D(7)=>
      OutputImg0_327_EXMPLR, D(6)=>OutputImg0_326_EXMPLR, D(5)=>
      OutputImg0_325_EXMPLR, D(4)=>OutputImg0_324_EXMPLR, D(3)=>
      OutputImg0_323_EXMPLR, D(2)=>OutputImg0_322_EXMPLR, D(1)=>
      OutputImg0_321_EXMPLR, D(0)=>OutputImg0_320_EXMPLR, EN=>nx23698, F(15)
      =>ImgReg0IN_319, F(14)=>ImgReg0IN_318, F(13)=>ImgReg0IN_317, F(12)=>
      ImgReg0IN_316, F(11)=>ImgReg0IN_315, F(10)=>ImgReg0IN_314, F(9)=>
      ImgReg0IN_313, F(8)=>ImgReg0IN_312, F(7)=>ImgReg0IN_311, F(6)=>
      ImgReg0IN_310, F(5)=>ImgReg0IN_309, F(4)=>ImgReg0IN_308, F(3)=>
      ImgReg0IN_307, F(2)=>ImgReg0IN_306, F(1)=>ImgReg0IN_305, F(0)=>
      ImgReg0IN_304);
   loop3_19_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_335_EXMPLR, D(14)=>OutputImg1_334_EXMPLR, D(13)=>
      OutputImg1_333_EXMPLR, D(12)=>OutputImg1_332_EXMPLR, D(11)=>
      OutputImg1_331_EXMPLR, D(10)=>OutputImg1_330_EXMPLR, D(9)=>
      OutputImg1_329_EXMPLR, D(8)=>OutputImg1_328_EXMPLR, D(7)=>
      OutputImg1_327_EXMPLR, D(6)=>OutputImg1_326_EXMPLR, D(5)=>
      OutputImg1_325_EXMPLR, D(4)=>OutputImg1_324_EXMPLR, D(3)=>
      OutputImg1_323_EXMPLR, D(2)=>OutputImg1_322_EXMPLR, D(1)=>
      OutputImg1_321_EXMPLR, D(0)=>OutputImg1_320_EXMPLR, EN=>nx23698, F(15)
      =>ImgReg1IN_319, F(14)=>ImgReg1IN_318, F(13)=>ImgReg1IN_317, F(12)=>
      ImgReg1IN_316, F(11)=>ImgReg1IN_315, F(10)=>ImgReg1IN_314, F(9)=>
      ImgReg1IN_313, F(8)=>ImgReg1IN_312, F(7)=>ImgReg1IN_311, F(6)=>
      ImgReg1IN_310, F(5)=>ImgReg1IN_309, F(4)=>ImgReg1IN_308, F(3)=>
      ImgReg1IN_307, F(2)=>ImgReg1IN_306, F(1)=>ImgReg1IN_305, F(0)=>
      ImgReg1IN_304);
   loop3_19_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_335_EXMPLR, D(14)=>OutputImg2_334_EXMPLR, D(13)=>
      OutputImg2_333_EXMPLR, D(12)=>OutputImg2_332_EXMPLR, D(11)=>
      OutputImg2_331_EXMPLR, D(10)=>OutputImg2_330_EXMPLR, D(9)=>
      OutputImg2_329_EXMPLR, D(8)=>OutputImg2_328_EXMPLR, D(7)=>
      OutputImg2_327_EXMPLR, D(6)=>OutputImg2_326_EXMPLR, D(5)=>
      OutputImg2_325_EXMPLR, D(4)=>OutputImg2_324_EXMPLR, D(3)=>
      OutputImg2_323_EXMPLR, D(2)=>OutputImg2_322_EXMPLR, D(1)=>
      OutputImg2_321_EXMPLR, D(0)=>OutputImg2_320_EXMPLR, EN=>nx23698, F(15)
      =>ImgReg2IN_319, F(14)=>ImgReg2IN_318, F(13)=>ImgReg2IN_317, F(12)=>
      ImgReg2IN_316, F(11)=>ImgReg2IN_315, F(10)=>ImgReg2IN_314, F(9)=>
      ImgReg2IN_313, F(8)=>ImgReg2IN_312, F(7)=>ImgReg2IN_311, F(6)=>
      ImgReg2IN_310, F(5)=>ImgReg2IN_309, F(4)=>ImgReg2IN_308, F(3)=>
      ImgReg2IN_307, F(2)=>ImgReg2IN_306, F(1)=>ImgReg2IN_305, F(0)=>
      ImgReg2IN_304);
   loop3_19_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_335_EXMPLR, D(14)=>OutputImg3_334_EXMPLR, D(13)=>
      OutputImg3_333_EXMPLR, D(12)=>OutputImg3_332_EXMPLR, D(11)=>
      OutputImg3_331_EXMPLR, D(10)=>OutputImg3_330_EXMPLR, D(9)=>
      OutputImg3_329_EXMPLR, D(8)=>OutputImg3_328_EXMPLR, D(7)=>
      OutputImg3_327_EXMPLR, D(6)=>OutputImg3_326_EXMPLR, D(5)=>
      OutputImg3_325_EXMPLR, D(4)=>OutputImg3_324_EXMPLR, D(3)=>
      OutputImg3_323_EXMPLR, D(2)=>OutputImg3_322_EXMPLR, D(1)=>
      OutputImg3_321_EXMPLR, D(0)=>OutputImg3_320_EXMPLR, EN=>nx23698, F(15)
      =>ImgReg3IN_319, F(14)=>ImgReg3IN_318, F(13)=>ImgReg3IN_317, F(12)=>
      ImgReg3IN_316, F(11)=>ImgReg3IN_315, F(10)=>ImgReg3IN_314, F(9)=>
      ImgReg3IN_313, F(8)=>ImgReg3IN_312, F(7)=>ImgReg3IN_311, F(6)=>
      ImgReg3IN_310, F(5)=>ImgReg3IN_309, F(4)=>ImgReg3IN_308, F(3)=>
      ImgReg3IN_307, F(2)=>ImgReg3IN_306, F(1)=>ImgReg3IN_305, F(0)=>
      ImgReg3IN_304);
   loop3_19_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_335_EXMPLR, D(14)=>OutputImg4_334_EXMPLR, D(13)=>
      OutputImg4_333_EXMPLR, D(12)=>OutputImg4_332_EXMPLR, D(11)=>
      OutputImg4_331_EXMPLR, D(10)=>OutputImg4_330_EXMPLR, D(9)=>
      OutputImg4_329_EXMPLR, D(8)=>OutputImg4_328_EXMPLR, D(7)=>
      OutputImg4_327_EXMPLR, D(6)=>OutputImg4_326_EXMPLR, D(5)=>
      OutputImg4_325_EXMPLR, D(4)=>OutputImg4_324_EXMPLR, D(3)=>
      OutputImg4_323_EXMPLR, D(2)=>OutputImg4_322_EXMPLR, D(1)=>
      OutputImg4_321_EXMPLR, D(0)=>OutputImg4_320_EXMPLR, EN=>nx23698, F(15)
      =>ImgReg4IN_319, F(14)=>ImgReg4IN_318, F(13)=>ImgReg4IN_317, F(12)=>
      ImgReg4IN_316, F(11)=>ImgReg4IN_315, F(10)=>ImgReg4IN_314, F(9)=>
      ImgReg4IN_313, F(8)=>ImgReg4IN_312, F(7)=>ImgReg4IN_311, F(6)=>
      ImgReg4IN_310, F(5)=>ImgReg4IN_309, F(4)=>ImgReg4IN_308, F(3)=>
      ImgReg4IN_307, F(2)=>ImgReg4IN_306, F(1)=>ImgReg4IN_305, F(0)=>
      ImgReg4IN_304);
   loop3_19_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_335_EXMPLR, D(14)=>OutputImg5_334_EXMPLR, D(13)=>
      OutputImg5_333_EXMPLR, D(12)=>OutputImg5_332_EXMPLR, D(11)=>
      OutputImg5_331_EXMPLR, D(10)=>OutputImg5_330_EXMPLR, D(9)=>
      OutputImg5_329_EXMPLR, D(8)=>OutputImg5_328_EXMPLR, D(7)=>
      OutputImg5_327_EXMPLR, D(6)=>OutputImg5_326_EXMPLR, D(5)=>
      OutputImg5_325_EXMPLR, D(4)=>OutputImg5_324_EXMPLR, D(3)=>
      OutputImg5_323_EXMPLR, D(2)=>OutputImg5_322_EXMPLR, D(1)=>
      OutputImg5_321_EXMPLR, D(0)=>OutputImg5_320_EXMPLR, EN=>nx23700, F(15)
      =>ImgReg5IN_319, F(14)=>ImgReg5IN_318, F(13)=>ImgReg5IN_317, F(12)=>
      ImgReg5IN_316, F(11)=>ImgReg5IN_315, F(10)=>ImgReg5IN_314, F(9)=>
      ImgReg5IN_313, F(8)=>ImgReg5IN_312, F(7)=>ImgReg5IN_311, F(6)=>
      ImgReg5IN_310, F(5)=>ImgReg5IN_309, F(4)=>ImgReg5IN_308, F(3)=>
      ImgReg5IN_307, F(2)=>ImgReg5IN_306, F(1)=>ImgReg5IN_305, F(0)=>
      ImgReg5IN_304);
   loop3_19_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(319), 
      D(14)=>DATA(318), D(13)=>DATA(317), D(12)=>DATA(316), D(11)=>DATA(315), 
      D(10)=>DATA(314), D(9)=>DATA(313), D(8)=>DATA(312), D(7)=>DATA(311), 
      D(6)=>DATA(310), D(5)=>DATA(309), D(4)=>DATA(308), D(3)=>DATA(307), 
      D(2)=>DATA(306), D(1)=>DATA(305), D(0)=>DATA(304), EN=>nx23658, F(15)
      =>ImgReg0IN_319, F(14)=>ImgReg0IN_318, F(13)=>ImgReg0IN_317, F(12)=>
      ImgReg0IN_316, F(11)=>ImgReg0IN_315, F(10)=>ImgReg0IN_314, F(9)=>
      ImgReg0IN_313, F(8)=>ImgReg0IN_312, F(7)=>ImgReg0IN_311, F(6)=>
      ImgReg0IN_310, F(5)=>ImgReg0IN_309, F(4)=>ImgReg0IN_308, F(3)=>
      ImgReg0IN_307, F(2)=>ImgReg0IN_306, F(1)=>ImgReg0IN_305, F(0)=>
      ImgReg0IN_304);
   loop3_19_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(319), 
      D(14)=>DATA(318), D(13)=>DATA(317), D(12)=>DATA(316), D(11)=>DATA(315), 
      D(10)=>DATA(314), D(9)=>DATA(313), D(8)=>DATA(312), D(7)=>DATA(311), 
      D(6)=>DATA(310), D(5)=>DATA(309), D(4)=>DATA(308), D(3)=>DATA(307), 
      D(2)=>DATA(306), D(1)=>DATA(305), D(0)=>DATA(304), EN=>nx23646, F(15)
      =>ImgReg1IN_319, F(14)=>ImgReg1IN_318, F(13)=>ImgReg1IN_317, F(12)=>
      ImgReg1IN_316, F(11)=>ImgReg1IN_315, F(10)=>ImgReg1IN_314, F(9)=>
      ImgReg1IN_313, F(8)=>ImgReg1IN_312, F(7)=>ImgReg1IN_311, F(6)=>
      ImgReg1IN_310, F(5)=>ImgReg1IN_309, F(4)=>ImgReg1IN_308, F(3)=>
      ImgReg1IN_307, F(2)=>ImgReg1IN_306, F(1)=>ImgReg1IN_305, F(0)=>
      ImgReg1IN_304);
   loop3_19_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(319), 
      D(14)=>DATA(318), D(13)=>DATA(317), D(12)=>DATA(316), D(11)=>DATA(315), 
      D(10)=>DATA(314), D(9)=>DATA(313), D(8)=>DATA(312), D(7)=>DATA(311), 
      D(6)=>DATA(310), D(5)=>DATA(309), D(4)=>DATA(308), D(3)=>DATA(307), 
      D(2)=>DATA(306), D(1)=>DATA(305), D(0)=>DATA(304), EN=>nx23634, F(15)
      =>ImgReg2IN_319, F(14)=>ImgReg2IN_318, F(13)=>ImgReg2IN_317, F(12)=>
      ImgReg2IN_316, F(11)=>ImgReg2IN_315, F(10)=>ImgReg2IN_314, F(9)=>
      ImgReg2IN_313, F(8)=>ImgReg2IN_312, F(7)=>ImgReg2IN_311, F(6)=>
      ImgReg2IN_310, F(5)=>ImgReg2IN_309, F(4)=>ImgReg2IN_308, F(3)=>
      ImgReg2IN_307, F(2)=>ImgReg2IN_306, F(1)=>ImgReg2IN_305, F(0)=>
      ImgReg2IN_304);
   loop3_19_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(319), 
      D(14)=>DATA(318), D(13)=>DATA(317), D(12)=>DATA(316), D(11)=>DATA(315), 
      D(10)=>DATA(314), D(9)=>DATA(313), D(8)=>DATA(312), D(7)=>DATA(311), 
      D(6)=>DATA(310), D(5)=>DATA(309), D(4)=>DATA(308), D(3)=>DATA(307), 
      D(2)=>DATA(306), D(1)=>DATA(305), D(0)=>DATA(304), EN=>nx23622, F(15)
      =>ImgReg3IN_319, F(14)=>ImgReg3IN_318, F(13)=>ImgReg3IN_317, F(12)=>
      ImgReg3IN_316, F(11)=>ImgReg3IN_315, F(10)=>ImgReg3IN_314, F(9)=>
      ImgReg3IN_313, F(8)=>ImgReg3IN_312, F(7)=>ImgReg3IN_311, F(6)=>
      ImgReg3IN_310, F(5)=>ImgReg3IN_309, F(4)=>ImgReg3IN_308, F(3)=>
      ImgReg3IN_307, F(2)=>ImgReg3IN_306, F(1)=>ImgReg3IN_305, F(0)=>
      ImgReg3IN_304);
   loop3_19_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(319), 
      D(14)=>DATA(318), D(13)=>DATA(317), D(12)=>DATA(316), D(11)=>DATA(315), 
      D(10)=>DATA(314), D(9)=>DATA(313), D(8)=>DATA(312), D(7)=>DATA(311), 
      D(6)=>DATA(310), D(5)=>DATA(309), D(4)=>DATA(308), D(3)=>DATA(307), 
      D(2)=>DATA(306), D(1)=>DATA(305), D(0)=>DATA(304), EN=>nx23610, F(15)
      =>ImgReg4IN_319, F(14)=>ImgReg4IN_318, F(13)=>ImgReg4IN_317, F(12)=>
      ImgReg4IN_316, F(11)=>ImgReg4IN_315, F(10)=>ImgReg4IN_314, F(9)=>
      ImgReg4IN_313, F(8)=>ImgReg4IN_312, F(7)=>ImgReg4IN_311, F(6)=>
      ImgReg4IN_310, F(5)=>ImgReg4IN_309, F(4)=>ImgReg4IN_308, F(3)=>
      ImgReg4IN_307, F(2)=>ImgReg4IN_306, F(1)=>ImgReg4IN_305, F(0)=>
      ImgReg4IN_304);
   loop3_19_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(319), 
      D(14)=>DATA(318), D(13)=>DATA(317), D(12)=>DATA(316), D(11)=>DATA(315), 
      D(10)=>DATA(314), D(9)=>DATA(313), D(8)=>DATA(312), D(7)=>DATA(311), 
      D(6)=>DATA(310), D(5)=>DATA(309), D(4)=>DATA(308), D(3)=>DATA(307), 
      D(2)=>DATA(306), D(1)=>DATA(305), D(0)=>DATA(304), EN=>nx23598, F(15)
      =>ImgReg5IN_319, F(14)=>ImgReg5IN_318, F(13)=>ImgReg5IN_317, F(12)=>
      ImgReg5IN_316, F(11)=>ImgReg5IN_315, F(10)=>ImgReg5IN_314, F(9)=>
      ImgReg5IN_313, F(8)=>ImgReg5IN_312, F(7)=>ImgReg5IN_311, F(6)=>
      ImgReg5IN_310, F(5)=>ImgReg5IN_309, F(4)=>ImgReg5IN_308, F(3)=>
      ImgReg5IN_307, F(2)=>ImgReg5IN_306, F(1)=>ImgReg5IN_305, F(0)=>
      ImgReg5IN_304);
   loop3_19_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_319_EXMPLR, D(14)=>OutputImg1_318_EXMPLR, D(13)=>
      OutputImg1_317_EXMPLR, D(12)=>OutputImg1_316_EXMPLR, D(11)=>
      OutputImg1_315_EXMPLR, D(10)=>OutputImg1_314_EXMPLR, D(9)=>
      OutputImg1_313_EXMPLR, D(8)=>OutputImg1_312_EXMPLR, D(7)=>
      OutputImg1_311_EXMPLR, D(6)=>OutputImg1_310_EXMPLR, D(5)=>
      OutputImg1_309_EXMPLR, D(4)=>OutputImg1_308_EXMPLR, D(3)=>
      OutputImg1_307_EXMPLR, D(2)=>OutputImg1_306_EXMPLR, D(1)=>
      OutputImg1_305_EXMPLR, D(0)=>OutputImg1_304_EXMPLR, EN=>nx23812, F(15)
      =>ImgReg0IN_319, F(14)=>ImgReg0IN_318, F(13)=>ImgReg0IN_317, F(12)=>
      ImgReg0IN_316, F(11)=>ImgReg0IN_315, F(10)=>ImgReg0IN_314, F(9)=>
      ImgReg0IN_313, F(8)=>ImgReg0IN_312, F(7)=>ImgReg0IN_311, F(6)=>
      ImgReg0IN_310, F(5)=>ImgReg0IN_309, F(4)=>ImgReg0IN_308, F(3)=>
      ImgReg0IN_307, F(2)=>ImgReg0IN_306, F(1)=>ImgReg0IN_305, F(0)=>
      ImgReg0IN_304);
   loop3_19_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_319_EXMPLR, D(14)=>OutputImg2_318_EXMPLR, D(13)=>
      OutputImg2_317_EXMPLR, D(12)=>OutputImg2_316_EXMPLR, D(11)=>
      OutputImg2_315_EXMPLR, D(10)=>OutputImg2_314_EXMPLR, D(9)=>
      OutputImg2_313_EXMPLR, D(8)=>OutputImg2_312_EXMPLR, D(7)=>
      OutputImg2_311_EXMPLR, D(6)=>OutputImg2_310_EXMPLR, D(5)=>
      OutputImg2_309_EXMPLR, D(4)=>OutputImg2_308_EXMPLR, D(3)=>
      OutputImg2_307_EXMPLR, D(2)=>OutputImg2_306_EXMPLR, D(1)=>
      OutputImg2_305_EXMPLR, D(0)=>OutputImg2_304_EXMPLR, EN=>nx23812, F(15)
      =>ImgReg1IN_319, F(14)=>ImgReg1IN_318, F(13)=>ImgReg1IN_317, F(12)=>
      ImgReg1IN_316, F(11)=>ImgReg1IN_315, F(10)=>ImgReg1IN_314, F(9)=>
      ImgReg1IN_313, F(8)=>ImgReg1IN_312, F(7)=>ImgReg1IN_311, F(6)=>
      ImgReg1IN_310, F(5)=>ImgReg1IN_309, F(4)=>ImgReg1IN_308, F(3)=>
      ImgReg1IN_307, F(2)=>ImgReg1IN_306, F(1)=>ImgReg1IN_305, F(0)=>
      ImgReg1IN_304);
   loop3_19_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_319_EXMPLR, D(14)=>OutputImg3_318_EXMPLR, D(13)=>
      OutputImg3_317_EXMPLR, D(12)=>OutputImg3_316_EXMPLR, D(11)=>
      OutputImg3_315_EXMPLR, D(10)=>OutputImg3_314_EXMPLR, D(9)=>
      OutputImg3_313_EXMPLR, D(8)=>OutputImg3_312_EXMPLR, D(7)=>
      OutputImg3_311_EXMPLR, D(6)=>OutputImg3_310_EXMPLR, D(5)=>
      OutputImg3_309_EXMPLR, D(4)=>OutputImg3_308_EXMPLR, D(3)=>
      OutputImg3_307_EXMPLR, D(2)=>OutputImg3_306_EXMPLR, D(1)=>
      OutputImg3_305_EXMPLR, D(0)=>OutputImg3_304_EXMPLR, EN=>nx23812, F(15)
      =>ImgReg2IN_319, F(14)=>ImgReg2IN_318, F(13)=>ImgReg2IN_317, F(12)=>
      ImgReg2IN_316, F(11)=>ImgReg2IN_315, F(10)=>ImgReg2IN_314, F(9)=>
      ImgReg2IN_313, F(8)=>ImgReg2IN_312, F(7)=>ImgReg2IN_311, F(6)=>
      ImgReg2IN_310, F(5)=>ImgReg2IN_309, F(4)=>ImgReg2IN_308, F(3)=>
      ImgReg2IN_307, F(2)=>ImgReg2IN_306, F(1)=>ImgReg2IN_305, F(0)=>
      ImgReg2IN_304);
   loop3_19_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_319_EXMPLR, D(14)=>OutputImg4_318_EXMPLR, D(13)=>
      OutputImg4_317_EXMPLR, D(12)=>OutputImg4_316_EXMPLR, D(11)=>
      OutputImg4_315_EXMPLR, D(10)=>OutputImg4_314_EXMPLR, D(9)=>
      OutputImg4_313_EXMPLR, D(8)=>OutputImg4_312_EXMPLR, D(7)=>
      OutputImg4_311_EXMPLR, D(6)=>OutputImg4_310_EXMPLR, D(5)=>
      OutputImg4_309_EXMPLR, D(4)=>OutputImg4_308_EXMPLR, D(3)=>
      OutputImg4_307_EXMPLR, D(2)=>OutputImg4_306_EXMPLR, D(1)=>
      OutputImg4_305_EXMPLR, D(0)=>OutputImg4_304_EXMPLR, EN=>nx23814, F(15)
      =>ImgReg3IN_319, F(14)=>ImgReg3IN_318, F(13)=>ImgReg3IN_317, F(12)=>
      ImgReg3IN_316, F(11)=>ImgReg3IN_315, F(10)=>ImgReg3IN_314, F(9)=>
      ImgReg3IN_313, F(8)=>ImgReg3IN_312, F(7)=>ImgReg3IN_311, F(6)=>
      ImgReg3IN_310, F(5)=>ImgReg3IN_309, F(4)=>ImgReg3IN_308, F(3)=>
      ImgReg3IN_307, F(2)=>ImgReg3IN_306, F(1)=>ImgReg3IN_305, F(0)=>
      ImgReg3IN_304);
   loop3_19_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_319_EXMPLR, D(14)=>OutputImg5_318_EXMPLR, D(13)=>
      OutputImg5_317_EXMPLR, D(12)=>OutputImg5_316_EXMPLR, D(11)=>
      OutputImg5_315_EXMPLR, D(10)=>OutputImg5_314_EXMPLR, D(9)=>
      OutputImg5_313_EXMPLR, D(8)=>OutputImg5_312_EXMPLR, D(7)=>
      OutputImg5_311_EXMPLR, D(6)=>OutputImg5_310_EXMPLR, D(5)=>
      OutputImg5_309_EXMPLR, D(4)=>OutputImg5_308_EXMPLR, D(3)=>
      OutputImg5_307_EXMPLR, D(2)=>OutputImg5_306_EXMPLR, D(1)=>
      OutputImg5_305_EXMPLR, D(0)=>OutputImg5_304_EXMPLR, EN=>nx23814, F(15)
      =>ImgReg4IN_319, F(14)=>ImgReg4IN_318, F(13)=>ImgReg4IN_317, F(12)=>
      ImgReg4IN_316, F(11)=>ImgReg4IN_315, F(10)=>ImgReg4IN_314, F(9)=>
      ImgReg4IN_313, F(8)=>ImgReg4IN_312, F(7)=>ImgReg4IN_311, F(6)=>
      ImgReg4IN_310, F(5)=>ImgReg4IN_309, F(4)=>ImgReg4IN_308, F(3)=>
      ImgReg4IN_307, F(2)=>ImgReg4IN_306, F(1)=>ImgReg4IN_305, F(0)=>
      ImgReg4IN_304);
   loop3_19_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_319, D(14)=>
      ImgReg0IN_318, D(13)=>ImgReg0IN_317, D(12)=>ImgReg0IN_316, D(11)=>
      ImgReg0IN_315, D(10)=>ImgReg0IN_314, D(9)=>ImgReg0IN_313, D(8)=>
      ImgReg0IN_312, D(7)=>ImgReg0IN_311, D(6)=>ImgReg0IN_310, D(5)=>
      ImgReg0IN_309, D(4)=>ImgReg0IN_308, D(3)=>ImgReg0IN_307, D(2)=>
      ImgReg0IN_306, D(1)=>ImgReg0IN_305, D(0)=>ImgReg0IN_304, CLK=>nx23942, 
      RST=>RST, EN=>nx23722, Q(15)=>OutputImg0_319_EXMPLR, Q(14)=>
      OutputImg0_318_EXMPLR, Q(13)=>OutputImg0_317_EXMPLR, Q(12)=>
      OutputImg0_316_EXMPLR, Q(11)=>OutputImg0_315_EXMPLR, Q(10)=>
      OutputImg0_314_EXMPLR, Q(9)=>OutputImg0_313_EXMPLR, Q(8)=>
      OutputImg0_312_EXMPLR, Q(7)=>OutputImg0_311_EXMPLR, Q(6)=>
      OutputImg0_310_EXMPLR, Q(5)=>OutputImg0_309_EXMPLR, Q(4)=>
      OutputImg0_308_EXMPLR, Q(3)=>OutputImg0_307_EXMPLR, Q(2)=>
      OutputImg0_306_EXMPLR, Q(1)=>OutputImg0_305_EXMPLR, Q(0)=>
      OutputImg0_304_EXMPLR);
   loop3_19_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_319, D(14)=>
      ImgReg1IN_318, D(13)=>ImgReg1IN_317, D(12)=>ImgReg1IN_316, D(11)=>
      ImgReg1IN_315, D(10)=>ImgReg1IN_314, D(9)=>ImgReg1IN_313, D(8)=>
      ImgReg1IN_312, D(7)=>ImgReg1IN_311, D(6)=>ImgReg1IN_310, D(5)=>
      ImgReg1IN_309, D(4)=>ImgReg1IN_308, D(3)=>ImgReg1IN_307, D(2)=>
      ImgReg1IN_306, D(1)=>ImgReg1IN_305, D(0)=>ImgReg1IN_304, CLK=>nx23944, 
      RST=>RST, EN=>nx23732, Q(15)=>OutputImg1_319_EXMPLR, Q(14)=>
      OutputImg1_318_EXMPLR, Q(13)=>OutputImg1_317_EXMPLR, Q(12)=>
      OutputImg1_316_EXMPLR, Q(11)=>OutputImg1_315_EXMPLR, Q(10)=>
      OutputImg1_314_EXMPLR, Q(9)=>OutputImg1_313_EXMPLR, Q(8)=>
      OutputImg1_312_EXMPLR, Q(7)=>OutputImg1_311_EXMPLR, Q(6)=>
      OutputImg1_310_EXMPLR, Q(5)=>OutputImg1_309_EXMPLR, Q(4)=>
      OutputImg1_308_EXMPLR, Q(3)=>OutputImg1_307_EXMPLR, Q(2)=>
      OutputImg1_306_EXMPLR, Q(1)=>OutputImg1_305_EXMPLR, Q(0)=>
      OutputImg1_304_EXMPLR);
   loop3_19_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_319, D(14)=>
      ImgReg2IN_318, D(13)=>ImgReg2IN_317, D(12)=>ImgReg2IN_316, D(11)=>
      ImgReg2IN_315, D(10)=>ImgReg2IN_314, D(9)=>ImgReg2IN_313, D(8)=>
      ImgReg2IN_312, D(7)=>ImgReg2IN_311, D(6)=>ImgReg2IN_310, D(5)=>
      ImgReg2IN_309, D(4)=>ImgReg2IN_308, D(3)=>ImgReg2IN_307, D(2)=>
      ImgReg2IN_306, D(1)=>ImgReg2IN_305, D(0)=>ImgReg2IN_304, CLK=>nx23944, 
      RST=>RST, EN=>nx23742, Q(15)=>OutputImg2_319_EXMPLR, Q(14)=>
      OutputImg2_318_EXMPLR, Q(13)=>OutputImg2_317_EXMPLR, Q(12)=>
      OutputImg2_316_EXMPLR, Q(11)=>OutputImg2_315_EXMPLR, Q(10)=>
      OutputImg2_314_EXMPLR, Q(9)=>OutputImg2_313_EXMPLR, Q(8)=>
      OutputImg2_312_EXMPLR, Q(7)=>OutputImg2_311_EXMPLR, Q(6)=>
      OutputImg2_310_EXMPLR, Q(5)=>OutputImg2_309_EXMPLR, Q(4)=>
      OutputImg2_308_EXMPLR, Q(3)=>OutputImg2_307_EXMPLR, Q(2)=>
      OutputImg2_306_EXMPLR, Q(1)=>OutputImg2_305_EXMPLR, Q(0)=>
      OutputImg2_304_EXMPLR);
   loop3_19_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_319, D(14)=>
      ImgReg3IN_318, D(13)=>ImgReg3IN_317, D(12)=>ImgReg3IN_316, D(11)=>
      ImgReg3IN_315, D(10)=>ImgReg3IN_314, D(9)=>ImgReg3IN_313, D(8)=>
      ImgReg3IN_312, D(7)=>ImgReg3IN_311, D(6)=>ImgReg3IN_310, D(5)=>
      ImgReg3IN_309, D(4)=>ImgReg3IN_308, D(3)=>ImgReg3IN_307, D(2)=>
      ImgReg3IN_306, D(1)=>ImgReg3IN_305, D(0)=>ImgReg3IN_304, CLK=>nx23946, 
      RST=>RST, EN=>nx23752, Q(15)=>OutputImg3_319_EXMPLR, Q(14)=>
      OutputImg3_318_EXMPLR, Q(13)=>OutputImg3_317_EXMPLR, Q(12)=>
      OutputImg3_316_EXMPLR, Q(11)=>OutputImg3_315_EXMPLR, Q(10)=>
      OutputImg3_314_EXMPLR, Q(9)=>OutputImg3_313_EXMPLR, Q(8)=>
      OutputImg3_312_EXMPLR, Q(7)=>OutputImg3_311_EXMPLR, Q(6)=>
      OutputImg3_310_EXMPLR, Q(5)=>OutputImg3_309_EXMPLR, Q(4)=>
      OutputImg3_308_EXMPLR, Q(3)=>OutputImg3_307_EXMPLR, Q(2)=>
      OutputImg3_306_EXMPLR, Q(1)=>OutputImg3_305_EXMPLR, Q(0)=>
      OutputImg3_304_EXMPLR);
   loop3_19_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_319, D(14)=>
      ImgReg4IN_318, D(13)=>ImgReg4IN_317, D(12)=>ImgReg4IN_316, D(11)=>
      ImgReg4IN_315, D(10)=>ImgReg4IN_314, D(9)=>ImgReg4IN_313, D(8)=>
      ImgReg4IN_312, D(7)=>ImgReg4IN_311, D(6)=>ImgReg4IN_310, D(5)=>
      ImgReg4IN_309, D(4)=>ImgReg4IN_308, D(3)=>ImgReg4IN_307, D(2)=>
      ImgReg4IN_306, D(1)=>ImgReg4IN_305, D(0)=>ImgReg4IN_304, CLK=>nx23946, 
      RST=>RST, EN=>nx23762, Q(15)=>OutputImg4_319_EXMPLR, Q(14)=>
      OutputImg4_318_EXMPLR, Q(13)=>OutputImg4_317_EXMPLR, Q(12)=>
      OutputImg4_316_EXMPLR, Q(11)=>OutputImg4_315_EXMPLR, Q(10)=>
      OutputImg4_314_EXMPLR, Q(9)=>OutputImg4_313_EXMPLR, Q(8)=>
      OutputImg4_312_EXMPLR, Q(7)=>OutputImg4_311_EXMPLR, Q(6)=>
      OutputImg4_310_EXMPLR, Q(5)=>OutputImg4_309_EXMPLR, Q(4)=>
      OutputImg4_308_EXMPLR, Q(3)=>OutputImg4_307_EXMPLR, Q(2)=>
      OutputImg4_306_EXMPLR, Q(1)=>OutputImg4_305_EXMPLR, Q(0)=>
      OutputImg4_304_EXMPLR);
   loop3_19_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_319, D(14)=>
      ImgReg5IN_318, D(13)=>ImgReg5IN_317, D(12)=>ImgReg5IN_316, D(11)=>
      ImgReg5IN_315, D(10)=>ImgReg5IN_314, D(9)=>ImgReg5IN_313, D(8)=>
      ImgReg5IN_312, D(7)=>ImgReg5IN_311, D(6)=>ImgReg5IN_310, D(5)=>
      ImgReg5IN_309, D(4)=>ImgReg5IN_308, D(3)=>ImgReg5IN_307, D(2)=>
      ImgReg5IN_306, D(1)=>ImgReg5IN_305, D(0)=>ImgReg5IN_304, CLK=>nx23948, 
      RST=>RST, EN=>nx23772, Q(15)=>OutputImg5_319_EXMPLR, Q(14)=>
      OutputImg5_318_EXMPLR, Q(13)=>OutputImg5_317_EXMPLR, Q(12)=>
      OutputImg5_316_EXMPLR, Q(11)=>OutputImg5_315_EXMPLR, Q(10)=>
      OutputImg5_314_EXMPLR, Q(9)=>OutputImg5_313_EXMPLR, Q(8)=>
      OutputImg5_312_EXMPLR, Q(7)=>OutputImg5_311_EXMPLR, Q(6)=>
      OutputImg5_310_EXMPLR, Q(5)=>OutputImg5_309_EXMPLR, Q(4)=>
      OutputImg5_308_EXMPLR, Q(3)=>OutputImg5_307_EXMPLR, Q(2)=>
      OutputImg5_306_EXMPLR, Q(1)=>OutputImg5_305_EXMPLR, Q(0)=>
      OutputImg5_304_EXMPLR);
   loop3_20_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_351_EXMPLR, D(14)=>OutputImg0_350_EXMPLR, D(13)=>
      OutputImg0_349_EXMPLR, D(12)=>OutputImg0_348_EXMPLR, D(11)=>
      OutputImg0_347_EXMPLR, D(10)=>OutputImg0_346_EXMPLR, D(9)=>
      OutputImg0_345_EXMPLR, D(8)=>OutputImg0_344_EXMPLR, D(7)=>
      OutputImg0_343_EXMPLR, D(6)=>OutputImg0_342_EXMPLR, D(5)=>
      OutputImg0_341_EXMPLR, D(4)=>OutputImg0_340_EXMPLR, D(3)=>
      OutputImg0_339_EXMPLR, D(2)=>OutputImg0_338_EXMPLR, D(1)=>
      OutputImg0_337_EXMPLR, D(0)=>OutputImg0_336_EXMPLR, EN=>nx23700, F(15)
      =>ImgReg0IN_335, F(14)=>ImgReg0IN_334, F(13)=>ImgReg0IN_333, F(12)=>
      ImgReg0IN_332, F(11)=>ImgReg0IN_331, F(10)=>ImgReg0IN_330, F(9)=>
      ImgReg0IN_329, F(8)=>ImgReg0IN_328, F(7)=>ImgReg0IN_327, F(6)=>
      ImgReg0IN_326, F(5)=>ImgReg0IN_325, F(4)=>ImgReg0IN_324, F(3)=>
      ImgReg0IN_323, F(2)=>ImgReg0IN_322, F(1)=>ImgReg0IN_321, F(0)=>
      ImgReg0IN_320);
   loop3_20_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_351_EXMPLR, D(14)=>OutputImg1_350_EXMPLR, D(13)=>
      OutputImg1_349_EXMPLR, D(12)=>OutputImg1_348_EXMPLR, D(11)=>
      OutputImg1_347_EXMPLR, D(10)=>OutputImg1_346_EXMPLR, D(9)=>
      OutputImg1_345_EXMPLR, D(8)=>OutputImg1_344_EXMPLR, D(7)=>
      OutputImg1_343_EXMPLR, D(6)=>OutputImg1_342_EXMPLR, D(5)=>
      OutputImg1_341_EXMPLR, D(4)=>OutputImg1_340_EXMPLR, D(3)=>
      OutputImg1_339_EXMPLR, D(2)=>OutputImg1_338_EXMPLR, D(1)=>
      OutputImg1_337_EXMPLR, D(0)=>OutputImg1_336_EXMPLR, EN=>nx23700, F(15)
      =>ImgReg1IN_335, F(14)=>ImgReg1IN_334, F(13)=>ImgReg1IN_333, F(12)=>
      ImgReg1IN_332, F(11)=>ImgReg1IN_331, F(10)=>ImgReg1IN_330, F(9)=>
      ImgReg1IN_329, F(8)=>ImgReg1IN_328, F(7)=>ImgReg1IN_327, F(6)=>
      ImgReg1IN_326, F(5)=>ImgReg1IN_325, F(4)=>ImgReg1IN_324, F(3)=>
      ImgReg1IN_323, F(2)=>ImgReg1IN_322, F(1)=>ImgReg1IN_321, F(0)=>
      ImgReg1IN_320);
   loop3_20_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_351_EXMPLR, D(14)=>OutputImg2_350_EXMPLR, D(13)=>
      OutputImg2_349_EXMPLR, D(12)=>OutputImg2_348_EXMPLR, D(11)=>
      OutputImg2_347_EXMPLR, D(10)=>OutputImg2_346_EXMPLR, D(9)=>
      OutputImg2_345_EXMPLR, D(8)=>OutputImg2_344_EXMPLR, D(7)=>
      OutputImg2_343_EXMPLR, D(6)=>OutputImg2_342_EXMPLR, D(5)=>
      OutputImg2_341_EXMPLR, D(4)=>OutputImg2_340_EXMPLR, D(3)=>
      OutputImg2_339_EXMPLR, D(2)=>OutputImg2_338_EXMPLR, D(1)=>
      OutputImg2_337_EXMPLR, D(0)=>OutputImg2_336_EXMPLR, EN=>nx23700, F(15)
      =>ImgReg2IN_335, F(14)=>ImgReg2IN_334, F(13)=>ImgReg2IN_333, F(12)=>
      ImgReg2IN_332, F(11)=>ImgReg2IN_331, F(10)=>ImgReg2IN_330, F(9)=>
      ImgReg2IN_329, F(8)=>ImgReg2IN_328, F(7)=>ImgReg2IN_327, F(6)=>
      ImgReg2IN_326, F(5)=>ImgReg2IN_325, F(4)=>ImgReg2IN_324, F(3)=>
      ImgReg2IN_323, F(2)=>ImgReg2IN_322, F(1)=>ImgReg2IN_321, F(0)=>
      ImgReg2IN_320);
   loop3_20_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_351_EXMPLR, D(14)=>OutputImg3_350_EXMPLR, D(13)=>
      OutputImg3_349_EXMPLR, D(12)=>OutputImg3_348_EXMPLR, D(11)=>
      OutputImg3_347_EXMPLR, D(10)=>OutputImg3_346_EXMPLR, D(9)=>
      OutputImg3_345_EXMPLR, D(8)=>OutputImg3_344_EXMPLR, D(7)=>
      OutputImg3_343_EXMPLR, D(6)=>OutputImg3_342_EXMPLR, D(5)=>
      OutputImg3_341_EXMPLR, D(4)=>OutputImg3_340_EXMPLR, D(3)=>
      OutputImg3_339_EXMPLR, D(2)=>OutputImg3_338_EXMPLR, D(1)=>
      OutputImg3_337_EXMPLR, D(0)=>OutputImg3_336_EXMPLR, EN=>nx23700, F(15)
      =>ImgReg3IN_335, F(14)=>ImgReg3IN_334, F(13)=>ImgReg3IN_333, F(12)=>
      ImgReg3IN_332, F(11)=>ImgReg3IN_331, F(10)=>ImgReg3IN_330, F(9)=>
      ImgReg3IN_329, F(8)=>ImgReg3IN_328, F(7)=>ImgReg3IN_327, F(6)=>
      ImgReg3IN_326, F(5)=>ImgReg3IN_325, F(4)=>ImgReg3IN_324, F(3)=>
      ImgReg3IN_323, F(2)=>ImgReg3IN_322, F(1)=>ImgReg3IN_321, F(0)=>
      ImgReg3IN_320);
   loop3_20_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_351_EXMPLR, D(14)=>OutputImg4_350_EXMPLR, D(13)=>
      OutputImg4_349_EXMPLR, D(12)=>OutputImg4_348_EXMPLR, D(11)=>
      OutputImg4_347_EXMPLR, D(10)=>OutputImg4_346_EXMPLR, D(9)=>
      OutputImg4_345_EXMPLR, D(8)=>OutputImg4_344_EXMPLR, D(7)=>
      OutputImg4_343_EXMPLR, D(6)=>OutputImg4_342_EXMPLR, D(5)=>
      OutputImg4_341_EXMPLR, D(4)=>OutputImg4_340_EXMPLR, D(3)=>
      OutputImg4_339_EXMPLR, D(2)=>OutputImg4_338_EXMPLR, D(1)=>
      OutputImg4_337_EXMPLR, D(0)=>OutputImg4_336_EXMPLR, EN=>nx23700, F(15)
      =>ImgReg4IN_335, F(14)=>ImgReg4IN_334, F(13)=>ImgReg4IN_333, F(12)=>
      ImgReg4IN_332, F(11)=>ImgReg4IN_331, F(10)=>ImgReg4IN_330, F(9)=>
      ImgReg4IN_329, F(8)=>ImgReg4IN_328, F(7)=>ImgReg4IN_327, F(6)=>
      ImgReg4IN_326, F(5)=>ImgReg4IN_325, F(4)=>ImgReg4IN_324, F(3)=>
      ImgReg4IN_323, F(2)=>ImgReg4IN_322, F(1)=>ImgReg4IN_321, F(0)=>
      ImgReg4IN_320);
   loop3_20_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_351_EXMPLR, D(14)=>OutputImg5_350_EXMPLR, D(13)=>
      OutputImg5_349_EXMPLR, D(12)=>OutputImg5_348_EXMPLR, D(11)=>
      OutputImg5_347_EXMPLR, D(10)=>OutputImg5_346_EXMPLR, D(9)=>
      OutputImg5_345_EXMPLR, D(8)=>OutputImg5_344_EXMPLR, D(7)=>
      OutputImg5_343_EXMPLR, D(6)=>OutputImg5_342_EXMPLR, D(5)=>
      OutputImg5_341_EXMPLR, D(4)=>OutputImg5_340_EXMPLR, D(3)=>
      OutputImg5_339_EXMPLR, D(2)=>OutputImg5_338_EXMPLR, D(1)=>
      OutputImg5_337_EXMPLR, D(0)=>OutputImg5_336_EXMPLR, EN=>nx23700, F(15)
      =>ImgReg5IN_335, F(14)=>ImgReg5IN_334, F(13)=>ImgReg5IN_333, F(12)=>
      ImgReg5IN_332, F(11)=>ImgReg5IN_331, F(10)=>ImgReg5IN_330, F(9)=>
      ImgReg5IN_329, F(8)=>ImgReg5IN_328, F(7)=>ImgReg5IN_327, F(6)=>
      ImgReg5IN_326, F(5)=>ImgReg5IN_325, F(4)=>ImgReg5IN_324, F(3)=>
      ImgReg5IN_323, F(2)=>ImgReg5IN_322, F(1)=>ImgReg5IN_321, F(0)=>
      ImgReg5IN_320);
   loop3_20_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(335), 
      D(14)=>DATA(334), D(13)=>DATA(333), D(12)=>DATA(332), D(11)=>DATA(331), 
      D(10)=>DATA(330), D(9)=>DATA(329), D(8)=>DATA(328), D(7)=>DATA(327), 
      D(6)=>DATA(326), D(5)=>DATA(325), D(4)=>DATA(324), D(3)=>DATA(323), 
      D(2)=>DATA(322), D(1)=>DATA(321), D(0)=>DATA(320), EN=>nx23658, F(15)
      =>ImgReg0IN_335, F(14)=>ImgReg0IN_334, F(13)=>ImgReg0IN_333, F(12)=>
      ImgReg0IN_332, F(11)=>ImgReg0IN_331, F(10)=>ImgReg0IN_330, F(9)=>
      ImgReg0IN_329, F(8)=>ImgReg0IN_328, F(7)=>ImgReg0IN_327, F(6)=>
      ImgReg0IN_326, F(5)=>ImgReg0IN_325, F(4)=>ImgReg0IN_324, F(3)=>
      ImgReg0IN_323, F(2)=>ImgReg0IN_322, F(1)=>ImgReg0IN_321, F(0)=>
      ImgReg0IN_320);
   loop3_20_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(335), 
      D(14)=>DATA(334), D(13)=>DATA(333), D(12)=>DATA(332), D(11)=>DATA(331), 
      D(10)=>DATA(330), D(9)=>DATA(329), D(8)=>DATA(328), D(7)=>DATA(327), 
      D(6)=>DATA(326), D(5)=>DATA(325), D(4)=>DATA(324), D(3)=>DATA(323), 
      D(2)=>DATA(322), D(1)=>DATA(321), D(0)=>DATA(320), EN=>nx23646, F(15)
      =>ImgReg1IN_335, F(14)=>ImgReg1IN_334, F(13)=>ImgReg1IN_333, F(12)=>
      ImgReg1IN_332, F(11)=>ImgReg1IN_331, F(10)=>ImgReg1IN_330, F(9)=>
      ImgReg1IN_329, F(8)=>ImgReg1IN_328, F(7)=>ImgReg1IN_327, F(6)=>
      ImgReg1IN_326, F(5)=>ImgReg1IN_325, F(4)=>ImgReg1IN_324, F(3)=>
      ImgReg1IN_323, F(2)=>ImgReg1IN_322, F(1)=>ImgReg1IN_321, F(0)=>
      ImgReg1IN_320);
   loop3_20_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(335), 
      D(14)=>DATA(334), D(13)=>DATA(333), D(12)=>DATA(332), D(11)=>DATA(331), 
      D(10)=>DATA(330), D(9)=>DATA(329), D(8)=>DATA(328), D(7)=>DATA(327), 
      D(6)=>DATA(326), D(5)=>DATA(325), D(4)=>DATA(324), D(3)=>DATA(323), 
      D(2)=>DATA(322), D(1)=>DATA(321), D(0)=>DATA(320), EN=>nx23634, F(15)
      =>ImgReg2IN_335, F(14)=>ImgReg2IN_334, F(13)=>ImgReg2IN_333, F(12)=>
      ImgReg2IN_332, F(11)=>ImgReg2IN_331, F(10)=>ImgReg2IN_330, F(9)=>
      ImgReg2IN_329, F(8)=>ImgReg2IN_328, F(7)=>ImgReg2IN_327, F(6)=>
      ImgReg2IN_326, F(5)=>ImgReg2IN_325, F(4)=>ImgReg2IN_324, F(3)=>
      ImgReg2IN_323, F(2)=>ImgReg2IN_322, F(1)=>ImgReg2IN_321, F(0)=>
      ImgReg2IN_320);
   loop3_20_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(335), 
      D(14)=>DATA(334), D(13)=>DATA(333), D(12)=>DATA(332), D(11)=>DATA(331), 
      D(10)=>DATA(330), D(9)=>DATA(329), D(8)=>DATA(328), D(7)=>DATA(327), 
      D(6)=>DATA(326), D(5)=>DATA(325), D(4)=>DATA(324), D(3)=>DATA(323), 
      D(2)=>DATA(322), D(1)=>DATA(321), D(0)=>DATA(320), EN=>nx23622, F(15)
      =>ImgReg3IN_335, F(14)=>ImgReg3IN_334, F(13)=>ImgReg3IN_333, F(12)=>
      ImgReg3IN_332, F(11)=>ImgReg3IN_331, F(10)=>ImgReg3IN_330, F(9)=>
      ImgReg3IN_329, F(8)=>ImgReg3IN_328, F(7)=>ImgReg3IN_327, F(6)=>
      ImgReg3IN_326, F(5)=>ImgReg3IN_325, F(4)=>ImgReg3IN_324, F(3)=>
      ImgReg3IN_323, F(2)=>ImgReg3IN_322, F(1)=>ImgReg3IN_321, F(0)=>
      ImgReg3IN_320);
   loop3_20_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(335), 
      D(14)=>DATA(334), D(13)=>DATA(333), D(12)=>DATA(332), D(11)=>DATA(331), 
      D(10)=>DATA(330), D(9)=>DATA(329), D(8)=>DATA(328), D(7)=>DATA(327), 
      D(6)=>DATA(326), D(5)=>DATA(325), D(4)=>DATA(324), D(3)=>DATA(323), 
      D(2)=>DATA(322), D(1)=>DATA(321), D(0)=>DATA(320), EN=>nx23610, F(15)
      =>ImgReg4IN_335, F(14)=>ImgReg4IN_334, F(13)=>ImgReg4IN_333, F(12)=>
      ImgReg4IN_332, F(11)=>ImgReg4IN_331, F(10)=>ImgReg4IN_330, F(9)=>
      ImgReg4IN_329, F(8)=>ImgReg4IN_328, F(7)=>ImgReg4IN_327, F(6)=>
      ImgReg4IN_326, F(5)=>ImgReg4IN_325, F(4)=>ImgReg4IN_324, F(3)=>
      ImgReg4IN_323, F(2)=>ImgReg4IN_322, F(1)=>ImgReg4IN_321, F(0)=>
      ImgReg4IN_320);
   loop3_20_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(335), 
      D(14)=>DATA(334), D(13)=>DATA(333), D(12)=>DATA(332), D(11)=>DATA(331), 
      D(10)=>DATA(330), D(9)=>DATA(329), D(8)=>DATA(328), D(7)=>DATA(327), 
      D(6)=>DATA(326), D(5)=>DATA(325), D(4)=>DATA(324), D(3)=>DATA(323), 
      D(2)=>DATA(322), D(1)=>DATA(321), D(0)=>DATA(320), EN=>nx23598, F(15)
      =>ImgReg5IN_335, F(14)=>ImgReg5IN_334, F(13)=>ImgReg5IN_333, F(12)=>
      ImgReg5IN_332, F(11)=>ImgReg5IN_331, F(10)=>ImgReg5IN_330, F(9)=>
      ImgReg5IN_329, F(8)=>ImgReg5IN_328, F(7)=>ImgReg5IN_327, F(6)=>
      ImgReg5IN_326, F(5)=>ImgReg5IN_325, F(4)=>ImgReg5IN_324, F(3)=>
      ImgReg5IN_323, F(2)=>ImgReg5IN_322, F(1)=>ImgReg5IN_321, F(0)=>
      ImgReg5IN_320);
   loop3_20_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_335_EXMPLR, D(14)=>OutputImg1_334_EXMPLR, D(13)=>
      OutputImg1_333_EXMPLR, D(12)=>OutputImg1_332_EXMPLR, D(11)=>
      OutputImg1_331_EXMPLR, D(10)=>OutputImg1_330_EXMPLR, D(9)=>
      OutputImg1_329_EXMPLR, D(8)=>OutputImg1_328_EXMPLR, D(7)=>
      OutputImg1_327_EXMPLR, D(6)=>OutputImg1_326_EXMPLR, D(5)=>
      OutputImg1_325_EXMPLR, D(4)=>OutputImg1_324_EXMPLR, D(3)=>
      OutputImg1_323_EXMPLR, D(2)=>OutputImg1_322_EXMPLR, D(1)=>
      OutputImg1_321_EXMPLR, D(0)=>OutputImg1_320_EXMPLR, EN=>nx23814, F(15)
      =>ImgReg0IN_335, F(14)=>ImgReg0IN_334, F(13)=>ImgReg0IN_333, F(12)=>
      ImgReg0IN_332, F(11)=>ImgReg0IN_331, F(10)=>ImgReg0IN_330, F(9)=>
      ImgReg0IN_329, F(8)=>ImgReg0IN_328, F(7)=>ImgReg0IN_327, F(6)=>
      ImgReg0IN_326, F(5)=>ImgReg0IN_325, F(4)=>ImgReg0IN_324, F(3)=>
      ImgReg0IN_323, F(2)=>ImgReg0IN_322, F(1)=>ImgReg0IN_321, F(0)=>
      ImgReg0IN_320);
   loop3_20_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_335_EXMPLR, D(14)=>OutputImg2_334_EXMPLR, D(13)=>
      OutputImg2_333_EXMPLR, D(12)=>OutputImg2_332_EXMPLR, D(11)=>
      OutputImg2_331_EXMPLR, D(10)=>OutputImg2_330_EXMPLR, D(9)=>
      OutputImg2_329_EXMPLR, D(8)=>OutputImg2_328_EXMPLR, D(7)=>
      OutputImg2_327_EXMPLR, D(6)=>OutputImg2_326_EXMPLR, D(5)=>
      OutputImg2_325_EXMPLR, D(4)=>OutputImg2_324_EXMPLR, D(3)=>
      OutputImg2_323_EXMPLR, D(2)=>OutputImg2_322_EXMPLR, D(1)=>
      OutputImg2_321_EXMPLR, D(0)=>OutputImg2_320_EXMPLR, EN=>nx23814, F(15)
      =>ImgReg1IN_335, F(14)=>ImgReg1IN_334, F(13)=>ImgReg1IN_333, F(12)=>
      ImgReg1IN_332, F(11)=>ImgReg1IN_331, F(10)=>ImgReg1IN_330, F(9)=>
      ImgReg1IN_329, F(8)=>ImgReg1IN_328, F(7)=>ImgReg1IN_327, F(6)=>
      ImgReg1IN_326, F(5)=>ImgReg1IN_325, F(4)=>ImgReg1IN_324, F(3)=>
      ImgReg1IN_323, F(2)=>ImgReg1IN_322, F(1)=>ImgReg1IN_321, F(0)=>
      ImgReg1IN_320);
   loop3_20_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_335_EXMPLR, D(14)=>OutputImg3_334_EXMPLR, D(13)=>
      OutputImg3_333_EXMPLR, D(12)=>OutputImg3_332_EXMPLR, D(11)=>
      OutputImg3_331_EXMPLR, D(10)=>OutputImg3_330_EXMPLR, D(9)=>
      OutputImg3_329_EXMPLR, D(8)=>OutputImg3_328_EXMPLR, D(7)=>
      OutputImg3_327_EXMPLR, D(6)=>OutputImg3_326_EXMPLR, D(5)=>
      OutputImg3_325_EXMPLR, D(4)=>OutputImg3_324_EXMPLR, D(3)=>
      OutputImg3_323_EXMPLR, D(2)=>OutputImg3_322_EXMPLR, D(1)=>
      OutputImg3_321_EXMPLR, D(0)=>OutputImg3_320_EXMPLR, EN=>nx23814, F(15)
      =>ImgReg2IN_335, F(14)=>ImgReg2IN_334, F(13)=>ImgReg2IN_333, F(12)=>
      ImgReg2IN_332, F(11)=>ImgReg2IN_331, F(10)=>ImgReg2IN_330, F(9)=>
      ImgReg2IN_329, F(8)=>ImgReg2IN_328, F(7)=>ImgReg2IN_327, F(6)=>
      ImgReg2IN_326, F(5)=>ImgReg2IN_325, F(4)=>ImgReg2IN_324, F(3)=>
      ImgReg2IN_323, F(2)=>ImgReg2IN_322, F(1)=>ImgReg2IN_321, F(0)=>
      ImgReg2IN_320);
   loop3_20_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_335_EXMPLR, D(14)=>OutputImg4_334_EXMPLR, D(13)=>
      OutputImg4_333_EXMPLR, D(12)=>OutputImg4_332_EXMPLR, D(11)=>
      OutputImg4_331_EXMPLR, D(10)=>OutputImg4_330_EXMPLR, D(9)=>
      OutputImg4_329_EXMPLR, D(8)=>OutputImg4_328_EXMPLR, D(7)=>
      OutputImg4_327_EXMPLR, D(6)=>OutputImg4_326_EXMPLR, D(5)=>
      OutputImg4_325_EXMPLR, D(4)=>OutputImg4_324_EXMPLR, D(3)=>
      OutputImg4_323_EXMPLR, D(2)=>OutputImg4_322_EXMPLR, D(1)=>
      OutputImg4_321_EXMPLR, D(0)=>OutputImg4_320_EXMPLR, EN=>nx23814, F(15)
      =>ImgReg3IN_335, F(14)=>ImgReg3IN_334, F(13)=>ImgReg3IN_333, F(12)=>
      ImgReg3IN_332, F(11)=>ImgReg3IN_331, F(10)=>ImgReg3IN_330, F(9)=>
      ImgReg3IN_329, F(8)=>ImgReg3IN_328, F(7)=>ImgReg3IN_327, F(6)=>
      ImgReg3IN_326, F(5)=>ImgReg3IN_325, F(4)=>ImgReg3IN_324, F(3)=>
      ImgReg3IN_323, F(2)=>ImgReg3IN_322, F(1)=>ImgReg3IN_321, F(0)=>
      ImgReg3IN_320);
   loop3_20_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_335_EXMPLR, D(14)=>OutputImg5_334_EXMPLR, D(13)=>
      OutputImg5_333_EXMPLR, D(12)=>OutputImg5_332_EXMPLR, D(11)=>
      OutputImg5_331_EXMPLR, D(10)=>OutputImg5_330_EXMPLR, D(9)=>
      OutputImg5_329_EXMPLR, D(8)=>OutputImg5_328_EXMPLR, D(7)=>
      OutputImg5_327_EXMPLR, D(6)=>OutputImg5_326_EXMPLR, D(5)=>
      OutputImg5_325_EXMPLR, D(4)=>OutputImg5_324_EXMPLR, D(3)=>
      OutputImg5_323_EXMPLR, D(2)=>OutputImg5_322_EXMPLR, D(1)=>
      OutputImg5_321_EXMPLR, D(0)=>OutputImg5_320_EXMPLR, EN=>nx23814, F(15)
      =>ImgReg4IN_335, F(14)=>ImgReg4IN_334, F(13)=>ImgReg4IN_333, F(12)=>
      ImgReg4IN_332, F(11)=>ImgReg4IN_331, F(10)=>ImgReg4IN_330, F(9)=>
      ImgReg4IN_329, F(8)=>ImgReg4IN_328, F(7)=>ImgReg4IN_327, F(6)=>
      ImgReg4IN_326, F(5)=>ImgReg4IN_325, F(4)=>ImgReg4IN_324, F(3)=>
      ImgReg4IN_323, F(2)=>ImgReg4IN_322, F(1)=>ImgReg4IN_321, F(0)=>
      ImgReg4IN_320);
   loop3_20_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_335, D(14)=>
      ImgReg0IN_334, D(13)=>ImgReg0IN_333, D(12)=>ImgReg0IN_332, D(11)=>
      ImgReg0IN_331, D(10)=>ImgReg0IN_330, D(9)=>ImgReg0IN_329, D(8)=>
      ImgReg0IN_328, D(7)=>ImgReg0IN_327, D(6)=>ImgReg0IN_326, D(5)=>
      ImgReg0IN_325, D(4)=>ImgReg0IN_324, D(3)=>ImgReg0IN_323, D(2)=>
      ImgReg0IN_322, D(1)=>ImgReg0IN_321, D(0)=>ImgReg0IN_320, CLK=>nx23948, 
      RST=>RST, EN=>nx23722, Q(15)=>OutputImg0_335_EXMPLR, Q(14)=>
      OutputImg0_334_EXMPLR, Q(13)=>OutputImg0_333_EXMPLR, Q(12)=>
      OutputImg0_332_EXMPLR, Q(11)=>OutputImg0_331_EXMPLR, Q(10)=>
      OutputImg0_330_EXMPLR, Q(9)=>OutputImg0_329_EXMPLR, Q(8)=>
      OutputImg0_328_EXMPLR, Q(7)=>OutputImg0_327_EXMPLR, Q(6)=>
      OutputImg0_326_EXMPLR, Q(5)=>OutputImg0_325_EXMPLR, Q(4)=>
      OutputImg0_324_EXMPLR, Q(3)=>OutputImg0_323_EXMPLR, Q(2)=>
      OutputImg0_322_EXMPLR, Q(1)=>OutputImg0_321_EXMPLR, Q(0)=>
      OutputImg0_320_EXMPLR);
   loop3_20_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_335, D(14)=>
      ImgReg1IN_334, D(13)=>ImgReg1IN_333, D(12)=>ImgReg1IN_332, D(11)=>
      ImgReg1IN_331, D(10)=>ImgReg1IN_330, D(9)=>ImgReg1IN_329, D(8)=>
      ImgReg1IN_328, D(7)=>ImgReg1IN_327, D(6)=>ImgReg1IN_326, D(5)=>
      ImgReg1IN_325, D(4)=>ImgReg1IN_324, D(3)=>ImgReg1IN_323, D(2)=>
      ImgReg1IN_322, D(1)=>ImgReg1IN_321, D(0)=>ImgReg1IN_320, CLK=>nx23950, 
      RST=>RST, EN=>nx23732, Q(15)=>OutputImg1_335_EXMPLR, Q(14)=>
      OutputImg1_334_EXMPLR, Q(13)=>OutputImg1_333_EXMPLR, Q(12)=>
      OutputImg1_332_EXMPLR, Q(11)=>OutputImg1_331_EXMPLR, Q(10)=>
      OutputImg1_330_EXMPLR, Q(9)=>OutputImg1_329_EXMPLR, Q(8)=>
      OutputImg1_328_EXMPLR, Q(7)=>OutputImg1_327_EXMPLR, Q(6)=>
      OutputImg1_326_EXMPLR, Q(5)=>OutputImg1_325_EXMPLR, Q(4)=>
      OutputImg1_324_EXMPLR, Q(3)=>OutputImg1_323_EXMPLR, Q(2)=>
      OutputImg1_322_EXMPLR, Q(1)=>OutputImg1_321_EXMPLR, Q(0)=>
      OutputImg1_320_EXMPLR);
   loop3_20_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_335, D(14)=>
      ImgReg2IN_334, D(13)=>ImgReg2IN_333, D(12)=>ImgReg2IN_332, D(11)=>
      ImgReg2IN_331, D(10)=>ImgReg2IN_330, D(9)=>ImgReg2IN_329, D(8)=>
      ImgReg2IN_328, D(7)=>ImgReg2IN_327, D(6)=>ImgReg2IN_326, D(5)=>
      ImgReg2IN_325, D(4)=>ImgReg2IN_324, D(3)=>ImgReg2IN_323, D(2)=>
      ImgReg2IN_322, D(1)=>ImgReg2IN_321, D(0)=>ImgReg2IN_320, CLK=>nx23950, 
      RST=>RST, EN=>nx23742, Q(15)=>OutputImg2_335_EXMPLR, Q(14)=>
      OutputImg2_334_EXMPLR, Q(13)=>OutputImg2_333_EXMPLR, Q(12)=>
      OutputImg2_332_EXMPLR, Q(11)=>OutputImg2_331_EXMPLR, Q(10)=>
      OutputImg2_330_EXMPLR, Q(9)=>OutputImg2_329_EXMPLR, Q(8)=>
      OutputImg2_328_EXMPLR, Q(7)=>OutputImg2_327_EXMPLR, Q(6)=>
      OutputImg2_326_EXMPLR, Q(5)=>OutputImg2_325_EXMPLR, Q(4)=>
      OutputImg2_324_EXMPLR, Q(3)=>OutputImg2_323_EXMPLR, Q(2)=>
      OutputImg2_322_EXMPLR, Q(1)=>OutputImg2_321_EXMPLR, Q(0)=>
      OutputImg2_320_EXMPLR);
   loop3_20_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_335, D(14)=>
      ImgReg3IN_334, D(13)=>ImgReg3IN_333, D(12)=>ImgReg3IN_332, D(11)=>
      ImgReg3IN_331, D(10)=>ImgReg3IN_330, D(9)=>ImgReg3IN_329, D(8)=>
      ImgReg3IN_328, D(7)=>ImgReg3IN_327, D(6)=>ImgReg3IN_326, D(5)=>
      ImgReg3IN_325, D(4)=>ImgReg3IN_324, D(3)=>ImgReg3IN_323, D(2)=>
      ImgReg3IN_322, D(1)=>ImgReg3IN_321, D(0)=>ImgReg3IN_320, CLK=>nx23952, 
      RST=>RST, EN=>nx23752, Q(15)=>OutputImg3_335_EXMPLR, Q(14)=>
      OutputImg3_334_EXMPLR, Q(13)=>OutputImg3_333_EXMPLR, Q(12)=>
      OutputImg3_332_EXMPLR, Q(11)=>OutputImg3_331_EXMPLR, Q(10)=>
      OutputImg3_330_EXMPLR, Q(9)=>OutputImg3_329_EXMPLR, Q(8)=>
      OutputImg3_328_EXMPLR, Q(7)=>OutputImg3_327_EXMPLR, Q(6)=>
      OutputImg3_326_EXMPLR, Q(5)=>OutputImg3_325_EXMPLR, Q(4)=>
      OutputImg3_324_EXMPLR, Q(3)=>OutputImg3_323_EXMPLR, Q(2)=>
      OutputImg3_322_EXMPLR, Q(1)=>OutputImg3_321_EXMPLR, Q(0)=>
      OutputImg3_320_EXMPLR);
   loop3_20_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_335, D(14)=>
      ImgReg4IN_334, D(13)=>ImgReg4IN_333, D(12)=>ImgReg4IN_332, D(11)=>
      ImgReg4IN_331, D(10)=>ImgReg4IN_330, D(9)=>ImgReg4IN_329, D(8)=>
      ImgReg4IN_328, D(7)=>ImgReg4IN_327, D(6)=>ImgReg4IN_326, D(5)=>
      ImgReg4IN_325, D(4)=>ImgReg4IN_324, D(3)=>ImgReg4IN_323, D(2)=>
      ImgReg4IN_322, D(1)=>ImgReg4IN_321, D(0)=>ImgReg4IN_320, CLK=>nx23952, 
      RST=>RST, EN=>nx23762, Q(15)=>OutputImg4_335_EXMPLR, Q(14)=>
      OutputImg4_334_EXMPLR, Q(13)=>OutputImg4_333_EXMPLR, Q(12)=>
      OutputImg4_332_EXMPLR, Q(11)=>OutputImg4_331_EXMPLR, Q(10)=>
      OutputImg4_330_EXMPLR, Q(9)=>OutputImg4_329_EXMPLR, Q(8)=>
      OutputImg4_328_EXMPLR, Q(7)=>OutputImg4_327_EXMPLR, Q(6)=>
      OutputImg4_326_EXMPLR, Q(5)=>OutputImg4_325_EXMPLR, Q(4)=>
      OutputImg4_324_EXMPLR, Q(3)=>OutputImg4_323_EXMPLR, Q(2)=>
      OutputImg4_322_EXMPLR, Q(1)=>OutputImg4_321_EXMPLR, Q(0)=>
      OutputImg4_320_EXMPLR);
   loop3_20_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_335, D(14)=>
      ImgReg5IN_334, D(13)=>ImgReg5IN_333, D(12)=>ImgReg5IN_332, D(11)=>
      ImgReg5IN_331, D(10)=>ImgReg5IN_330, D(9)=>ImgReg5IN_329, D(8)=>
      ImgReg5IN_328, D(7)=>ImgReg5IN_327, D(6)=>ImgReg5IN_326, D(5)=>
      ImgReg5IN_325, D(4)=>ImgReg5IN_324, D(3)=>ImgReg5IN_323, D(2)=>
      ImgReg5IN_322, D(1)=>ImgReg5IN_321, D(0)=>ImgReg5IN_320, CLK=>nx23954, 
      RST=>RST, EN=>nx23772, Q(15)=>OutputImg5_335_EXMPLR, Q(14)=>
      OutputImg5_334_EXMPLR, Q(13)=>OutputImg5_333_EXMPLR, Q(12)=>
      OutputImg5_332_EXMPLR, Q(11)=>OutputImg5_331_EXMPLR, Q(10)=>
      OutputImg5_330_EXMPLR, Q(9)=>OutputImg5_329_EXMPLR, Q(8)=>
      OutputImg5_328_EXMPLR, Q(7)=>OutputImg5_327_EXMPLR, Q(6)=>
      OutputImg5_326_EXMPLR, Q(5)=>OutputImg5_325_EXMPLR, Q(4)=>
      OutputImg5_324_EXMPLR, Q(3)=>OutputImg5_323_EXMPLR, Q(2)=>
      OutputImg5_322_EXMPLR, Q(1)=>OutputImg5_321_EXMPLR, Q(0)=>
      OutputImg5_320_EXMPLR);
   loop3_21_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_367_EXMPLR, D(14)=>OutputImg0_366_EXMPLR, D(13)=>
      OutputImg0_365_EXMPLR, D(12)=>OutputImg0_364_EXMPLR, D(11)=>
      OutputImg0_363_EXMPLR, D(10)=>OutputImg0_362_EXMPLR, D(9)=>
      OutputImg0_361_EXMPLR, D(8)=>OutputImg0_360_EXMPLR, D(7)=>
      OutputImg0_359_EXMPLR, D(6)=>OutputImg0_358_EXMPLR, D(5)=>
      OutputImg0_357_EXMPLR, D(4)=>OutputImg0_356_EXMPLR, D(3)=>
      OutputImg0_355_EXMPLR, D(2)=>OutputImg0_354_EXMPLR, D(1)=>
      OutputImg0_353_EXMPLR, D(0)=>OutputImg0_352_EXMPLR, EN=>nx23702, F(15)
      =>ImgReg0IN_351, F(14)=>ImgReg0IN_350, F(13)=>ImgReg0IN_349, F(12)=>
      ImgReg0IN_348, F(11)=>ImgReg0IN_347, F(10)=>ImgReg0IN_346, F(9)=>
      ImgReg0IN_345, F(8)=>ImgReg0IN_344, F(7)=>ImgReg0IN_343, F(6)=>
      ImgReg0IN_342, F(5)=>ImgReg0IN_341, F(4)=>ImgReg0IN_340, F(3)=>
      ImgReg0IN_339, F(2)=>ImgReg0IN_338, F(1)=>ImgReg0IN_337, F(0)=>
      ImgReg0IN_336);
   loop3_21_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_367_EXMPLR, D(14)=>OutputImg1_366_EXMPLR, D(13)=>
      OutputImg1_365_EXMPLR, D(12)=>OutputImg1_364_EXMPLR, D(11)=>
      OutputImg1_363_EXMPLR, D(10)=>OutputImg1_362_EXMPLR, D(9)=>
      OutputImg1_361_EXMPLR, D(8)=>OutputImg1_360_EXMPLR, D(7)=>
      OutputImg1_359_EXMPLR, D(6)=>OutputImg1_358_EXMPLR, D(5)=>
      OutputImg1_357_EXMPLR, D(4)=>OutputImg1_356_EXMPLR, D(3)=>
      OutputImg1_355_EXMPLR, D(2)=>OutputImg1_354_EXMPLR, D(1)=>
      OutputImg1_353_EXMPLR, D(0)=>OutputImg1_352_EXMPLR, EN=>nx23702, F(15)
      =>ImgReg1IN_351, F(14)=>ImgReg1IN_350, F(13)=>ImgReg1IN_349, F(12)=>
      ImgReg1IN_348, F(11)=>ImgReg1IN_347, F(10)=>ImgReg1IN_346, F(9)=>
      ImgReg1IN_345, F(8)=>ImgReg1IN_344, F(7)=>ImgReg1IN_343, F(6)=>
      ImgReg1IN_342, F(5)=>ImgReg1IN_341, F(4)=>ImgReg1IN_340, F(3)=>
      ImgReg1IN_339, F(2)=>ImgReg1IN_338, F(1)=>ImgReg1IN_337, F(0)=>
      ImgReg1IN_336);
   loop3_21_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_367_EXMPLR, D(14)=>OutputImg2_366_EXMPLR, D(13)=>
      OutputImg2_365_EXMPLR, D(12)=>OutputImg2_364_EXMPLR, D(11)=>
      OutputImg2_363_EXMPLR, D(10)=>OutputImg2_362_EXMPLR, D(9)=>
      OutputImg2_361_EXMPLR, D(8)=>OutputImg2_360_EXMPLR, D(7)=>
      OutputImg2_359_EXMPLR, D(6)=>OutputImg2_358_EXMPLR, D(5)=>
      OutputImg2_357_EXMPLR, D(4)=>OutputImg2_356_EXMPLR, D(3)=>
      OutputImg2_355_EXMPLR, D(2)=>OutputImg2_354_EXMPLR, D(1)=>
      OutputImg2_353_EXMPLR, D(0)=>OutputImg2_352_EXMPLR, EN=>nx23702, F(15)
      =>ImgReg2IN_351, F(14)=>ImgReg2IN_350, F(13)=>ImgReg2IN_349, F(12)=>
      ImgReg2IN_348, F(11)=>ImgReg2IN_347, F(10)=>ImgReg2IN_346, F(9)=>
      ImgReg2IN_345, F(8)=>ImgReg2IN_344, F(7)=>ImgReg2IN_343, F(6)=>
      ImgReg2IN_342, F(5)=>ImgReg2IN_341, F(4)=>ImgReg2IN_340, F(3)=>
      ImgReg2IN_339, F(2)=>ImgReg2IN_338, F(1)=>ImgReg2IN_337, F(0)=>
      ImgReg2IN_336);
   loop3_21_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_367_EXMPLR, D(14)=>OutputImg3_366_EXMPLR, D(13)=>
      OutputImg3_365_EXMPLR, D(12)=>OutputImg3_364_EXMPLR, D(11)=>
      OutputImg3_363_EXMPLR, D(10)=>OutputImg3_362_EXMPLR, D(9)=>
      OutputImg3_361_EXMPLR, D(8)=>OutputImg3_360_EXMPLR, D(7)=>
      OutputImg3_359_EXMPLR, D(6)=>OutputImg3_358_EXMPLR, D(5)=>
      OutputImg3_357_EXMPLR, D(4)=>OutputImg3_356_EXMPLR, D(3)=>
      OutputImg3_355_EXMPLR, D(2)=>OutputImg3_354_EXMPLR, D(1)=>
      OutputImg3_353_EXMPLR, D(0)=>OutputImg3_352_EXMPLR, EN=>nx23702, F(15)
      =>ImgReg3IN_351, F(14)=>ImgReg3IN_350, F(13)=>ImgReg3IN_349, F(12)=>
      ImgReg3IN_348, F(11)=>ImgReg3IN_347, F(10)=>ImgReg3IN_346, F(9)=>
      ImgReg3IN_345, F(8)=>ImgReg3IN_344, F(7)=>ImgReg3IN_343, F(6)=>
      ImgReg3IN_342, F(5)=>ImgReg3IN_341, F(4)=>ImgReg3IN_340, F(3)=>
      ImgReg3IN_339, F(2)=>ImgReg3IN_338, F(1)=>ImgReg3IN_337, F(0)=>
      ImgReg3IN_336);
   loop3_21_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_367_EXMPLR, D(14)=>OutputImg4_366_EXMPLR, D(13)=>
      OutputImg4_365_EXMPLR, D(12)=>OutputImg4_364_EXMPLR, D(11)=>
      OutputImg4_363_EXMPLR, D(10)=>OutputImg4_362_EXMPLR, D(9)=>
      OutputImg4_361_EXMPLR, D(8)=>OutputImg4_360_EXMPLR, D(7)=>
      OutputImg4_359_EXMPLR, D(6)=>OutputImg4_358_EXMPLR, D(5)=>
      OutputImg4_357_EXMPLR, D(4)=>OutputImg4_356_EXMPLR, D(3)=>
      OutputImg4_355_EXMPLR, D(2)=>OutputImg4_354_EXMPLR, D(1)=>
      OutputImg4_353_EXMPLR, D(0)=>OutputImg4_352_EXMPLR, EN=>nx23702, F(15)
      =>ImgReg4IN_351, F(14)=>ImgReg4IN_350, F(13)=>ImgReg4IN_349, F(12)=>
      ImgReg4IN_348, F(11)=>ImgReg4IN_347, F(10)=>ImgReg4IN_346, F(9)=>
      ImgReg4IN_345, F(8)=>ImgReg4IN_344, F(7)=>ImgReg4IN_343, F(6)=>
      ImgReg4IN_342, F(5)=>ImgReg4IN_341, F(4)=>ImgReg4IN_340, F(3)=>
      ImgReg4IN_339, F(2)=>ImgReg4IN_338, F(1)=>ImgReg4IN_337, F(0)=>
      ImgReg4IN_336);
   loop3_21_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_367_EXMPLR, D(14)=>OutputImg5_366_EXMPLR, D(13)=>
      OutputImg5_365_EXMPLR, D(12)=>OutputImg5_364_EXMPLR, D(11)=>
      OutputImg5_363_EXMPLR, D(10)=>OutputImg5_362_EXMPLR, D(9)=>
      OutputImg5_361_EXMPLR, D(8)=>OutputImg5_360_EXMPLR, D(7)=>
      OutputImg5_359_EXMPLR, D(6)=>OutputImg5_358_EXMPLR, D(5)=>
      OutputImg5_357_EXMPLR, D(4)=>OutputImg5_356_EXMPLR, D(3)=>
      OutputImg5_355_EXMPLR, D(2)=>OutputImg5_354_EXMPLR, D(1)=>
      OutputImg5_353_EXMPLR, D(0)=>OutputImg5_352_EXMPLR, EN=>nx23702, F(15)
      =>ImgReg5IN_351, F(14)=>ImgReg5IN_350, F(13)=>ImgReg5IN_349, F(12)=>
      ImgReg5IN_348, F(11)=>ImgReg5IN_347, F(10)=>ImgReg5IN_346, F(9)=>
      ImgReg5IN_345, F(8)=>ImgReg5IN_344, F(7)=>ImgReg5IN_343, F(6)=>
      ImgReg5IN_342, F(5)=>ImgReg5IN_341, F(4)=>ImgReg5IN_340, F(3)=>
      ImgReg5IN_339, F(2)=>ImgReg5IN_338, F(1)=>ImgReg5IN_337, F(0)=>
      ImgReg5IN_336);
   loop3_21_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(351), 
      D(14)=>DATA(350), D(13)=>DATA(349), D(12)=>DATA(348), D(11)=>DATA(347), 
      D(10)=>DATA(346), D(9)=>DATA(345), D(8)=>DATA(344), D(7)=>DATA(343), 
      D(6)=>DATA(342), D(5)=>DATA(341), D(4)=>DATA(340), D(3)=>DATA(339), 
      D(2)=>DATA(338), D(1)=>DATA(337), D(0)=>DATA(336), EN=>nx23660, F(15)
      =>ImgReg0IN_351, F(14)=>ImgReg0IN_350, F(13)=>ImgReg0IN_349, F(12)=>
      ImgReg0IN_348, F(11)=>ImgReg0IN_347, F(10)=>ImgReg0IN_346, F(9)=>
      ImgReg0IN_345, F(8)=>ImgReg0IN_344, F(7)=>ImgReg0IN_343, F(6)=>
      ImgReg0IN_342, F(5)=>ImgReg0IN_341, F(4)=>ImgReg0IN_340, F(3)=>
      ImgReg0IN_339, F(2)=>ImgReg0IN_338, F(1)=>ImgReg0IN_337, F(0)=>
      ImgReg0IN_336);
   loop3_21_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(351), 
      D(14)=>DATA(350), D(13)=>DATA(349), D(12)=>DATA(348), D(11)=>DATA(347), 
      D(10)=>DATA(346), D(9)=>DATA(345), D(8)=>DATA(344), D(7)=>DATA(343), 
      D(6)=>DATA(342), D(5)=>DATA(341), D(4)=>DATA(340), D(3)=>DATA(339), 
      D(2)=>DATA(338), D(1)=>DATA(337), D(0)=>DATA(336), EN=>nx23648, F(15)
      =>ImgReg1IN_351, F(14)=>ImgReg1IN_350, F(13)=>ImgReg1IN_349, F(12)=>
      ImgReg1IN_348, F(11)=>ImgReg1IN_347, F(10)=>ImgReg1IN_346, F(9)=>
      ImgReg1IN_345, F(8)=>ImgReg1IN_344, F(7)=>ImgReg1IN_343, F(6)=>
      ImgReg1IN_342, F(5)=>ImgReg1IN_341, F(4)=>ImgReg1IN_340, F(3)=>
      ImgReg1IN_339, F(2)=>ImgReg1IN_338, F(1)=>ImgReg1IN_337, F(0)=>
      ImgReg1IN_336);
   loop3_21_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(351), 
      D(14)=>DATA(350), D(13)=>DATA(349), D(12)=>DATA(348), D(11)=>DATA(347), 
      D(10)=>DATA(346), D(9)=>DATA(345), D(8)=>DATA(344), D(7)=>DATA(343), 
      D(6)=>DATA(342), D(5)=>DATA(341), D(4)=>DATA(340), D(3)=>DATA(339), 
      D(2)=>DATA(338), D(1)=>DATA(337), D(0)=>DATA(336), EN=>nx23636, F(15)
      =>ImgReg2IN_351, F(14)=>ImgReg2IN_350, F(13)=>ImgReg2IN_349, F(12)=>
      ImgReg2IN_348, F(11)=>ImgReg2IN_347, F(10)=>ImgReg2IN_346, F(9)=>
      ImgReg2IN_345, F(8)=>ImgReg2IN_344, F(7)=>ImgReg2IN_343, F(6)=>
      ImgReg2IN_342, F(5)=>ImgReg2IN_341, F(4)=>ImgReg2IN_340, F(3)=>
      ImgReg2IN_339, F(2)=>ImgReg2IN_338, F(1)=>ImgReg2IN_337, F(0)=>
      ImgReg2IN_336);
   loop3_21_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(351), 
      D(14)=>DATA(350), D(13)=>DATA(349), D(12)=>DATA(348), D(11)=>DATA(347), 
      D(10)=>DATA(346), D(9)=>DATA(345), D(8)=>DATA(344), D(7)=>DATA(343), 
      D(6)=>DATA(342), D(5)=>DATA(341), D(4)=>DATA(340), D(3)=>DATA(339), 
      D(2)=>DATA(338), D(1)=>DATA(337), D(0)=>DATA(336), EN=>nx23624, F(15)
      =>ImgReg3IN_351, F(14)=>ImgReg3IN_350, F(13)=>ImgReg3IN_349, F(12)=>
      ImgReg3IN_348, F(11)=>ImgReg3IN_347, F(10)=>ImgReg3IN_346, F(9)=>
      ImgReg3IN_345, F(8)=>ImgReg3IN_344, F(7)=>ImgReg3IN_343, F(6)=>
      ImgReg3IN_342, F(5)=>ImgReg3IN_341, F(4)=>ImgReg3IN_340, F(3)=>
      ImgReg3IN_339, F(2)=>ImgReg3IN_338, F(1)=>ImgReg3IN_337, F(0)=>
      ImgReg3IN_336);
   loop3_21_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(351), 
      D(14)=>DATA(350), D(13)=>DATA(349), D(12)=>DATA(348), D(11)=>DATA(347), 
      D(10)=>DATA(346), D(9)=>DATA(345), D(8)=>DATA(344), D(7)=>DATA(343), 
      D(6)=>DATA(342), D(5)=>DATA(341), D(4)=>DATA(340), D(3)=>DATA(339), 
      D(2)=>DATA(338), D(1)=>DATA(337), D(0)=>DATA(336), EN=>nx23612, F(15)
      =>ImgReg4IN_351, F(14)=>ImgReg4IN_350, F(13)=>ImgReg4IN_349, F(12)=>
      ImgReg4IN_348, F(11)=>ImgReg4IN_347, F(10)=>ImgReg4IN_346, F(9)=>
      ImgReg4IN_345, F(8)=>ImgReg4IN_344, F(7)=>ImgReg4IN_343, F(6)=>
      ImgReg4IN_342, F(5)=>ImgReg4IN_341, F(4)=>ImgReg4IN_340, F(3)=>
      ImgReg4IN_339, F(2)=>ImgReg4IN_338, F(1)=>ImgReg4IN_337, F(0)=>
      ImgReg4IN_336);
   loop3_21_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(351), 
      D(14)=>DATA(350), D(13)=>DATA(349), D(12)=>DATA(348), D(11)=>DATA(347), 
      D(10)=>DATA(346), D(9)=>DATA(345), D(8)=>DATA(344), D(7)=>DATA(343), 
      D(6)=>DATA(342), D(5)=>DATA(341), D(4)=>DATA(340), D(3)=>DATA(339), 
      D(2)=>DATA(338), D(1)=>DATA(337), D(0)=>DATA(336), EN=>nx23600, F(15)
      =>ImgReg5IN_351, F(14)=>ImgReg5IN_350, F(13)=>ImgReg5IN_349, F(12)=>
      ImgReg5IN_348, F(11)=>ImgReg5IN_347, F(10)=>ImgReg5IN_346, F(9)=>
      ImgReg5IN_345, F(8)=>ImgReg5IN_344, F(7)=>ImgReg5IN_343, F(6)=>
      ImgReg5IN_342, F(5)=>ImgReg5IN_341, F(4)=>ImgReg5IN_340, F(3)=>
      ImgReg5IN_339, F(2)=>ImgReg5IN_338, F(1)=>ImgReg5IN_337, F(0)=>
      ImgReg5IN_336);
   loop3_21_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_351_EXMPLR, D(14)=>OutputImg1_350_EXMPLR, D(13)=>
      OutputImg1_349_EXMPLR, D(12)=>OutputImg1_348_EXMPLR, D(11)=>
      OutputImg1_347_EXMPLR, D(10)=>OutputImg1_346_EXMPLR, D(9)=>
      OutputImg1_345_EXMPLR, D(8)=>OutputImg1_344_EXMPLR, D(7)=>
      OutputImg1_343_EXMPLR, D(6)=>OutputImg1_342_EXMPLR, D(5)=>
      OutputImg1_341_EXMPLR, D(4)=>OutputImg1_340_EXMPLR, D(3)=>
      OutputImg1_339_EXMPLR, D(2)=>OutputImg1_338_EXMPLR, D(1)=>
      OutputImg1_337_EXMPLR, D(0)=>OutputImg1_336_EXMPLR, EN=>nx23816, F(15)
      =>ImgReg0IN_351, F(14)=>ImgReg0IN_350, F(13)=>ImgReg0IN_349, F(12)=>
      ImgReg0IN_348, F(11)=>ImgReg0IN_347, F(10)=>ImgReg0IN_346, F(9)=>
      ImgReg0IN_345, F(8)=>ImgReg0IN_344, F(7)=>ImgReg0IN_343, F(6)=>
      ImgReg0IN_342, F(5)=>ImgReg0IN_341, F(4)=>ImgReg0IN_340, F(3)=>
      ImgReg0IN_339, F(2)=>ImgReg0IN_338, F(1)=>ImgReg0IN_337, F(0)=>
      ImgReg0IN_336);
   loop3_21_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_351_EXMPLR, D(14)=>OutputImg2_350_EXMPLR, D(13)=>
      OutputImg2_349_EXMPLR, D(12)=>OutputImg2_348_EXMPLR, D(11)=>
      OutputImg2_347_EXMPLR, D(10)=>OutputImg2_346_EXMPLR, D(9)=>
      OutputImg2_345_EXMPLR, D(8)=>OutputImg2_344_EXMPLR, D(7)=>
      OutputImg2_343_EXMPLR, D(6)=>OutputImg2_342_EXMPLR, D(5)=>
      OutputImg2_341_EXMPLR, D(4)=>OutputImg2_340_EXMPLR, D(3)=>
      OutputImg2_339_EXMPLR, D(2)=>OutputImg2_338_EXMPLR, D(1)=>
      OutputImg2_337_EXMPLR, D(0)=>OutputImg2_336_EXMPLR, EN=>nx23816, F(15)
      =>ImgReg1IN_351, F(14)=>ImgReg1IN_350, F(13)=>ImgReg1IN_349, F(12)=>
      ImgReg1IN_348, F(11)=>ImgReg1IN_347, F(10)=>ImgReg1IN_346, F(9)=>
      ImgReg1IN_345, F(8)=>ImgReg1IN_344, F(7)=>ImgReg1IN_343, F(6)=>
      ImgReg1IN_342, F(5)=>ImgReg1IN_341, F(4)=>ImgReg1IN_340, F(3)=>
      ImgReg1IN_339, F(2)=>ImgReg1IN_338, F(1)=>ImgReg1IN_337, F(0)=>
      ImgReg1IN_336);
   loop3_21_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_351_EXMPLR, D(14)=>OutputImg3_350_EXMPLR, D(13)=>
      OutputImg3_349_EXMPLR, D(12)=>OutputImg3_348_EXMPLR, D(11)=>
      OutputImg3_347_EXMPLR, D(10)=>OutputImg3_346_EXMPLR, D(9)=>
      OutputImg3_345_EXMPLR, D(8)=>OutputImg3_344_EXMPLR, D(7)=>
      OutputImg3_343_EXMPLR, D(6)=>OutputImg3_342_EXMPLR, D(5)=>
      OutputImg3_341_EXMPLR, D(4)=>OutputImg3_340_EXMPLR, D(3)=>
      OutputImg3_339_EXMPLR, D(2)=>OutputImg3_338_EXMPLR, D(1)=>
      OutputImg3_337_EXMPLR, D(0)=>OutputImg3_336_EXMPLR, EN=>nx23816, F(15)
      =>ImgReg2IN_351, F(14)=>ImgReg2IN_350, F(13)=>ImgReg2IN_349, F(12)=>
      ImgReg2IN_348, F(11)=>ImgReg2IN_347, F(10)=>ImgReg2IN_346, F(9)=>
      ImgReg2IN_345, F(8)=>ImgReg2IN_344, F(7)=>ImgReg2IN_343, F(6)=>
      ImgReg2IN_342, F(5)=>ImgReg2IN_341, F(4)=>ImgReg2IN_340, F(3)=>
      ImgReg2IN_339, F(2)=>ImgReg2IN_338, F(1)=>ImgReg2IN_337, F(0)=>
      ImgReg2IN_336);
   loop3_21_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_351_EXMPLR, D(14)=>OutputImg4_350_EXMPLR, D(13)=>
      OutputImg4_349_EXMPLR, D(12)=>OutputImg4_348_EXMPLR, D(11)=>
      OutputImg4_347_EXMPLR, D(10)=>OutputImg4_346_EXMPLR, D(9)=>
      OutputImg4_345_EXMPLR, D(8)=>OutputImg4_344_EXMPLR, D(7)=>
      OutputImg4_343_EXMPLR, D(6)=>OutputImg4_342_EXMPLR, D(5)=>
      OutputImg4_341_EXMPLR, D(4)=>OutputImg4_340_EXMPLR, D(3)=>
      OutputImg4_339_EXMPLR, D(2)=>OutputImg4_338_EXMPLR, D(1)=>
      OutputImg4_337_EXMPLR, D(0)=>OutputImg4_336_EXMPLR, EN=>nx23816, F(15)
      =>ImgReg3IN_351, F(14)=>ImgReg3IN_350, F(13)=>ImgReg3IN_349, F(12)=>
      ImgReg3IN_348, F(11)=>ImgReg3IN_347, F(10)=>ImgReg3IN_346, F(9)=>
      ImgReg3IN_345, F(8)=>ImgReg3IN_344, F(7)=>ImgReg3IN_343, F(6)=>
      ImgReg3IN_342, F(5)=>ImgReg3IN_341, F(4)=>ImgReg3IN_340, F(3)=>
      ImgReg3IN_339, F(2)=>ImgReg3IN_338, F(1)=>ImgReg3IN_337, F(0)=>
      ImgReg3IN_336);
   loop3_21_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_351_EXMPLR, D(14)=>OutputImg5_350_EXMPLR, D(13)=>
      OutputImg5_349_EXMPLR, D(12)=>OutputImg5_348_EXMPLR, D(11)=>
      OutputImg5_347_EXMPLR, D(10)=>OutputImg5_346_EXMPLR, D(9)=>
      OutputImg5_345_EXMPLR, D(8)=>OutputImg5_344_EXMPLR, D(7)=>
      OutputImg5_343_EXMPLR, D(6)=>OutputImg5_342_EXMPLR, D(5)=>
      OutputImg5_341_EXMPLR, D(4)=>OutputImg5_340_EXMPLR, D(3)=>
      OutputImg5_339_EXMPLR, D(2)=>OutputImg5_338_EXMPLR, D(1)=>
      OutputImg5_337_EXMPLR, D(0)=>OutputImg5_336_EXMPLR, EN=>nx23816, F(15)
      =>ImgReg4IN_351, F(14)=>ImgReg4IN_350, F(13)=>ImgReg4IN_349, F(12)=>
      ImgReg4IN_348, F(11)=>ImgReg4IN_347, F(10)=>ImgReg4IN_346, F(9)=>
      ImgReg4IN_345, F(8)=>ImgReg4IN_344, F(7)=>ImgReg4IN_343, F(6)=>
      ImgReg4IN_342, F(5)=>ImgReg4IN_341, F(4)=>ImgReg4IN_340, F(3)=>
      ImgReg4IN_339, F(2)=>ImgReg4IN_338, F(1)=>ImgReg4IN_337, F(0)=>
      ImgReg4IN_336);
   loop3_21_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_351, D(14)=>
      ImgReg0IN_350, D(13)=>ImgReg0IN_349, D(12)=>ImgReg0IN_348, D(11)=>
      ImgReg0IN_347, D(10)=>ImgReg0IN_346, D(9)=>ImgReg0IN_345, D(8)=>
      ImgReg0IN_344, D(7)=>ImgReg0IN_343, D(6)=>ImgReg0IN_342, D(5)=>
      ImgReg0IN_341, D(4)=>ImgReg0IN_340, D(3)=>ImgReg0IN_339, D(2)=>
      ImgReg0IN_338, D(1)=>ImgReg0IN_337, D(0)=>ImgReg0IN_336, CLK=>nx23954, 
      RST=>RST, EN=>nx23724, Q(15)=>OutputImg0_351_EXMPLR, Q(14)=>
      OutputImg0_350_EXMPLR, Q(13)=>OutputImg0_349_EXMPLR, Q(12)=>
      OutputImg0_348_EXMPLR, Q(11)=>OutputImg0_347_EXMPLR, Q(10)=>
      OutputImg0_346_EXMPLR, Q(9)=>OutputImg0_345_EXMPLR, Q(8)=>
      OutputImg0_344_EXMPLR, Q(7)=>OutputImg0_343_EXMPLR, Q(6)=>
      OutputImg0_342_EXMPLR, Q(5)=>OutputImg0_341_EXMPLR, Q(4)=>
      OutputImg0_340_EXMPLR, Q(3)=>OutputImg0_339_EXMPLR, Q(2)=>
      OutputImg0_338_EXMPLR, Q(1)=>OutputImg0_337_EXMPLR, Q(0)=>
      OutputImg0_336_EXMPLR);
   loop3_21_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_351, D(14)=>
      ImgReg1IN_350, D(13)=>ImgReg1IN_349, D(12)=>ImgReg1IN_348, D(11)=>
      ImgReg1IN_347, D(10)=>ImgReg1IN_346, D(9)=>ImgReg1IN_345, D(8)=>
      ImgReg1IN_344, D(7)=>ImgReg1IN_343, D(6)=>ImgReg1IN_342, D(5)=>
      ImgReg1IN_341, D(4)=>ImgReg1IN_340, D(3)=>ImgReg1IN_339, D(2)=>
      ImgReg1IN_338, D(1)=>ImgReg1IN_337, D(0)=>ImgReg1IN_336, CLK=>nx23956, 
      RST=>RST, EN=>nx23734, Q(15)=>OutputImg1_351_EXMPLR, Q(14)=>
      OutputImg1_350_EXMPLR, Q(13)=>OutputImg1_349_EXMPLR, Q(12)=>
      OutputImg1_348_EXMPLR, Q(11)=>OutputImg1_347_EXMPLR, Q(10)=>
      OutputImg1_346_EXMPLR, Q(9)=>OutputImg1_345_EXMPLR, Q(8)=>
      OutputImg1_344_EXMPLR, Q(7)=>OutputImg1_343_EXMPLR, Q(6)=>
      OutputImg1_342_EXMPLR, Q(5)=>OutputImg1_341_EXMPLR, Q(4)=>
      OutputImg1_340_EXMPLR, Q(3)=>OutputImg1_339_EXMPLR, Q(2)=>
      OutputImg1_338_EXMPLR, Q(1)=>OutputImg1_337_EXMPLR, Q(0)=>
      OutputImg1_336_EXMPLR);
   loop3_21_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_351, D(14)=>
      ImgReg2IN_350, D(13)=>ImgReg2IN_349, D(12)=>ImgReg2IN_348, D(11)=>
      ImgReg2IN_347, D(10)=>ImgReg2IN_346, D(9)=>ImgReg2IN_345, D(8)=>
      ImgReg2IN_344, D(7)=>ImgReg2IN_343, D(6)=>ImgReg2IN_342, D(5)=>
      ImgReg2IN_341, D(4)=>ImgReg2IN_340, D(3)=>ImgReg2IN_339, D(2)=>
      ImgReg2IN_338, D(1)=>ImgReg2IN_337, D(0)=>ImgReg2IN_336, CLK=>nx23956, 
      RST=>RST, EN=>nx23744, Q(15)=>OutputImg2_351_EXMPLR, Q(14)=>
      OutputImg2_350_EXMPLR, Q(13)=>OutputImg2_349_EXMPLR, Q(12)=>
      OutputImg2_348_EXMPLR, Q(11)=>OutputImg2_347_EXMPLR, Q(10)=>
      OutputImg2_346_EXMPLR, Q(9)=>OutputImg2_345_EXMPLR, Q(8)=>
      OutputImg2_344_EXMPLR, Q(7)=>OutputImg2_343_EXMPLR, Q(6)=>
      OutputImg2_342_EXMPLR, Q(5)=>OutputImg2_341_EXMPLR, Q(4)=>
      OutputImg2_340_EXMPLR, Q(3)=>OutputImg2_339_EXMPLR, Q(2)=>
      OutputImg2_338_EXMPLR, Q(1)=>OutputImg2_337_EXMPLR, Q(0)=>
      OutputImg2_336_EXMPLR);
   loop3_21_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_351, D(14)=>
      ImgReg3IN_350, D(13)=>ImgReg3IN_349, D(12)=>ImgReg3IN_348, D(11)=>
      ImgReg3IN_347, D(10)=>ImgReg3IN_346, D(9)=>ImgReg3IN_345, D(8)=>
      ImgReg3IN_344, D(7)=>ImgReg3IN_343, D(6)=>ImgReg3IN_342, D(5)=>
      ImgReg3IN_341, D(4)=>ImgReg3IN_340, D(3)=>ImgReg3IN_339, D(2)=>
      ImgReg3IN_338, D(1)=>ImgReg3IN_337, D(0)=>ImgReg3IN_336, CLK=>nx23958, 
      RST=>RST, EN=>nx23754, Q(15)=>OutputImg3_351_EXMPLR, Q(14)=>
      OutputImg3_350_EXMPLR, Q(13)=>OutputImg3_349_EXMPLR, Q(12)=>
      OutputImg3_348_EXMPLR, Q(11)=>OutputImg3_347_EXMPLR, Q(10)=>
      OutputImg3_346_EXMPLR, Q(9)=>OutputImg3_345_EXMPLR, Q(8)=>
      OutputImg3_344_EXMPLR, Q(7)=>OutputImg3_343_EXMPLR, Q(6)=>
      OutputImg3_342_EXMPLR, Q(5)=>OutputImg3_341_EXMPLR, Q(4)=>
      OutputImg3_340_EXMPLR, Q(3)=>OutputImg3_339_EXMPLR, Q(2)=>
      OutputImg3_338_EXMPLR, Q(1)=>OutputImg3_337_EXMPLR, Q(0)=>
      OutputImg3_336_EXMPLR);
   loop3_21_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_351, D(14)=>
      ImgReg4IN_350, D(13)=>ImgReg4IN_349, D(12)=>ImgReg4IN_348, D(11)=>
      ImgReg4IN_347, D(10)=>ImgReg4IN_346, D(9)=>ImgReg4IN_345, D(8)=>
      ImgReg4IN_344, D(7)=>ImgReg4IN_343, D(6)=>ImgReg4IN_342, D(5)=>
      ImgReg4IN_341, D(4)=>ImgReg4IN_340, D(3)=>ImgReg4IN_339, D(2)=>
      ImgReg4IN_338, D(1)=>ImgReg4IN_337, D(0)=>ImgReg4IN_336, CLK=>nx23958, 
      RST=>RST, EN=>nx23764, Q(15)=>OutputImg4_351_EXMPLR, Q(14)=>
      OutputImg4_350_EXMPLR, Q(13)=>OutputImg4_349_EXMPLR, Q(12)=>
      OutputImg4_348_EXMPLR, Q(11)=>OutputImg4_347_EXMPLR, Q(10)=>
      OutputImg4_346_EXMPLR, Q(9)=>OutputImg4_345_EXMPLR, Q(8)=>
      OutputImg4_344_EXMPLR, Q(7)=>OutputImg4_343_EXMPLR, Q(6)=>
      OutputImg4_342_EXMPLR, Q(5)=>OutputImg4_341_EXMPLR, Q(4)=>
      OutputImg4_340_EXMPLR, Q(3)=>OutputImg4_339_EXMPLR, Q(2)=>
      OutputImg4_338_EXMPLR, Q(1)=>OutputImg4_337_EXMPLR, Q(0)=>
      OutputImg4_336_EXMPLR);
   loop3_21_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_351, D(14)=>
      ImgReg5IN_350, D(13)=>ImgReg5IN_349, D(12)=>ImgReg5IN_348, D(11)=>
      ImgReg5IN_347, D(10)=>ImgReg5IN_346, D(9)=>ImgReg5IN_345, D(8)=>
      ImgReg5IN_344, D(7)=>ImgReg5IN_343, D(6)=>ImgReg5IN_342, D(5)=>
      ImgReg5IN_341, D(4)=>ImgReg5IN_340, D(3)=>ImgReg5IN_339, D(2)=>
      ImgReg5IN_338, D(1)=>ImgReg5IN_337, D(0)=>ImgReg5IN_336, CLK=>nx23960, 
      RST=>RST, EN=>nx23774, Q(15)=>OutputImg5_351_EXMPLR, Q(14)=>
      OutputImg5_350_EXMPLR, Q(13)=>OutputImg5_349_EXMPLR, Q(12)=>
      OutputImg5_348_EXMPLR, Q(11)=>OutputImg5_347_EXMPLR, Q(10)=>
      OutputImg5_346_EXMPLR, Q(9)=>OutputImg5_345_EXMPLR, Q(8)=>
      OutputImg5_344_EXMPLR, Q(7)=>OutputImg5_343_EXMPLR, Q(6)=>
      OutputImg5_342_EXMPLR, Q(5)=>OutputImg5_341_EXMPLR, Q(4)=>
      OutputImg5_340_EXMPLR, Q(3)=>OutputImg5_339_EXMPLR, Q(2)=>
      OutputImg5_338_EXMPLR, Q(1)=>OutputImg5_337_EXMPLR, Q(0)=>
      OutputImg5_336_EXMPLR);
   loop3_22_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_383_EXMPLR, D(14)=>OutputImg0_382_EXMPLR, D(13)=>
      OutputImg0_381_EXMPLR, D(12)=>OutputImg0_380_EXMPLR, D(11)=>
      OutputImg0_379_EXMPLR, D(10)=>OutputImg0_378_EXMPLR, D(9)=>
      OutputImg0_377_EXMPLR, D(8)=>OutputImg0_376_EXMPLR, D(7)=>
      OutputImg0_375_EXMPLR, D(6)=>OutputImg0_374_EXMPLR, D(5)=>
      OutputImg0_373_EXMPLR, D(4)=>OutputImg0_372_EXMPLR, D(3)=>
      OutputImg0_371_EXMPLR, D(2)=>OutputImg0_370_EXMPLR, D(1)=>
      OutputImg0_369_EXMPLR, D(0)=>OutputImg0_368_EXMPLR, EN=>nx23702, F(15)
      =>ImgReg0IN_367, F(14)=>ImgReg0IN_366, F(13)=>ImgReg0IN_365, F(12)=>
      ImgReg0IN_364, F(11)=>ImgReg0IN_363, F(10)=>ImgReg0IN_362, F(9)=>
      ImgReg0IN_361, F(8)=>ImgReg0IN_360, F(7)=>ImgReg0IN_359, F(6)=>
      ImgReg0IN_358, F(5)=>ImgReg0IN_357, F(4)=>ImgReg0IN_356, F(3)=>
      ImgReg0IN_355, F(2)=>ImgReg0IN_354, F(1)=>ImgReg0IN_353, F(0)=>
      ImgReg0IN_352);
   loop3_22_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_383_EXMPLR, D(14)=>OutputImg1_382_EXMPLR, D(13)=>
      OutputImg1_381_EXMPLR, D(12)=>OutputImg1_380_EXMPLR, D(11)=>
      OutputImg1_379_EXMPLR, D(10)=>OutputImg1_378_EXMPLR, D(9)=>
      OutputImg1_377_EXMPLR, D(8)=>OutputImg1_376_EXMPLR, D(7)=>
      OutputImg1_375_EXMPLR, D(6)=>OutputImg1_374_EXMPLR, D(5)=>
      OutputImg1_373_EXMPLR, D(4)=>OutputImg1_372_EXMPLR, D(3)=>
      OutputImg1_371_EXMPLR, D(2)=>OutputImg1_370_EXMPLR, D(1)=>
      OutputImg1_369_EXMPLR, D(0)=>OutputImg1_368_EXMPLR, EN=>nx23704, F(15)
      =>ImgReg1IN_367, F(14)=>ImgReg1IN_366, F(13)=>ImgReg1IN_365, F(12)=>
      ImgReg1IN_364, F(11)=>ImgReg1IN_363, F(10)=>ImgReg1IN_362, F(9)=>
      ImgReg1IN_361, F(8)=>ImgReg1IN_360, F(7)=>ImgReg1IN_359, F(6)=>
      ImgReg1IN_358, F(5)=>ImgReg1IN_357, F(4)=>ImgReg1IN_356, F(3)=>
      ImgReg1IN_355, F(2)=>ImgReg1IN_354, F(1)=>ImgReg1IN_353, F(0)=>
      ImgReg1IN_352);
   loop3_22_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_383_EXMPLR, D(14)=>OutputImg2_382_EXMPLR, D(13)=>
      OutputImg2_381_EXMPLR, D(12)=>OutputImg2_380_EXMPLR, D(11)=>
      OutputImg2_379_EXMPLR, D(10)=>OutputImg2_378_EXMPLR, D(9)=>
      OutputImg2_377_EXMPLR, D(8)=>OutputImg2_376_EXMPLR, D(7)=>
      OutputImg2_375_EXMPLR, D(6)=>OutputImg2_374_EXMPLR, D(5)=>
      OutputImg2_373_EXMPLR, D(4)=>OutputImg2_372_EXMPLR, D(3)=>
      OutputImg2_371_EXMPLR, D(2)=>OutputImg2_370_EXMPLR, D(1)=>
      OutputImg2_369_EXMPLR, D(0)=>OutputImg2_368_EXMPLR, EN=>nx23704, F(15)
      =>ImgReg2IN_367, F(14)=>ImgReg2IN_366, F(13)=>ImgReg2IN_365, F(12)=>
      ImgReg2IN_364, F(11)=>ImgReg2IN_363, F(10)=>ImgReg2IN_362, F(9)=>
      ImgReg2IN_361, F(8)=>ImgReg2IN_360, F(7)=>ImgReg2IN_359, F(6)=>
      ImgReg2IN_358, F(5)=>ImgReg2IN_357, F(4)=>ImgReg2IN_356, F(3)=>
      ImgReg2IN_355, F(2)=>ImgReg2IN_354, F(1)=>ImgReg2IN_353, F(0)=>
      ImgReg2IN_352);
   loop3_22_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_383_EXMPLR, D(14)=>OutputImg3_382_EXMPLR, D(13)=>
      OutputImg3_381_EXMPLR, D(12)=>OutputImg3_380_EXMPLR, D(11)=>
      OutputImg3_379_EXMPLR, D(10)=>OutputImg3_378_EXMPLR, D(9)=>
      OutputImg3_377_EXMPLR, D(8)=>OutputImg3_376_EXMPLR, D(7)=>
      OutputImg3_375_EXMPLR, D(6)=>OutputImg3_374_EXMPLR, D(5)=>
      OutputImg3_373_EXMPLR, D(4)=>OutputImg3_372_EXMPLR, D(3)=>
      OutputImg3_371_EXMPLR, D(2)=>OutputImg3_370_EXMPLR, D(1)=>
      OutputImg3_369_EXMPLR, D(0)=>OutputImg3_368_EXMPLR, EN=>nx23704, F(15)
      =>ImgReg3IN_367, F(14)=>ImgReg3IN_366, F(13)=>ImgReg3IN_365, F(12)=>
      ImgReg3IN_364, F(11)=>ImgReg3IN_363, F(10)=>ImgReg3IN_362, F(9)=>
      ImgReg3IN_361, F(8)=>ImgReg3IN_360, F(7)=>ImgReg3IN_359, F(6)=>
      ImgReg3IN_358, F(5)=>ImgReg3IN_357, F(4)=>ImgReg3IN_356, F(3)=>
      ImgReg3IN_355, F(2)=>ImgReg3IN_354, F(1)=>ImgReg3IN_353, F(0)=>
      ImgReg3IN_352);
   loop3_22_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_383_EXMPLR, D(14)=>OutputImg4_382_EXMPLR, D(13)=>
      OutputImg4_381_EXMPLR, D(12)=>OutputImg4_380_EXMPLR, D(11)=>
      OutputImg4_379_EXMPLR, D(10)=>OutputImg4_378_EXMPLR, D(9)=>
      OutputImg4_377_EXMPLR, D(8)=>OutputImg4_376_EXMPLR, D(7)=>
      OutputImg4_375_EXMPLR, D(6)=>OutputImg4_374_EXMPLR, D(5)=>
      OutputImg4_373_EXMPLR, D(4)=>OutputImg4_372_EXMPLR, D(3)=>
      OutputImg4_371_EXMPLR, D(2)=>OutputImg4_370_EXMPLR, D(1)=>
      OutputImg4_369_EXMPLR, D(0)=>OutputImg4_368_EXMPLR, EN=>nx23704, F(15)
      =>ImgReg4IN_367, F(14)=>ImgReg4IN_366, F(13)=>ImgReg4IN_365, F(12)=>
      ImgReg4IN_364, F(11)=>ImgReg4IN_363, F(10)=>ImgReg4IN_362, F(9)=>
      ImgReg4IN_361, F(8)=>ImgReg4IN_360, F(7)=>ImgReg4IN_359, F(6)=>
      ImgReg4IN_358, F(5)=>ImgReg4IN_357, F(4)=>ImgReg4IN_356, F(3)=>
      ImgReg4IN_355, F(2)=>ImgReg4IN_354, F(1)=>ImgReg4IN_353, F(0)=>
      ImgReg4IN_352);
   loop3_22_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_383_EXMPLR, D(14)=>OutputImg5_382_EXMPLR, D(13)=>
      OutputImg5_381_EXMPLR, D(12)=>OutputImg5_380_EXMPLR, D(11)=>
      OutputImg5_379_EXMPLR, D(10)=>OutputImg5_378_EXMPLR, D(9)=>
      OutputImg5_377_EXMPLR, D(8)=>OutputImg5_376_EXMPLR, D(7)=>
      OutputImg5_375_EXMPLR, D(6)=>OutputImg5_374_EXMPLR, D(5)=>
      OutputImg5_373_EXMPLR, D(4)=>OutputImg5_372_EXMPLR, D(3)=>
      OutputImg5_371_EXMPLR, D(2)=>OutputImg5_370_EXMPLR, D(1)=>
      OutputImg5_369_EXMPLR, D(0)=>OutputImg5_368_EXMPLR, EN=>nx23704, F(15)
      =>ImgReg5IN_367, F(14)=>ImgReg5IN_366, F(13)=>ImgReg5IN_365, F(12)=>
      ImgReg5IN_364, F(11)=>ImgReg5IN_363, F(10)=>ImgReg5IN_362, F(9)=>
      ImgReg5IN_361, F(8)=>ImgReg5IN_360, F(7)=>ImgReg5IN_359, F(6)=>
      ImgReg5IN_358, F(5)=>ImgReg5IN_357, F(4)=>ImgReg5IN_356, F(3)=>
      ImgReg5IN_355, F(2)=>ImgReg5IN_354, F(1)=>ImgReg5IN_353, F(0)=>
      ImgReg5IN_352);
   loop3_22_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(367), 
      D(14)=>DATA(366), D(13)=>DATA(365), D(12)=>DATA(364), D(11)=>DATA(363), 
      D(10)=>DATA(362), D(9)=>DATA(361), D(8)=>DATA(360), D(7)=>DATA(359), 
      D(6)=>DATA(358), D(5)=>DATA(357), D(4)=>DATA(356), D(3)=>DATA(355), 
      D(2)=>DATA(354), D(1)=>DATA(353), D(0)=>DATA(352), EN=>nx23660, F(15)
      =>ImgReg0IN_367, F(14)=>ImgReg0IN_366, F(13)=>ImgReg0IN_365, F(12)=>
      ImgReg0IN_364, F(11)=>ImgReg0IN_363, F(10)=>ImgReg0IN_362, F(9)=>
      ImgReg0IN_361, F(8)=>ImgReg0IN_360, F(7)=>ImgReg0IN_359, F(6)=>
      ImgReg0IN_358, F(5)=>ImgReg0IN_357, F(4)=>ImgReg0IN_356, F(3)=>
      ImgReg0IN_355, F(2)=>ImgReg0IN_354, F(1)=>ImgReg0IN_353, F(0)=>
      ImgReg0IN_352);
   loop3_22_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(367), 
      D(14)=>DATA(366), D(13)=>DATA(365), D(12)=>DATA(364), D(11)=>DATA(363), 
      D(10)=>DATA(362), D(9)=>DATA(361), D(8)=>DATA(360), D(7)=>DATA(359), 
      D(6)=>DATA(358), D(5)=>DATA(357), D(4)=>DATA(356), D(3)=>DATA(355), 
      D(2)=>DATA(354), D(1)=>DATA(353), D(0)=>DATA(352), EN=>nx23648, F(15)
      =>ImgReg1IN_367, F(14)=>ImgReg1IN_366, F(13)=>ImgReg1IN_365, F(12)=>
      ImgReg1IN_364, F(11)=>ImgReg1IN_363, F(10)=>ImgReg1IN_362, F(9)=>
      ImgReg1IN_361, F(8)=>ImgReg1IN_360, F(7)=>ImgReg1IN_359, F(6)=>
      ImgReg1IN_358, F(5)=>ImgReg1IN_357, F(4)=>ImgReg1IN_356, F(3)=>
      ImgReg1IN_355, F(2)=>ImgReg1IN_354, F(1)=>ImgReg1IN_353, F(0)=>
      ImgReg1IN_352);
   loop3_22_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(367), 
      D(14)=>DATA(366), D(13)=>DATA(365), D(12)=>DATA(364), D(11)=>DATA(363), 
      D(10)=>DATA(362), D(9)=>DATA(361), D(8)=>DATA(360), D(7)=>DATA(359), 
      D(6)=>DATA(358), D(5)=>DATA(357), D(4)=>DATA(356), D(3)=>DATA(355), 
      D(2)=>DATA(354), D(1)=>DATA(353), D(0)=>DATA(352), EN=>nx23636, F(15)
      =>ImgReg2IN_367, F(14)=>ImgReg2IN_366, F(13)=>ImgReg2IN_365, F(12)=>
      ImgReg2IN_364, F(11)=>ImgReg2IN_363, F(10)=>ImgReg2IN_362, F(9)=>
      ImgReg2IN_361, F(8)=>ImgReg2IN_360, F(7)=>ImgReg2IN_359, F(6)=>
      ImgReg2IN_358, F(5)=>ImgReg2IN_357, F(4)=>ImgReg2IN_356, F(3)=>
      ImgReg2IN_355, F(2)=>ImgReg2IN_354, F(1)=>ImgReg2IN_353, F(0)=>
      ImgReg2IN_352);
   loop3_22_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(367), 
      D(14)=>DATA(366), D(13)=>DATA(365), D(12)=>DATA(364), D(11)=>DATA(363), 
      D(10)=>DATA(362), D(9)=>DATA(361), D(8)=>DATA(360), D(7)=>DATA(359), 
      D(6)=>DATA(358), D(5)=>DATA(357), D(4)=>DATA(356), D(3)=>DATA(355), 
      D(2)=>DATA(354), D(1)=>DATA(353), D(0)=>DATA(352), EN=>nx23624, F(15)
      =>ImgReg3IN_367, F(14)=>ImgReg3IN_366, F(13)=>ImgReg3IN_365, F(12)=>
      ImgReg3IN_364, F(11)=>ImgReg3IN_363, F(10)=>ImgReg3IN_362, F(9)=>
      ImgReg3IN_361, F(8)=>ImgReg3IN_360, F(7)=>ImgReg3IN_359, F(6)=>
      ImgReg3IN_358, F(5)=>ImgReg3IN_357, F(4)=>ImgReg3IN_356, F(3)=>
      ImgReg3IN_355, F(2)=>ImgReg3IN_354, F(1)=>ImgReg3IN_353, F(0)=>
      ImgReg3IN_352);
   loop3_22_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(367), 
      D(14)=>DATA(366), D(13)=>DATA(365), D(12)=>DATA(364), D(11)=>DATA(363), 
      D(10)=>DATA(362), D(9)=>DATA(361), D(8)=>DATA(360), D(7)=>DATA(359), 
      D(6)=>DATA(358), D(5)=>DATA(357), D(4)=>DATA(356), D(3)=>DATA(355), 
      D(2)=>DATA(354), D(1)=>DATA(353), D(0)=>DATA(352), EN=>nx23612, F(15)
      =>ImgReg4IN_367, F(14)=>ImgReg4IN_366, F(13)=>ImgReg4IN_365, F(12)=>
      ImgReg4IN_364, F(11)=>ImgReg4IN_363, F(10)=>ImgReg4IN_362, F(9)=>
      ImgReg4IN_361, F(8)=>ImgReg4IN_360, F(7)=>ImgReg4IN_359, F(6)=>
      ImgReg4IN_358, F(5)=>ImgReg4IN_357, F(4)=>ImgReg4IN_356, F(3)=>
      ImgReg4IN_355, F(2)=>ImgReg4IN_354, F(1)=>ImgReg4IN_353, F(0)=>
      ImgReg4IN_352);
   loop3_22_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(367), 
      D(14)=>DATA(366), D(13)=>DATA(365), D(12)=>DATA(364), D(11)=>DATA(363), 
      D(10)=>DATA(362), D(9)=>DATA(361), D(8)=>DATA(360), D(7)=>DATA(359), 
      D(6)=>DATA(358), D(5)=>DATA(357), D(4)=>DATA(356), D(3)=>DATA(355), 
      D(2)=>DATA(354), D(1)=>DATA(353), D(0)=>DATA(352), EN=>nx23600, F(15)
      =>ImgReg5IN_367, F(14)=>ImgReg5IN_366, F(13)=>ImgReg5IN_365, F(12)=>
      ImgReg5IN_364, F(11)=>ImgReg5IN_363, F(10)=>ImgReg5IN_362, F(9)=>
      ImgReg5IN_361, F(8)=>ImgReg5IN_360, F(7)=>ImgReg5IN_359, F(6)=>
      ImgReg5IN_358, F(5)=>ImgReg5IN_357, F(4)=>ImgReg5IN_356, F(3)=>
      ImgReg5IN_355, F(2)=>ImgReg5IN_354, F(1)=>ImgReg5IN_353, F(0)=>
      ImgReg5IN_352);
   loop3_22_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_367_EXMPLR, D(14)=>OutputImg1_366_EXMPLR, D(13)=>
      OutputImg1_365_EXMPLR, D(12)=>OutputImg1_364_EXMPLR, D(11)=>
      OutputImg1_363_EXMPLR, D(10)=>OutputImg1_362_EXMPLR, D(9)=>
      OutputImg1_361_EXMPLR, D(8)=>OutputImg1_360_EXMPLR, D(7)=>
      OutputImg1_359_EXMPLR, D(6)=>OutputImg1_358_EXMPLR, D(5)=>
      OutputImg1_357_EXMPLR, D(4)=>OutputImg1_356_EXMPLR, D(3)=>
      OutputImg1_355_EXMPLR, D(2)=>OutputImg1_354_EXMPLR, D(1)=>
      OutputImg1_353_EXMPLR, D(0)=>OutputImg1_352_EXMPLR, EN=>nx23816, F(15)
      =>ImgReg0IN_367, F(14)=>ImgReg0IN_366, F(13)=>ImgReg0IN_365, F(12)=>
      ImgReg0IN_364, F(11)=>ImgReg0IN_363, F(10)=>ImgReg0IN_362, F(9)=>
      ImgReg0IN_361, F(8)=>ImgReg0IN_360, F(7)=>ImgReg0IN_359, F(6)=>
      ImgReg0IN_358, F(5)=>ImgReg0IN_357, F(4)=>ImgReg0IN_356, F(3)=>
      ImgReg0IN_355, F(2)=>ImgReg0IN_354, F(1)=>ImgReg0IN_353, F(0)=>
      ImgReg0IN_352);
   loop3_22_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_367_EXMPLR, D(14)=>OutputImg2_366_EXMPLR, D(13)=>
      OutputImg2_365_EXMPLR, D(12)=>OutputImg2_364_EXMPLR, D(11)=>
      OutputImg2_363_EXMPLR, D(10)=>OutputImg2_362_EXMPLR, D(9)=>
      OutputImg2_361_EXMPLR, D(8)=>OutputImg2_360_EXMPLR, D(7)=>
      OutputImg2_359_EXMPLR, D(6)=>OutputImg2_358_EXMPLR, D(5)=>
      OutputImg2_357_EXMPLR, D(4)=>OutputImg2_356_EXMPLR, D(3)=>
      OutputImg2_355_EXMPLR, D(2)=>OutputImg2_354_EXMPLR, D(1)=>
      OutputImg2_353_EXMPLR, D(0)=>OutputImg2_352_EXMPLR, EN=>nx23816, F(15)
      =>ImgReg1IN_367, F(14)=>ImgReg1IN_366, F(13)=>ImgReg1IN_365, F(12)=>
      ImgReg1IN_364, F(11)=>ImgReg1IN_363, F(10)=>ImgReg1IN_362, F(9)=>
      ImgReg1IN_361, F(8)=>ImgReg1IN_360, F(7)=>ImgReg1IN_359, F(6)=>
      ImgReg1IN_358, F(5)=>ImgReg1IN_357, F(4)=>ImgReg1IN_356, F(3)=>
      ImgReg1IN_355, F(2)=>ImgReg1IN_354, F(1)=>ImgReg1IN_353, F(0)=>
      ImgReg1IN_352);
   loop3_22_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_367_EXMPLR, D(14)=>OutputImg3_366_EXMPLR, D(13)=>
      OutputImg3_365_EXMPLR, D(12)=>OutputImg3_364_EXMPLR, D(11)=>
      OutputImg3_363_EXMPLR, D(10)=>OutputImg3_362_EXMPLR, D(9)=>
      OutputImg3_361_EXMPLR, D(8)=>OutputImg3_360_EXMPLR, D(7)=>
      OutputImg3_359_EXMPLR, D(6)=>OutputImg3_358_EXMPLR, D(5)=>
      OutputImg3_357_EXMPLR, D(4)=>OutputImg3_356_EXMPLR, D(3)=>
      OutputImg3_355_EXMPLR, D(2)=>OutputImg3_354_EXMPLR, D(1)=>
      OutputImg3_353_EXMPLR, D(0)=>OutputImg3_352_EXMPLR, EN=>nx23818, F(15)
      =>ImgReg2IN_367, F(14)=>ImgReg2IN_366, F(13)=>ImgReg2IN_365, F(12)=>
      ImgReg2IN_364, F(11)=>ImgReg2IN_363, F(10)=>ImgReg2IN_362, F(9)=>
      ImgReg2IN_361, F(8)=>ImgReg2IN_360, F(7)=>ImgReg2IN_359, F(6)=>
      ImgReg2IN_358, F(5)=>ImgReg2IN_357, F(4)=>ImgReg2IN_356, F(3)=>
      ImgReg2IN_355, F(2)=>ImgReg2IN_354, F(1)=>ImgReg2IN_353, F(0)=>
      ImgReg2IN_352);
   loop3_22_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_367_EXMPLR, D(14)=>OutputImg4_366_EXMPLR, D(13)=>
      OutputImg4_365_EXMPLR, D(12)=>OutputImg4_364_EXMPLR, D(11)=>
      OutputImg4_363_EXMPLR, D(10)=>OutputImg4_362_EXMPLR, D(9)=>
      OutputImg4_361_EXMPLR, D(8)=>OutputImg4_360_EXMPLR, D(7)=>
      OutputImg4_359_EXMPLR, D(6)=>OutputImg4_358_EXMPLR, D(5)=>
      OutputImg4_357_EXMPLR, D(4)=>OutputImg4_356_EXMPLR, D(3)=>
      OutputImg4_355_EXMPLR, D(2)=>OutputImg4_354_EXMPLR, D(1)=>
      OutputImg4_353_EXMPLR, D(0)=>OutputImg4_352_EXMPLR, EN=>nx23818, F(15)
      =>ImgReg3IN_367, F(14)=>ImgReg3IN_366, F(13)=>ImgReg3IN_365, F(12)=>
      ImgReg3IN_364, F(11)=>ImgReg3IN_363, F(10)=>ImgReg3IN_362, F(9)=>
      ImgReg3IN_361, F(8)=>ImgReg3IN_360, F(7)=>ImgReg3IN_359, F(6)=>
      ImgReg3IN_358, F(5)=>ImgReg3IN_357, F(4)=>ImgReg3IN_356, F(3)=>
      ImgReg3IN_355, F(2)=>ImgReg3IN_354, F(1)=>ImgReg3IN_353, F(0)=>
      ImgReg3IN_352);
   loop3_22_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_367_EXMPLR, D(14)=>OutputImg5_366_EXMPLR, D(13)=>
      OutputImg5_365_EXMPLR, D(12)=>OutputImg5_364_EXMPLR, D(11)=>
      OutputImg5_363_EXMPLR, D(10)=>OutputImg5_362_EXMPLR, D(9)=>
      OutputImg5_361_EXMPLR, D(8)=>OutputImg5_360_EXMPLR, D(7)=>
      OutputImg5_359_EXMPLR, D(6)=>OutputImg5_358_EXMPLR, D(5)=>
      OutputImg5_357_EXMPLR, D(4)=>OutputImg5_356_EXMPLR, D(3)=>
      OutputImg5_355_EXMPLR, D(2)=>OutputImg5_354_EXMPLR, D(1)=>
      OutputImg5_353_EXMPLR, D(0)=>OutputImg5_352_EXMPLR, EN=>nx23818, F(15)
      =>ImgReg4IN_367, F(14)=>ImgReg4IN_366, F(13)=>ImgReg4IN_365, F(12)=>
      ImgReg4IN_364, F(11)=>ImgReg4IN_363, F(10)=>ImgReg4IN_362, F(9)=>
      ImgReg4IN_361, F(8)=>ImgReg4IN_360, F(7)=>ImgReg4IN_359, F(6)=>
      ImgReg4IN_358, F(5)=>ImgReg4IN_357, F(4)=>ImgReg4IN_356, F(3)=>
      ImgReg4IN_355, F(2)=>ImgReg4IN_354, F(1)=>ImgReg4IN_353, F(0)=>
      ImgReg4IN_352);
   loop3_22_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_367, D(14)=>
      ImgReg0IN_366, D(13)=>ImgReg0IN_365, D(12)=>ImgReg0IN_364, D(11)=>
      ImgReg0IN_363, D(10)=>ImgReg0IN_362, D(9)=>ImgReg0IN_361, D(8)=>
      ImgReg0IN_360, D(7)=>ImgReg0IN_359, D(6)=>ImgReg0IN_358, D(5)=>
      ImgReg0IN_357, D(4)=>ImgReg0IN_356, D(3)=>ImgReg0IN_355, D(2)=>
      ImgReg0IN_354, D(1)=>ImgReg0IN_353, D(0)=>ImgReg0IN_352, CLK=>nx23960, 
      RST=>RST, EN=>nx23724, Q(15)=>OutputImg0_367_EXMPLR, Q(14)=>
      OutputImg0_366_EXMPLR, Q(13)=>OutputImg0_365_EXMPLR, Q(12)=>
      OutputImg0_364_EXMPLR, Q(11)=>OutputImg0_363_EXMPLR, Q(10)=>
      OutputImg0_362_EXMPLR, Q(9)=>OutputImg0_361_EXMPLR, Q(8)=>
      OutputImg0_360_EXMPLR, Q(7)=>OutputImg0_359_EXMPLR, Q(6)=>
      OutputImg0_358_EXMPLR, Q(5)=>OutputImg0_357_EXMPLR, Q(4)=>
      OutputImg0_356_EXMPLR, Q(3)=>OutputImg0_355_EXMPLR, Q(2)=>
      OutputImg0_354_EXMPLR, Q(1)=>OutputImg0_353_EXMPLR, Q(0)=>
      OutputImg0_352_EXMPLR);
   loop3_22_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_367, D(14)=>
      ImgReg1IN_366, D(13)=>ImgReg1IN_365, D(12)=>ImgReg1IN_364, D(11)=>
      ImgReg1IN_363, D(10)=>ImgReg1IN_362, D(9)=>ImgReg1IN_361, D(8)=>
      ImgReg1IN_360, D(7)=>ImgReg1IN_359, D(6)=>ImgReg1IN_358, D(5)=>
      ImgReg1IN_357, D(4)=>ImgReg1IN_356, D(3)=>ImgReg1IN_355, D(2)=>
      ImgReg1IN_354, D(1)=>ImgReg1IN_353, D(0)=>ImgReg1IN_352, CLK=>nx23962, 
      RST=>RST, EN=>nx23734, Q(15)=>OutputImg1_367_EXMPLR, Q(14)=>
      OutputImg1_366_EXMPLR, Q(13)=>OutputImg1_365_EXMPLR, Q(12)=>
      OutputImg1_364_EXMPLR, Q(11)=>OutputImg1_363_EXMPLR, Q(10)=>
      OutputImg1_362_EXMPLR, Q(9)=>OutputImg1_361_EXMPLR, Q(8)=>
      OutputImg1_360_EXMPLR, Q(7)=>OutputImg1_359_EXMPLR, Q(6)=>
      OutputImg1_358_EXMPLR, Q(5)=>OutputImg1_357_EXMPLR, Q(4)=>
      OutputImg1_356_EXMPLR, Q(3)=>OutputImg1_355_EXMPLR, Q(2)=>
      OutputImg1_354_EXMPLR, Q(1)=>OutputImg1_353_EXMPLR, Q(0)=>
      OutputImg1_352_EXMPLR);
   loop3_22_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_367, D(14)=>
      ImgReg2IN_366, D(13)=>ImgReg2IN_365, D(12)=>ImgReg2IN_364, D(11)=>
      ImgReg2IN_363, D(10)=>ImgReg2IN_362, D(9)=>ImgReg2IN_361, D(8)=>
      ImgReg2IN_360, D(7)=>ImgReg2IN_359, D(6)=>ImgReg2IN_358, D(5)=>
      ImgReg2IN_357, D(4)=>ImgReg2IN_356, D(3)=>ImgReg2IN_355, D(2)=>
      ImgReg2IN_354, D(1)=>ImgReg2IN_353, D(0)=>ImgReg2IN_352, CLK=>nx23962, 
      RST=>RST, EN=>nx23744, Q(15)=>OutputImg2_367_EXMPLR, Q(14)=>
      OutputImg2_366_EXMPLR, Q(13)=>OutputImg2_365_EXMPLR, Q(12)=>
      OutputImg2_364_EXMPLR, Q(11)=>OutputImg2_363_EXMPLR, Q(10)=>
      OutputImg2_362_EXMPLR, Q(9)=>OutputImg2_361_EXMPLR, Q(8)=>
      OutputImg2_360_EXMPLR, Q(7)=>OutputImg2_359_EXMPLR, Q(6)=>
      OutputImg2_358_EXMPLR, Q(5)=>OutputImg2_357_EXMPLR, Q(4)=>
      OutputImg2_356_EXMPLR, Q(3)=>OutputImg2_355_EXMPLR, Q(2)=>
      OutputImg2_354_EXMPLR, Q(1)=>OutputImg2_353_EXMPLR, Q(0)=>
      OutputImg2_352_EXMPLR);
   loop3_22_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_367, D(14)=>
      ImgReg3IN_366, D(13)=>ImgReg3IN_365, D(12)=>ImgReg3IN_364, D(11)=>
      ImgReg3IN_363, D(10)=>ImgReg3IN_362, D(9)=>ImgReg3IN_361, D(8)=>
      ImgReg3IN_360, D(7)=>ImgReg3IN_359, D(6)=>ImgReg3IN_358, D(5)=>
      ImgReg3IN_357, D(4)=>ImgReg3IN_356, D(3)=>ImgReg3IN_355, D(2)=>
      ImgReg3IN_354, D(1)=>ImgReg3IN_353, D(0)=>ImgReg3IN_352, CLK=>nx23964, 
      RST=>RST, EN=>nx23754, Q(15)=>OutputImg3_367_EXMPLR, Q(14)=>
      OutputImg3_366_EXMPLR, Q(13)=>OutputImg3_365_EXMPLR, Q(12)=>
      OutputImg3_364_EXMPLR, Q(11)=>OutputImg3_363_EXMPLR, Q(10)=>
      OutputImg3_362_EXMPLR, Q(9)=>OutputImg3_361_EXMPLR, Q(8)=>
      OutputImg3_360_EXMPLR, Q(7)=>OutputImg3_359_EXMPLR, Q(6)=>
      OutputImg3_358_EXMPLR, Q(5)=>OutputImg3_357_EXMPLR, Q(4)=>
      OutputImg3_356_EXMPLR, Q(3)=>OutputImg3_355_EXMPLR, Q(2)=>
      OutputImg3_354_EXMPLR, Q(1)=>OutputImg3_353_EXMPLR, Q(0)=>
      OutputImg3_352_EXMPLR);
   loop3_22_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_367, D(14)=>
      ImgReg4IN_366, D(13)=>ImgReg4IN_365, D(12)=>ImgReg4IN_364, D(11)=>
      ImgReg4IN_363, D(10)=>ImgReg4IN_362, D(9)=>ImgReg4IN_361, D(8)=>
      ImgReg4IN_360, D(7)=>ImgReg4IN_359, D(6)=>ImgReg4IN_358, D(5)=>
      ImgReg4IN_357, D(4)=>ImgReg4IN_356, D(3)=>ImgReg4IN_355, D(2)=>
      ImgReg4IN_354, D(1)=>ImgReg4IN_353, D(0)=>ImgReg4IN_352, CLK=>nx23964, 
      RST=>RST, EN=>nx23764, Q(15)=>OutputImg4_367_EXMPLR, Q(14)=>
      OutputImg4_366_EXMPLR, Q(13)=>OutputImg4_365_EXMPLR, Q(12)=>
      OutputImg4_364_EXMPLR, Q(11)=>OutputImg4_363_EXMPLR, Q(10)=>
      OutputImg4_362_EXMPLR, Q(9)=>OutputImg4_361_EXMPLR, Q(8)=>
      OutputImg4_360_EXMPLR, Q(7)=>OutputImg4_359_EXMPLR, Q(6)=>
      OutputImg4_358_EXMPLR, Q(5)=>OutputImg4_357_EXMPLR, Q(4)=>
      OutputImg4_356_EXMPLR, Q(3)=>OutputImg4_355_EXMPLR, Q(2)=>
      OutputImg4_354_EXMPLR, Q(1)=>OutputImg4_353_EXMPLR, Q(0)=>
      OutputImg4_352_EXMPLR);
   loop3_22_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_367, D(14)=>
      ImgReg5IN_366, D(13)=>ImgReg5IN_365, D(12)=>ImgReg5IN_364, D(11)=>
      ImgReg5IN_363, D(10)=>ImgReg5IN_362, D(9)=>ImgReg5IN_361, D(8)=>
      ImgReg5IN_360, D(7)=>ImgReg5IN_359, D(6)=>ImgReg5IN_358, D(5)=>
      ImgReg5IN_357, D(4)=>ImgReg5IN_356, D(3)=>ImgReg5IN_355, D(2)=>
      ImgReg5IN_354, D(1)=>ImgReg5IN_353, D(0)=>ImgReg5IN_352, CLK=>nx23966, 
      RST=>RST, EN=>nx23774, Q(15)=>OutputImg5_367_EXMPLR, Q(14)=>
      OutputImg5_366_EXMPLR, Q(13)=>OutputImg5_365_EXMPLR, Q(12)=>
      OutputImg5_364_EXMPLR, Q(11)=>OutputImg5_363_EXMPLR, Q(10)=>
      OutputImg5_362_EXMPLR, Q(9)=>OutputImg5_361_EXMPLR, Q(8)=>
      OutputImg5_360_EXMPLR, Q(7)=>OutputImg5_359_EXMPLR, Q(6)=>
      OutputImg5_358_EXMPLR, Q(5)=>OutputImg5_357_EXMPLR, Q(4)=>
      OutputImg5_356_EXMPLR, Q(3)=>OutputImg5_355_EXMPLR, Q(2)=>
      OutputImg5_354_EXMPLR, Q(1)=>OutputImg5_353_EXMPLR, Q(0)=>
      OutputImg5_352_EXMPLR);
   loop3_23_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_399_EXMPLR, D(14)=>OutputImg0_398_EXMPLR, D(13)=>
      OutputImg0_397_EXMPLR, D(12)=>OutputImg0_396_EXMPLR, D(11)=>
      OutputImg0_395_EXMPLR, D(10)=>OutputImg0_394_EXMPLR, D(9)=>
      OutputImg0_393_EXMPLR, D(8)=>OutputImg0_392_EXMPLR, D(7)=>
      OutputImg0_391_EXMPLR, D(6)=>OutputImg0_390_EXMPLR, D(5)=>
      OutputImg0_389_EXMPLR, D(4)=>OutputImg0_388_EXMPLR, D(3)=>
      OutputImg0_387_EXMPLR, D(2)=>OutputImg0_386_EXMPLR, D(1)=>
      OutputImg0_385_EXMPLR, D(0)=>OutputImg0_384_EXMPLR, EN=>nx23704, F(15)
      =>ImgReg0IN_383, F(14)=>ImgReg0IN_382, F(13)=>ImgReg0IN_381, F(12)=>
      ImgReg0IN_380, F(11)=>ImgReg0IN_379, F(10)=>ImgReg0IN_378, F(9)=>
      ImgReg0IN_377, F(8)=>ImgReg0IN_376, F(7)=>ImgReg0IN_375, F(6)=>
      ImgReg0IN_374, F(5)=>ImgReg0IN_373, F(4)=>ImgReg0IN_372, F(3)=>
      ImgReg0IN_371, F(2)=>ImgReg0IN_370, F(1)=>ImgReg0IN_369, F(0)=>
      ImgReg0IN_368);
   loop3_23_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_399_EXMPLR, D(14)=>OutputImg1_398_EXMPLR, D(13)=>
      OutputImg1_397_EXMPLR, D(12)=>OutputImg1_396_EXMPLR, D(11)=>
      OutputImg1_395_EXMPLR, D(10)=>OutputImg1_394_EXMPLR, D(9)=>
      OutputImg1_393_EXMPLR, D(8)=>OutputImg1_392_EXMPLR, D(7)=>
      OutputImg1_391_EXMPLR, D(6)=>OutputImg1_390_EXMPLR, D(5)=>
      OutputImg1_389_EXMPLR, D(4)=>OutputImg1_388_EXMPLR, D(3)=>
      OutputImg1_387_EXMPLR, D(2)=>OutputImg1_386_EXMPLR, D(1)=>
      OutputImg1_385_EXMPLR, D(0)=>OutputImg1_384_EXMPLR, EN=>nx23704, F(15)
      =>ImgReg1IN_383, F(14)=>ImgReg1IN_382, F(13)=>ImgReg1IN_381, F(12)=>
      ImgReg1IN_380, F(11)=>ImgReg1IN_379, F(10)=>ImgReg1IN_378, F(9)=>
      ImgReg1IN_377, F(8)=>ImgReg1IN_376, F(7)=>ImgReg1IN_375, F(6)=>
      ImgReg1IN_374, F(5)=>ImgReg1IN_373, F(4)=>ImgReg1IN_372, F(3)=>
      ImgReg1IN_371, F(2)=>ImgReg1IN_370, F(1)=>ImgReg1IN_369, F(0)=>
      ImgReg1IN_368);
   loop3_23_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_399_EXMPLR, D(14)=>OutputImg2_398_EXMPLR, D(13)=>
      OutputImg2_397_EXMPLR, D(12)=>OutputImg2_396_EXMPLR, D(11)=>
      OutputImg2_395_EXMPLR, D(10)=>OutputImg2_394_EXMPLR, D(9)=>
      OutputImg2_393_EXMPLR, D(8)=>OutputImg2_392_EXMPLR, D(7)=>
      OutputImg2_391_EXMPLR, D(6)=>OutputImg2_390_EXMPLR, D(5)=>
      OutputImg2_389_EXMPLR, D(4)=>OutputImg2_388_EXMPLR, D(3)=>
      OutputImg2_387_EXMPLR, D(2)=>OutputImg2_386_EXMPLR, D(1)=>
      OutputImg2_385_EXMPLR, D(0)=>OutputImg2_384_EXMPLR, EN=>nx23706, F(15)
      =>ImgReg2IN_383, F(14)=>ImgReg2IN_382, F(13)=>ImgReg2IN_381, F(12)=>
      ImgReg2IN_380, F(11)=>ImgReg2IN_379, F(10)=>ImgReg2IN_378, F(9)=>
      ImgReg2IN_377, F(8)=>ImgReg2IN_376, F(7)=>ImgReg2IN_375, F(6)=>
      ImgReg2IN_374, F(5)=>ImgReg2IN_373, F(4)=>ImgReg2IN_372, F(3)=>
      ImgReg2IN_371, F(2)=>ImgReg2IN_370, F(1)=>ImgReg2IN_369, F(0)=>
      ImgReg2IN_368);
   loop3_23_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_399_EXMPLR, D(14)=>OutputImg3_398_EXMPLR, D(13)=>
      OutputImg3_397_EXMPLR, D(12)=>OutputImg3_396_EXMPLR, D(11)=>
      OutputImg3_395_EXMPLR, D(10)=>OutputImg3_394_EXMPLR, D(9)=>
      OutputImg3_393_EXMPLR, D(8)=>OutputImg3_392_EXMPLR, D(7)=>
      OutputImg3_391_EXMPLR, D(6)=>OutputImg3_390_EXMPLR, D(5)=>
      OutputImg3_389_EXMPLR, D(4)=>OutputImg3_388_EXMPLR, D(3)=>
      OutputImg3_387_EXMPLR, D(2)=>OutputImg3_386_EXMPLR, D(1)=>
      OutputImg3_385_EXMPLR, D(0)=>OutputImg3_384_EXMPLR, EN=>nx23706, F(15)
      =>ImgReg3IN_383, F(14)=>ImgReg3IN_382, F(13)=>ImgReg3IN_381, F(12)=>
      ImgReg3IN_380, F(11)=>ImgReg3IN_379, F(10)=>ImgReg3IN_378, F(9)=>
      ImgReg3IN_377, F(8)=>ImgReg3IN_376, F(7)=>ImgReg3IN_375, F(6)=>
      ImgReg3IN_374, F(5)=>ImgReg3IN_373, F(4)=>ImgReg3IN_372, F(3)=>
      ImgReg3IN_371, F(2)=>ImgReg3IN_370, F(1)=>ImgReg3IN_369, F(0)=>
      ImgReg3IN_368);
   loop3_23_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_399_EXMPLR, D(14)=>OutputImg4_398_EXMPLR, D(13)=>
      OutputImg4_397_EXMPLR, D(12)=>OutputImg4_396_EXMPLR, D(11)=>
      OutputImg4_395_EXMPLR, D(10)=>OutputImg4_394_EXMPLR, D(9)=>
      OutputImg4_393_EXMPLR, D(8)=>OutputImg4_392_EXMPLR, D(7)=>
      OutputImg4_391_EXMPLR, D(6)=>OutputImg4_390_EXMPLR, D(5)=>
      OutputImg4_389_EXMPLR, D(4)=>OutputImg4_388_EXMPLR, D(3)=>
      OutputImg4_387_EXMPLR, D(2)=>OutputImg4_386_EXMPLR, D(1)=>
      OutputImg4_385_EXMPLR, D(0)=>OutputImg4_384_EXMPLR, EN=>nx23706, F(15)
      =>ImgReg4IN_383, F(14)=>ImgReg4IN_382, F(13)=>ImgReg4IN_381, F(12)=>
      ImgReg4IN_380, F(11)=>ImgReg4IN_379, F(10)=>ImgReg4IN_378, F(9)=>
      ImgReg4IN_377, F(8)=>ImgReg4IN_376, F(7)=>ImgReg4IN_375, F(6)=>
      ImgReg4IN_374, F(5)=>ImgReg4IN_373, F(4)=>ImgReg4IN_372, F(3)=>
      ImgReg4IN_371, F(2)=>ImgReg4IN_370, F(1)=>ImgReg4IN_369, F(0)=>
      ImgReg4IN_368);
   loop3_23_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_399_EXMPLR, D(14)=>OutputImg5_398_EXMPLR, D(13)=>
      OutputImg5_397_EXMPLR, D(12)=>OutputImg5_396_EXMPLR, D(11)=>
      OutputImg5_395_EXMPLR, D(10)=>OutputImg5_394_EXMPLR, D(9)=>
      OutputImg5_393_EXMPLR, D(8)=>OutputImg5_392_EXMPLR, D(7)=>
      OutputImg5_391_EXMPLR, D(6)=>OutputImg5_390_EXMPLR, D(5)=>
      OutputImg5_389_EXMPLR, D(4)=>OutputImg5_388_EXMPLR, D(3)=>
      OutputImg5_387_EXMPLR, D(2)=>OutputImg5_386_EXMPLR, D(1)=>
      OutputImg5_385_EXMPLR, D(0)=>OutputImg5_384_EXMPLR, EN=>nx23706, F(15)
      =>ImgReg5IN_383, F(14)=>ImgReg5IN_382, F(13)=>ImgReg5IN_381, F(12)=>
      ImgReg5IN_380, F(11)=>ImgReg5IN_379, F(10)=>ImgReg5IN_378, F(9)=>
      ImgReg5IN_377, F(8)=>ImgReg5IN_376, F(7)=>ImgReg5IN_375, F(6)=>
      ImgReg5IN_374, F(5)=>ImgReg5IN_373, F(4)=>ImgReg5IN_372, F(3)=>
      ImgReg5IN_371, F(2)=>ImgReg5IN_370, F(1)=>ImgReg5IN_369, F(0)=>
      ImgReg5IN_368);
   loop3_23_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(383), 
      D(14)=>DATA(382), D(13)=>DATA(381), D(12)=>DATA(380), D(11)=>DATA(379), 
      D(10)=>DATA(378), D(9)=>DATA(377), D(8)=>DATA(376), D(7)=>DATA(375), 
      D(6)=>DATA(374), D(5)=>DATA(373), D(4)=>DATA(372), D(3)=>DATA(371), 
      D(2)=>DATA(370), D(1)=>DATA(369), D(0)=>DATA(368), EN=>nx23660, F(15)
      =>ImgReg0IN_383, F(14)=>ImgReg0IN_382, F(13)=>ImgReg0IN_381, F(12)=>
      ImgReg0IN_380, F(11)=>ImgReg0IN_379, F(10)=>ImgReg0IN_378, F(9)=>
      ImgReg0IN_377, F(8)=>ImgReg0IN_376, F(7)=>ImgReg0IN_375, F(6)=>
      ImgReg0IN_374, F(5)=>ImgReg0IN_373, F(4)=>ImgReg0IN_372, F(3)=>
      ImgReg0IN_371, F(2)=>ImgReg0IN_370, F(1)=>ImgReg0IN_369, F(0)=>
      ImgReg0IN_368);
   loop3_23_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(383), 
      D(14)=>DATA(382), D(13)=>DATA(381), D(12)=>DATA(380), D(11)=>DATA(379), 
      D(10)=>DATA(378), D(9)=>DATA(377), D(8)=>DATA(376), D(7)=>DATA(375), 
      D(6)=>DATA(374), D(5)=>DATA(373), D(4)=>DATA(372), D(3)=>DATA(371), 
      D(2)=>DATA(370), D(1)=>DATA(369), D(0)=>DATA(368), EN=>nx23648, F(15)
      =>ImgReg1IN_383, F(14)=>ImgReg1IN_382, F(13)=>ImgReg1IN_381, F(12)=>
      ImgReg1IN_380, F(11)=>ImgReg1IN_379, F(10)=>ImgReg1IN_378, F(9)=>
      ImgReg1IN_377, F(8)=>ImgReg1IN_376, F(7)=>ImgReg1IN_375, F(6)=>
      ImgReg1IN_374, F(5)=>ImgReg1IN_373, F(4)=>ImgReg1IN_372, F(3)=>
      ImgReg1IN_371, F(2)=>ImgReg1IN_370, F(1)=>ImgReg1IN_369, F(0)=>
      ImgReg1IN_368);
   loop3_23_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(383), 
      D(14)=>DATA(382), D(13)=>DATA(381), D(12)=>DATA(380), D(11)=>DATA(379), 
      D(10)=>DATA(378), D(9)=>DATA(377), D(8)=>DATA(376), D(7)=>DATA(375), 
      D(6)=>DATA(374), D(5)=>DATA(373), D(4)=>DATA(372), D(3)=>DATA(371), 
      D(2)=>DATA(370), D(1)=>DATA(369), D(0)=>DATA(368), EN=>nx23636, F(15)
      =>ImgReg2IN_383, F(14)=>ImgReg2IN_382, F(13)=>ImgReg2IN_381, F(12)=>
      ImgReg2IN_380, F(11)=>ImgReg2IN_379, F(10)=>ImgReg2IN_378, F(9)=>
      ImgReg2IN_377, F(8)=>ImgReg2IN_376, F(7)=>ImgReg2IN_375, F(6)=>
      ImgReg2IN_374, F(5)=>ImgReg2IN_373, F(4)=>ImgReg2IN_372, F(3)=>
      ImgReg2IN_371, F(2)=>ImgReg2IN_370, F(1)=>ImgReg2IN_369, F(0)=>
      ImgReg2IN_368);
   loop3_23_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(383), 
      D(14)=>DATA(382), D(13)=>DATA(381), D(12)=>DATA(380), D(11)=>DATA(379), 
      D(10)=>DATA(378), D(9)=>DATA(377), D(8)=>DATA(376), D(7)=>DATA(375), 
      D(6)=>DATA(374), D(5)=>DATA(373), D(4)=>DATA(372), D(3)=>DATA(371), 
      D(2)=>DATA(370), D(1)=>DATA(369), D(0)=>DATA(368), EN=>nx23624, F(15)
      =>ImgReg3IN_383, F(14)=>ImgReg3IN_382, F(13)=>ImgReg3IN_381, F(12)=>
      ImgReg3IN_380, F(11)=>ImgReg3IN_379, F(10)=>ImgReg3IN_378, F(9)=>
      ImgReg3IN_377, F(8)=>ImgReg3IN_376, F(7)=>ImgReg3IN_375, F(6)=>
      ImgReg3IN_374, F(5)=>ImgReg3IN_373, F(4)=>ImgReg3IN_372, F(3)=>
      ImgReg3IN_371, F(2)=>ImgReg3IN_370, F(1)=>ImgReg3IN_369, F(0)=>
      ImgReg3IN_368);
   loop3_23_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(383), 
      D(14)=>DATA(382), D(13)=>DATA(381), D(12)=>DATA(380), D(11)=>DATA(379), 
      D(10)=>DATA(378), D(9)=>DATA(377), D(8)=>DATA(376), D(7)=>DATA(375), 
      D(6)=>DATA(374), D(5)=>DATA(373), D(4)=>DATA(372), D(3)=>DATA(371), 
      D(2)=>DATA(370), D(1)=>DATA(369), D(0)=>DATA(368), EN=>nx23612, F(15)
      =>ImgReg4IN_383, F(14)=>ImgReg4IN_382, F(13)=>ImgReg4IN_381, F(12)=>
      ImgReg4IN_380, F(11)=>ImgReg4IN_379, F(10)=>ImgReg4IN_378, F(9)=>
      ImgReg4IN_377, F(8)=>ImgReg4IN_376, F(7)=>ImgReg4IN_375, F(6)=>
      ImgReg4IN_374, F(5)=>ImgReg4IN_373, F(4)=>ImgReg4IN_372, F(3)=>
      ImgReg4IN_371, F(2)=>ImgReg4IN_370, F(1)=>ImgReg4IN_369, F(0)=>
      ImgReg4IN_368);
   loop3_23_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(383), 
      D(14)=>DATA(382), D(13)=>DATA(381), D(12)=>DATA(380), D(11)=>DATA(379), 
      D(10)=>DATA(378), D(9)=>DATA(377), D(8)=>DATA(376), D(7)=>DATA(375), 
      D(6)=>DATA(374), D(5)=>DATA(373), D(4)=>DATA(372), D(3)=>DATA(371), 
      D(2)=>DATA(370), D(1)=>DATA(369), D(0)=>DATA(368), EN=>nx23600, F(15)
      =>ImgReg5IN_383, F(14)=>ImgReg5IN_382, F(13)=>ImgReg5IN_381, F(12)=>
      ImgReg5IN_380, F(11)=>ImgReg5IN_379, F(10)=>ImgReg5IN_378, F(9)=>
      ImgReg5IN_377, F(8)=>ImgReg5IN_376, F(7)=>ImgReg5IN_375, F(6)=>
      ImgReg5IN_374, F(5)=>ImgReg5IN_373, F(4)=>ImgReg5IN_372, F(3)=>
      ImgReg5IN_371, F(2)=>ImgReg5IN_370, F(1)=>ImgReg5IN_369, F(0)=>
      ImgReg5IN_368);
   loop3_23_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_383_EXMPLR, D(14)=>OutputImg1_382_EXMPLR, D(13)=>
      OutputImg1_381_EXMPLR, D(12)=>OutputImg1_380_EXMPLR, D(11)=>
      OutputImg1_379_EXMPLR, D(10)=>OutputImg1_378_EXMPLR, D(9)=>
      OutputImg1_377_EXMPLR, D(8)=>OutputImg1_376_EXMPLR, D(7)=>
      OutputImg1_375_EXMPLR, D(6)=>OutputImg1_374_EXMPLR, D(5)=>
      OutputImg1_373_EXMPLR, D(4)=>OutputImg1_372_EXMPLR, D(3)=>
      OutputImg1_371_EXMPLR, D(2)=>OutputImg1_370_EXMPLR, D(1)=>
      OutputImg1_369_EXMPLR, D(0)=>OutputImg1_368_EXMPLR, EN=>nx23818, F(15)
      =>ImgReg0IN_383, F(14)=>ImgReg0IN_382, F(13)=>ImgReg0IN_381, F(12)=>
      ImgReg0IN_380, F(11)=>ImgReg0IN_379, F(10)=>ImgReg0IN_378, F(9)=>
      ImgReg0IN_377, F(8)=>ImgReg0IN_376, F(7)=>ImgReg0IN_375, F(6)=>
      ImgReg0IN_374, F(5)=>ImgReg0IN_373, F(4)=>ImgReg0IN_372, F(3)=>
      ImgReg0IN_371, F(2)=>ImgReg0IN_370, F(1)=>ImgReg0IN_369, F(0)=>
      ImgReg0IN_368);
   loop3_23_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_383_EXMPLR, D(14)=>OutputImg2_382_EXMPLR, D(13)=>
      OutputImg2_381_EXMPLR, D(12)=>OutputImg2_380_EXMPLR, D(11)=>
      OutputImg2_379_EXMPLR, D(10)=>OutputImg2_378_EXMPLR, D(9)=>
      OutputImg2_377_EXMPLR, D(8)=>OutputImg2_376_EXMPLR, D(7)=>
      OutputImg2_375_EXMPLR, D(6)=>OutputImg2_374_EXMPLR, D(5)=>
      OutputImg2_373_EXMPLR, D(4)=>OutputImg2_372_EXMPLR, D(3)=>
      OutputImg2_371_EXMPLR, D(2)=>OutputImg2_370_EXMPLR, D(1)=>
      OutputImg2_369_EXMPLR, D(0)=>OutputImg2_368_EXMPLR, EN=>nx23818, F(15)
      =>ImgReg1IN_383, F(14)=>ImgReg1IN_382, F(13)=>ImgReg1IN_381, F(12)=>
      ImgReg1IN_380, F(11)=>ImgReg1IN_379, F(10)=>ImgReg1IN_378, F(9)=>
      ImgReg1IN_377, F(8)=>ImgReg1IN_376, F(7)=>ImgReg1IN_375, F(6)=>
      ImgReg1IN_374, F(5)=>ImgReg1IN_373, F(4)=>ImgReg1IN_372, F(3)=>
      ImgReg1IN_371, F(2)=>ImgReg1IN_370, F(1)=>ImgReg1IN_369, F(0)=>
      ImgReg1IN_368);
   loop3_23_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_383_EXMPLR, D(14)=>OutputImg3_382_EXMPLR, D(13)=>
      OutputImg3_381_EXMPLR, D(12)=>OutputImg3_380_EXMPLR, D(11)=>
      OutputImg3_379_EXMPLR, D(10)=>OutputImg3_378_EXMPLR, D(9)=>
      OutputImg3_377_EXMPLR, D(8)=>OutputImg3_376_EXMPLR, D(7)=>
      OutputImg3_375_EXMPLR, D(6)=>OutputImg3_374_EXMPLR, D(5)=>
      OutputImg3_373_EXMPLR, D(4)=>OutputImg3_372_EXMPLR, D(3)=>
      OutputImg3_371_EXMPLR, D(2)=>OutputImg3_370_EXMPLR, D(1)=>
      OutputImg3_369_EXMPLR, D(0)=>OutputImg3_368_EXMPLR, EN=>nx23818, F(15)
      =>ImgReg2IN_383, F(14)=>ImgReg2IN_382, F(13)=>ImgReg2IN_381, F(12)=>
      ImgReg2IN_380, F(11)=>ImgReg2IN_379, F(10)=>ImgReg2IN_378, F(9)=>
      ImgReg2IN_377, F(8)=>ImgReg2IN_376, F(7)=>ImgReg2IN_375, F(6)=>
      ImgReg2IN_374, F(5)=>ImgReg2IN_373, F(4)=>ImgReg2IN_372, F(3)=>
      ImgReg2IN_371, F(2)=>ImgReg2IN_370, F(1)=>ImgReg2IN_369, F(0)=>
      ImgReg2IN_368);
   loop3_23_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_383_EXMPLR, D(14)=>OutputImg4_382_EXMPLR, D(13)=>
      OutputImg4_381_EXMPLR, D(12)=>OutputImg4_380_EXMPLR, D(11)=>
      OutputImg4_379_EXMPLR, D(10)=>OutputImg4_378_EXMPLR, D(9)=>
      OutputImg4_377_EXMPLR, D(8)=>OutputImg4_376_EXMPLR, D(7)=>
      OutputImg4_375_EXMPLR, D(6)=>OutputImg4_374_EXMPLR, D(5)=>
      OutputImg4_373_EXMPLR, D(4)=>OutputImg4_372_EXMPLR, D(3)=>
      OutputImg4_371_EXMPLR, D(2)=>OutputImg4_370_EXMPLR, D(1)=>
      OutputImg4_369_EXMPLR, D(0)=>OutputImg4_368_EXMPLR, EN=>nx23818, F(15)
      =>ImgReg3IN_383, F(14)=>ImgReg3IN_382, F(13)=>ImgReg3IN_381, F(12)=>
      ImgReg3IN_380, F(11)=>ImgReg3IN_379, F(10)=>ImgReg3IN_378, F(9)=>
      ImgReg3IN_377, F(8)=>ImgReg3IN_376, F(7)=>ImgReg3IN_375, F(6)=>
      ImgReg3IN_374, F(5)=>ImgReg3IN_373, F(4)=>ImgReg3IN_372, F(3)=>
      ImgReg3IN_371, F(2)=>ImgReg3IN_370, F(1)=>ImgReg3IN_369, F(0)=>
      ImgReg3IN_368);
   loop3_23_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_383_EXMPLR, D(14)=>OutputImg5_382_EXMPLR, D(13)=>
      OutputImg5_381_EXMPLR, D(12)=>OutputImg5_380_EXMPLR, D(11)=>
      OutputImg5_379_EXMPLR, D(10)=>OutputImg5_378_EXMPLR, D(9)=>
      OutputImg5_377_EXMPLR, D(8)=>OutputImg5_376_EXMPLR, D(7)=>
      OutputImg5_375_EXMPLR, D(6)=>OutputImg5_374_EXMPLR, D(5)=>
      OutputImg5_373_EXMPLR, D(4)=>OutputImg5_372_EXMPLR, D(3)=>
      OutputImg5_371_EXMPLR, D(2)=>OutputImg5_370_EXMPLR, D(1)=>
      OutputImg5_369_EXMPLR, D(0)=>OutputImg5_368_EXMPLR, EN=>nx23820, F(15)
      =>ImgReg4IN_383, F(14)=>ImgReg4IN_382, F(13)=>ImgReg4IN_381, F(12)=>
      ImgReg4IN_380, F(11)=>ImgReg4IN_379, F(10)=>ImgReg4IN_378, F(9)=>
      ImgReg4IN_377, F(8)=>ImgReg4IN_376, F(7)=>ImgReg4IN_375, F(6)=>
      ImgReg4IN_374, F(5)=>ImgReg4IN_373, F(4)=>ImgReg4IN_372, F(3)=>
      ImgReg4IN_371, F(2)=>ImgReg4IN_370, F(1)=>ImgReg4IN_369, F(0)=>
      ImgReg4IN_368);
   loop3_23_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_383, D(14)=>
      ImgReg0IN_382, D(13)=>ImgReg0IN_381, D(12)=>ImgReg0IN_380, D(11)=>
      ImgReg0IN_379, D(10)=>ImgReg0IN_378, D(9)=>ImgReg0IN_377, D(8)=>
      ImgReg0IN_376, D(7)=>ImgReg0IN_375, D(6)=>ImgReg0IN_374, D(5)=>
      ImgReg0IN_373, D(4)=>ImgReg0IN_372, D(3)=>ImgReg0IN_371, D(2)=>
      ImgReg0IN_370, D(1)=>ImgReg0IN_369, D(0)=>ImgReg0IN_368, CLK=>nx23966, 
      RST=>RST, EN=>nx23724, Q(15)=>OutputImg0_383_EXMPLR, Q(14)=>
      OutputImg0_382_EXMPLR, Q(13)=>OutputImg0_381_EXMPLR, Q(12)=>
      OutputImg0_380_EXMPLR, Q(11)=>OutputImg0_379_EXMPLR, Q(10)=>
      OutputImg0_378_EXMPLR, Q(9)=>OutputImg0_377_EXMPLR, Q(8)=>
      OutputImg0_376_EXMPLR, Q(7)=>OutputImg0_375_EXMPLR, Q(6)=>
      OutputImg0_374_EXMPLR, Q(5)=>OutputImg0_373_EXMPLR, Q(4)=>
      OutputImg0_372_EXMPLR, Q(3)=>OutputImg0_371_EXMPLR, Q(2)=>
      OutputImg0_370_EXMPLR, Q(1)=>OutputImg0_369_EXMPLR, Q(0)=>
      OutputImg0_368_EXMPLR);
   loop3_23_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_383, D(14)=>
      ImgReg1IN_382, D(13)=>ImgReg1IN_381, D(12)=>ImgReg1IN_380, D(11)=>
      ImgReg1IN_379, D(10)=>ImgReg1IN_378, D(9)=>ImgReg1IN_377, D(8)=>
      ImgReg1IN_376, D(7)=>ImgReg1IN_375, D(6)=>ImgReg1IN_374, D(5)=>
      ImgReg1IN_373, D(4)=>ImgReg1IN_372, D(3)=>ImgReg1IN_371, D(2)=>
      ImgReg1IN_370, D(1)=>ImgReg1IN_369, D(0)=>ImgReg1IN_368, CLK=>nx23968, 
      RST=>RST, EN=>nx23734, Q(15)=>OutputImg1_383_EXMPLR, Q(14)=>
      OutputImg1_382_EXMPLR, Q(13)=>OutputImg1_381_EXMPLR, Q(12)=>
      OutputImg1_380_EXMPLR, Q(11)=>OutputImg1_379_EXMPLR, Q(10)=>
      OutputImg1_378_EXMPLR, Q(9)=>OutputImg1_377_EXMPLR, Q(8)=>
      OutputImg1_376_EXMPLR, Q(7)=>OutputImg1_375_EXMPLR, Q(6)=>
      OutputImg1_374_EXMPLR, Q(5)=>OutputImg1_373_EXMPLR, Q(4)=>
      OutputImg1_372_EXMPLR, Q(3)=>OutputImg1_371_EXMPLR, Q(2)=>
      OutputImg1_370_EXMPLR, Q(1)=>OutputImg1_369_EXMPLR, Q(0)=>
      OutputImg1_368_EXMPLR);
   loop3_23_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_383, D(14)=>
      ImgReg2IN_382, D(13)=>ImgReg2IN_381, D(12)=>ImgReg2IN_380, D(11)=>
      ImgReg2IN_379, D(10)=>ImgReg2IN_378, D(9)=>ImgReg2IN_377, D(8)=>
      ImgReg2IN_376, D(7)=>ImgReg2IN_375, D(6)=>ImgReg2IN_374, D(5)=>
      ImgReg2IN_373, D(4)=>ImgReg2IN_372, D(3)=>ImgReg2IN_371, D(2)=>
      ImgReg2IN_370, D(1)=>ImgReg2IN_369, D(0)=>ImgReg2IN_368, CLK=>nx23968, 
      RST=>RST, EN=>nx23744, Q(15)=>OutputImg2_383_EXMPLR, Q(14)=>
      OutputImg2_382_EXMPLR, Q(13)=>OutputImg2_381_EXMPLR, Q(12)=>
      OutputImg2_380_EXMPLR, Q(11)=>OutputImg2_379_EXMPLR, Q(10)=>
      OutputImg2_378_EXMPLR, Q(9)=>OutputImg2_377_EXMPLR, Q(8)=>
      OutputImg2_376_EXMPLR, Q(7)=>OutputImg2_375_EXMPLR, Q(6)=>
      OutputImg2_374_EXMPLR, Q(5)=>OutputImg2_373_EXMPLR, Q(4)=>
      OutputImg2_372_EXMPLR, Q(3)=>OutputImg2_371_EXMPLR, Q(2)=>
      OutputImg2_370_EXMPLR, Q(1)=>OutputImg2_369_EXMPLR, Q(0)=>
      OutputImg2_368_EXMPLR);
   loop3_23_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_383, D(14)=>
      ImgReg3IN_382, D(13)=>ImgReg3IN_381, D(12)=>ImgReg3IN_380, D(11)=>
      ImgReg3IN_379, D(10)=>ImgReg3IN_378, D(9)=>ImgReg3IN_377, D(8)=>
      ImgReg3IN_376, D(7)=>ImgReg3IN_375, D(6)=>ImgReg3IN_374, D(5)=>
      ImgReg3IN_373, D(4)=>ImgReg3IN_372, D(3)=>ImgReg3IN_371, D(2)=>
      ImgReg3IN_370, D(1)=>ImgReg3IN_369, D(0)=>ImgReg3IN_368, CLK=>nx23970, 
      RST=>RST, EN=>nx23754, Q(15)=>OutputImg3_383_EXMPLR, Q(14)=>
      OutputImg3_382_EXMPLR, Q(13)=>OutputImg3_381_EXMPLR, Q(12)=>
      OutputImg3_380_EXMPLR, Q(11)=>OutputImg3_379_EXMPLR, Q(10)=>
      OutputImg3_378_EXMPLR, Q(9)=>OutputImg3_377_EXMPLR, Q(8)=>
      OutputImg3_376_EXMPLR, Q(7)=>OutputImg3_375_EXMPLR, Q(6)=>
      OutputImg3_374_EXMPLR, Q(5)=>OutputImg3_373_EXMPLR, Q(4)=>
      OutputImg3_372_EXMPLR, Q(3)=>OutputImg3_371_EXMPLR, Q(2)=>
      OutputImg3_370_EXMPLR, Q(1)=>OutputImg3_369_EXMPLR, Q(0)=>
      OutputImg3_368_EXMPLR);
   loop3_23_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_383, D(14)=>
      ImgReg4IN_382, D(13)=>ImgReg4IN_381, D(12)=>ImgReg4IN_380, D(11)=>
      ImgReg4IN_379, D(10)=>ImgReg4IN_378, D(9)=>ImgReg4IN_377, D(8)=>
      ImgReg4IN_376, D(7)=>ImgReg4IN_375, D(6)=>ImgReg4IN_374, D(5)=>
      ImgReg4IN_373, D(4)=>ImgReg4IN_372, D(3)=>ImgReg4IN_371, D(2)=>
      ImgReg4IN_370, D(1)=>ImgReg4IN_369, D(0)=>ImgReg4IN_368, CLK=>nx23970, 
      RST=>RST, EN=>nx23764, Q(15)=>OutputImg4_383_EXMPLR, Q(14)=>
      OutputImg4_382_EXMPLR, Q(13)=>OutputImg4_381_EXMPLR, Q(12)=>
      OutputImg4_380_EXMPLR, Q(11)=>OutputImg4_379_EXMPLR, Q(10)=>
      OutputImg4_378_EXMPLR, Q(9)=>OutputImg4_377_EXMPLR, Q(8)=>
      OutputImg4_376_EXMPLR, Q(7)=>OutputImg4_375_EXMPLR, Q(6)=>
      OutputImg4_374_EXMPLR, Q(5)=>OutputImg4_373_EXMPLR, Q(4)=>
      OutputImg4_372_EXMPLR, Q(3)=>OutputImg4_371_EXMPLR, Q(2)=>
      OutputImg4_370_EXMPLR, Q(1)=>OutputImg4_369_EXMPLR, Q(0)=>
      OutputImg4_368_EXMPLR);
   loop3_23_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_383, D(14)=>
      ImgReg5IN_382, D(13)=>ImgReg5IN_381, D(12)=>ImgReg5IN_380, D(11)=>
      ImgReg5IN_379, D(10)=>ImgReg5IN_378, D(9)=>ImgReg5IN_377, D(8)=>
      ImgReg5IN_376, D(7)=>ImgReg5IN_375, D(6)=>ImgReg5IN_374, D(5)=>
      ImgReg5IN_373, D(4)=>ImgReg5IN_372, D(3)=>ImgReg5IN_371, D(2)=>
      ImgReg5IN_370, D(1)=>ImgReg5IN_369, D(0)=>ImgReg5IN_368, CLK=>nx23972, 
      RST=>RST, EN=>nx23774, Q(15)=>OutputImg5_383_EXMPLR, Q(14)=>
      OutputImg5_382_EXMPLR, Q(13)=>OutputImg5_381_EXMPLR, Q(12)=>
      OutputImg5_380_EXMPLR, Q(11)=>OutputImg5_379_EXMPLR, Q(10)=>
      OutputImg5_378_EXMPLR, Q(9)=>OutputImg5_377_EXMPLR, Q(8)=>
      OutputImg5_376_EXMPLR, Q(7)=>OutputImg5_375_EXMPLR, Q(6)=>
      OutputImg5_374_EXMPLR, Q(5)=>OutputImg5_373_EXMPLR, Q(4)=>
      OutputImg5_372_EXMPLR, Q(3)=>OutputImg5_371_EXMPLR, Q(2)=>
      OutputImg5_370_EXMPLR, Q(1)=>OutputImg5_369_EXMPLR, Q(0)=>
      OutputImg5_368_EXMPLR);
   loop3_24_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_415_EXMPLR, D(14)=>OutputImg0_414_EXMPLR, D(13)=>
      OutputImg0_413_EXMPLR, D(12)=>OutputImg0_412_EXMPLR, D(11)=>
      OutputImg0_411_EXMPLR, D(10)=>OutputImg0_410_EXMPLR, D(9)=>
      OutputImg0_409_EXMPLR, D(8)=>OutputImg0_408_EXMPLR, D(7)=>
      OutputImg0_407_EXMPLR, D(6)=>OutputImg0_406_EXMPLR, D(5)=>
      OutputImg0_405_EXMPLR, D(4)=>OutputImg0_404_EXMPLR, D(3)=>
      OutputImg0_403_EXMPLR, D(2)=>OutputImg0_402_EXMPLR, D(1)=>
      OutputImg0_401_EXMPLR, D(0)=>OutputImg0_400_EXMPLR, EN=>nx23706, F(15)
      =>ImgReg0IN_399, F(14)=>ImgReg0IN_398, F(13)=>ImgReg0IN_397, F(12)=>
      ImgReg0IN_396, F(11)=>ImgReg0IN_395, F(10)=>ImgReg0IN_394, F(9)=>
      ImgReg0IN_393, F(8)=>ImgReg0IN_392, F(7)=>ImgReg0IN_391, F(6)=>
      ImgReg0IN_390, F(5)=>ImgReg0IN_389, F(4)=>ImgReg0IN_388, F(3)=>
      ImgReg0IN_387, F(2)=>ImgReg0IN_386, F(1)=>ImgReg0IN_385, F(0)=>
      ImgReg0IN_384);
   loop3_24_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_415_EXMPLR, D(14)=>OutputImg1_414_EXMPLR, D(13)=>
      OutputImg1_413_EXMPLR, D(12)=>OutputImg1_412_EXMPLR, D(11)=>
      OutputImg1_411_EXMPLR, D(10)=>OutputImg1_410_EXMPLR, D(9)=>
      OutputImg1_409_EXMPLR, D(8)=>OutputImg1_408_EXMPLR, D(7)=>
      OutputImg1_407_EXMPLR, D(6)=>OutputImg1_406_EXMPLR, D(5)=>
      OutputImg1_405_EXMPLR, D(4)=>OutputImg1_404_EXMPLR, D(3)=>
      OutputImg1_403_EXMPLR, D(2)=>OutputImg1_402_EXMPLR, D(1)=>
      OutputImg1_401_EXMPLR, D(0)=>OutputImg1_400_EXMPLR, EN=>nx23706, F(15)
      =>ImgReg1IN_399, F(14)=>ImgReg1IN_398, F(13)=>ImgReg1IN_397, F(12)=>
      ImgReg1IN_396, F(11)=>ImgReg1IN_395, F(10)=>ImgReg1IN_394, F(9)=>
      ImgReg1IN_393, F(8)=>ImgReg1IN_392, F(7)=>ImgReg1IN_391, F(6)=>
      ImgReg1IN_390, F(5)=>ImgReg1IN_389, F(4)=>ImgReg1IN_388, F(3)=>
      ImgReg1IN_387, F(2)=>ImgReg1IN_386, F(1)=>ImgReg1IN_385, F(0)=>
      ImgReg1IN_384);
   loop3_24_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_415_EXMPLR, D(14)=>OutputImg2_414_EXMPLR, D(13)=>
      OutputImg2_413_EXMPLR, D(12)=>OutputImg2_412_EXMPLR, D(11)=>
      OutputImg2_411_EXMPLR, D(10)=>OutputImg2_410_EXMPLR, D(9)=>
      OutputImg2_409_EXMPLR, D(8)=>OutputImg2_408_EXMPLR, D(7)=>
      OutputImg2_407_EXMPLR, D(6)=>OutputImg2_406_EXMPLR, D(5)=>
      OutputImg2_405_EXMPLR, D(4)=>OutputImg2_404_EXMPLR, D(3)=>
      OutputImg2_403_EXMPLR, D(2)=>OutputImg2_402_EXMPLR, D(1)=>
      OutputImg2_401_EXMPLR, D(0)=>OutputImg2_400_EXMPLR, EN=>nx23706, F(15)
      =>ImgReg2IN_399, F(14)=>ImgReg2IN_398, F(13)=>ImgReg2IN_397, F(12)=>
      ImgReg2IN_396, F(11)=>ImgReg2IN_395, F(10)=>ImgReg2IN_394, F(9)=>
      ImgReg2IN_393, F(8)=>ImgReg2IN_392, F(7)=>ImgReg2IN_391, F(6)=>
      ImgReg2IN_390, F(5)=>ImgReg2IN_389, F(4)=>ImgReg2IN_388, F(3)=>
      ImgReg2IN_387, F(2)=>ImgReg2IN_386, F(1)=>ImgReg2IN_385, F(0)=>
      ImgReg2IN_384);
   loop3_24_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_415_EXMPLR, D(14)=>OutputImg3_414_EXMPLR, D(13)=>
      OutputImg3_413_EXMPLR, D(12)=>OutputImg3_412_EXMPLR, D(11)=>
      OutputImg3_411_EXMPLR, D(10)=>OutputImg3_410_EXMPLR, D(9)=>
      OutputImg3_409_EXMPLR, D(8)=>OutputImg3_408_EXMPLR, D(7)=>
      OutputImg3_407_EXMPLR, D(6)=>OutputImg3_406_EXMPLR, D(5)=>
      OutputImg3_405_EXMPLR, D(4)=>OutputImg3_404_EXMPLR, D(3)=>
      OutputImg3_403_EXMPLR, D(2)=>OutputImg3_402_EXMPLR, D(1)=>
      OutputImg3_401_EXMPLR, D(0)=>OutputImg3_400_EXMPLR, EN=>nx23708, F(15)
      =>ImgReg3IN_399, F(14)=>ImgReg3IN_398, F(13)=>ImgReg3IN_397, F(12)=>
      ImgReg3IN_396, F(11)=>ImgReg3IN_395, F(10)=>ImgReg3IN_394, F(9)=>
      ImgReg3IN_393, F(8)=>ImgReg3IN_392, F(7)=>ImgReg3IN_391, F(6)=>
      ImgReg3IN_390, F(5)=>ImgReg3IN_389, F(4)=>ImgReg3IN_388, F(3)=>
      ImgReg3IN_387, F(2)=>ImgReg3IN_386, F(1)=>ImgReg3IN_385, F(0)=>
      ImgReg3IN_384);
   loop3_24_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_415_EXMPLR, D(14)=>OutputImg4_414_EXMPLR, D(13)=>
      OutputImg4_413_EXMPLR, D(12)=>OutputImg4_412_EXMPLR, D(11)=>
      OutputImg4_411_EXMPLR, D(10)=>OutputImg4_410_EXMPLR, D(9)=>
      OutputImg4_409_EXMPLR, D(8)=>OutputImg4_408_EXMPLR, D(7)=>
      OutputImg4_407_EXMPLR, D(6)=>OutputImg4_406_EXMPLR, D(5)=>
      OutputImg4_405_EXMPLR, D(4)=>OutputImg4_404_EXMPLR, D(3)=>
      OutputImg4_403_EXMPLR, D(2)=>OutputImg4_402_EXMPLR, D(1)=>
      OutputImg4_401_EXMPLR, D(0)=>OutputImg4_400_EXMPLR, EN=>nx23708, F(15)
      =>ImgReg4IN_399, F(14)=>ImgReg4IN_398, F(13)=>ImgReg4IN_397, F(12)=>
      ImgReg4IN_396, F(11)=>ImgReg4IN_395, F(10)=>ImgReg4IN_394, F(9)=>
      ImgReg4IN_393, F(8)=>ImgReg4IN_392, F(7)=>ImgReg4IN_391, F(6)=>
      ImgReg4IN_390, F(5)=>ImgReg4IN_389, F(4)=>ImgReg4IN_388, F(3)=>
      ImgReg4IN_387, F(2)=>ImgReg4IN_386, F(1)=>ImgReg4IN_385, F(0)=>
      ImgReg4IN_384);
   loop3_24_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_415_EXMPLR, D(14)=>OutputImg5_414_EXMPLR, D(13)=>
      OutputImg5_413_EXMPLR, D(12)=>OutputImg5_412_EXMPLR, D(11)=>
      OutputImg5_411_EXMPLR, D(10)=>OutputImg5_410_EXMPLR, D(9)=>
      OutputImg5_409_EXMPLR, D(8)=>OutputImg5_408_EXMPLR, D(7)=>
      OutputImg5_407_EXMPLR, D(6)=>OutputImg5_406_EXMPLR, D(5)=>
      OutputImg5_405_EXMPLR, D(4)=>OutputImg5_404_EXMPLR, D(3)=>
      OutputImg5_403_EXMPLR, D(2)=>OutputImg5_402_EXMPLR, D(1)=>
      OutputImg5_401_EXMPLR, D(0)=>OutputImg5_400_EXMPLR, EN=>nx23708, F(15)
      =>ImgReg5IN_399, F(14)=>ImgReg5IN_398, F(13)=>ImgReg5IN_397, F(12)=>
      ImgReg5IN_396, F(11)=>ImgReg5IN_395, F(10)=>ImgReg5IN_394, F(9)=>
      ImgReg5IN_393, F(8)=>ImgReg5IN_392, F(7)=>ImgReg5IN_391, F(6)=>
      ImgReg5IN_390, F(5)=>ImgReg5IN_389, F(4)=>ImgReg5IN_388, F(3)=>
      ImgReg5IN_387, F(2)=>ImgReg5IN_386, F(1)=>ImgReg5IN_385, F(0)=>
      ImgReg5IN_384);
   loop3_24_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(399), 
      D(14)=>DATA(398), D(13)=>DATA(397), D(12)=>DATA(396), D(11)=>DATA(395), 
      D(10)=>DATA(394), D(9)=>DATA(393), D(8)=>DATA(392), D(7)=>DATA(391), 
      D(6)=>DATA(390), D(5)=>DATA(389), D(4)=>DATA(388), D(3)=>DATA(387), 
      D(2)=>DATA(386), D(1)=>DATA(385), D(0)=>DATA(384), EN=>nx23660, F(15)
      =>ImgReg0IN_399, F(14)=>ImgReg0IN_398, F(13)=>ImgReg0IN_397, F(12)=>
      ImgReg0IN_396, F(11)=>ImgReg0IN_395, F(10)=>ImgReg0IN_394, F(9)=>
      ImgReg0IN_393, F(8)=>ImgReg0IN_392, F(7)=>ImgReg0IN_391, F(6)=>
      ImgReg0IN_390, F(5)=>ImgReg0IN_389, F(4)=>ImgReg0IN_388, F(3)=>
      ImgReg0IN_387, F(2)=>ImgReg0IN_386, F(1)=>ImgReg0IN_385, F(0)=>
      ImgReg0IN_384);
   loop3_24_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(399), 
      D(14)=>DATA(398), D(13)=>DATA(397), D(12)=>DATA(396), D(11)=>DATA(395), 
      D(10)=>DATA(394), D(9)=>DATA(393), D(8)=>DATA(392), D(7)=>DATA(391), 
      D(6)=>DATA(390), D(5)=>DATA(389), D(4)=>DATA(388), D(3)=>DATA(387), 
      D(2)=>DATA(386), D(1)=>DATA(385), D(0)=>DATA(384), EN=>nx23648, F(15)
      =>ImgReg1IN_399, F(14)=>ImgReg1IN_398, F(13)=>ImgReg1IN_397, F(12)=>
      ImgReg1IN_396, F(11)=>ImgReg1IN_395, F(10)=>ImgReg1IN_394, F(9)=>
      ImgReg1IN_393, F(8)=>ImgReg1IN_392, F(7)=>ImgReg1IN_391, F(6)=>
      ImgReg1IN_390, F(5)=>ImgReg1IN_389, F(4)=>ImgReg1IN_388, F(3)=>
      ImgReg1IN_387, F(2)=>ImgReg1IN_386, F(1)=>ImgReg1IN_385, F(0)=>
      ImgReg1IN_384);
   loop3_24_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(399), 
      D(14)=>DATA(398), D(13)=>DATA(397), D(12)=>DATA(396), D(11)=>DATA(395), 
      D(10)=>DATA(394), D(9)=>DATA(393), D(8)=>DATA(392), D(7)=>DATA(391), 
      D(6)=>DATA(390), D(5)=>DATA(389), D(4)=>DATA(388), D(3)=>DATA(387), 
      D(2)=>DATA(386), D(1)=>DATA(385), D(0)=>DATA(384), EN=>nx23636, F(15)
      =>ImgReg2IN_399, F(14)=>ImgReg2IN_398, F(13)=>ImgReg2IN_397, F(12)=>
      ImgReg2IN_396, F(11)=>ImgReg2IN_395, F(10)=>ImgReg2IN_394, F(9)=>
      ImgReg2IN_393, F(8)=>ImgReg2IN_392, F(7)=>ImgReg2IN_391, F(6)=>
      ImgReg2IN_390, F(5)=>ImgReg2IN_389, F(4)=>ImgReg2IN_388, F(3)=>
      ImgReg2IN_387, F(2)=>ImgReg2IN_386, F(1)=>ImgReg2IN_385, F(0)=>
      ImgReg2IN_384);
   loop3_24_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(399), 
      D(14)=>DATA(398), D(13)=>DATA(397), D(12)=>DATA(396), D(11)=>DATA(395), 
      D(10)=>DATA(394), D(9)=>DATA(393), D(8)=>DATA(392), D(7)=>DATA(391), 
      D(6)=>DATA(390), D(5)=>DATA(389), D(4)=>DATA(388), D(3)=>DATA(387), 
      D(2)=>DATA(386), D(1)=>DATA(385), D(0)=>DATA(384), EN=>nx23624, F(15)
      =>ImgReg3IN_399, F(14)=>ImgReg3IN_398, F(13)=>ImgReg3IN_397, F(12)=>
      ImgReg3IN_396, F(11)=>ImgReg3IN_395, F(10)=>ImgReg3IN_394, F(9)=>
      ImgReg3IN_393, F(8)=>ImgReg3IN_392, F(7)=>ImgReg3IN_391, F(6)=>
      ImgReg3IN_390, F(5)=>ImgReg3IN_389, F(4)=>ImgReg3IN_388, F(3)=>
      ImgReg3IN_387, F(2)=>ImgReg3IN_386, F(1)=>ImgReg3IN_385, F(0)=>
      ImgReg3IN_384);
   loop3_24_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(399), 
      D(14)=>DATA(398), D(13)=>DATA(397), D(12)=>DATA(396), D(11)=>DATA(395), 
      D(10)=>DATA(394), D(9)=>DATA(393), D(8)=>DATA(392), D(7)=>DATA(391), 
      D(6)=>DATA(390), D(5)=>DATA(389), D(4)=>DATA(388), D(3)=>DATA(387), 
      D(2)=>DATA(386), D(1)=>DATA(385), D(0)=>DATA(384), EN=>nx23612, F(15)
      =>ImgReg4IN_399, F(14)=>ImgReg4IN_398, F(13)=>ImgReg4IN_397, F(12)=>
      ImgReg4IN_396, F(11)=>ImgReg4IN_395, F(10)=>ImgReg4IN_394, F(9)=>
      ImgReg4IN_393, F(8)=>ImgReg4IN_392, F(7)=>ImgReg4IN_391, F(6)=>
      ImgReg4IN_390, F(5)=>ImgReg4IN_389, F(4)=>ImgReg4IN_388, F(3)=>
      ImgReg4IN_387, F(2)=>ImgReg4IN_386, F(1)=>ImgReg4IN_385, F(0)=>
      ImgReg4IN_384);
   loop3_24_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(399), 
      D(14)=>DATA(398), D(13)=>DATA(397), D(12)=>DATA(396), D(11)=>DATA(395), 
      D(10)=>DATA(394), D(9)=>DATA(393), D(8)=>DATA(392), D(7)=>DATA(391), 
      D(6)=>DATA(390), D(5)=>DATA(389), D(4)=>DATA(388), D(3)=>DATA(387), 
      D(2)=>DATA(386), D(1)=>DATA(385), D(0)=>DATA(384), EN=>nx23600, F(15)
      =>ImgReg5IN_399, F(14)=>ImgReg5IN_398, F(13)=>ImgReg5IN_397, F(12)=>
      ImgReg5IN_396, F(11)=>ImgReg5IN_395, F(10)=>ImgReg5IN_394, F(9)=>
      ImgReg5IN_393, F(8)=>ImgReg5IN_392, F(7)=>ImgReg5IN_391, F(6)=>
      ImgReg5IN_390, F(5)=>ImgReg5IN_389, F(4)=>ImgReg5IN_388, F(3)=>
      ImgReg5IN_387, F(2)=>ImgReg5IN_386, F(1)=>ImgReg5IN_385, F(0)=>
      ImgReg5IN_384);
   loop3_24_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_399_EXMPLR, D(14)=>OutputImg1_398_EXMPLR, D(13)=>
      OutputImg1_397_EXMPLR, D(12)=>OutputImg1_396_EXMPLR, D(11)=>
      OutputImg1_395_EXMPLR, D(10)=>OutputImg1_394_EXMPLR, D(9)=>
      OutputImg1_393_EXMPLR, D(8)=>OutputImg1_392_EXMPLR, D(7)=>
      OutputImg1_391_EXMPLR, D(6)=>OutputImg1_390_EXMPLR, D(5)=>
      OutputImg1_389_EXMPLR, D(4)=>OutputImg1_388_EXMPLR, D(3)=>
      OutputImg1_387_EXMPLR, D(2)=>OutputImg1_386_EXMPLR, D(1)=>
      OutputImg1_385_EXMPLR, D(0)=>OutputImg1_384_EXMPLR, EN=>nx23820, F(15)
      =>ImgReg0IN_399, F(14)=>ImgReg0IN_398, F(13)=>ImgReg0IN_397, F(12)=>
      ImgReg0IN_396, F(11)=>ImgReg0IN_395, F(10)=>ImgReg0IN_394, F(9)=>
      ImgReg0IN_393, F(8)=>ImgReg0IN_392, F(7)=>ImgReg0IN_391, F(6)=>
      ImgReg0IN_390, F(5)=>ImgReg0IN_389, F(4)=>ImgReg0IN_388, F(3)=>
      ImgReg0IN_387, F(2)=>ImgReg0IN_386, F(1)=>ImgReg0IN_385, F(0)=>
      ImgReg0IN_384);
   loop3_24_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_399_EXMPLR, D(14)=>OutputImg2_398_EXMPLR, D(13)=>
      OutputImg2_397_EXMPLR, D(12)=>OutputImg2_396_EXMPLR, D(11)=>
      OutputImg2_395_EXMPLR, D(10)=>OutputImg2_394_EXMPLR, D(9)=>
      OutputImg2_393_EXMPLR, D(8)=>OutputImg2_392_EXMPLR, D(7)=>
      OutputImg2_391_EXMPLR, D(6)=>OutputImg2_390_EXMPLR, D(5)=>
      OutputImg2_389_EXMPLR, D(4)=>OutputImg2_388_EXMPLR, D(3)=>
      OutputImg2_387_EXMPLR, D(2)=>OutputImg2_386_EXMPLR, D(1)=>
      OutputImg2_385_EXMPLR, D(0)=>OutputImg2_384_EXMPLR, EN=>nx23820, F(15)
      =>ImgReg1IN_399, F(14)=>ImgReg1IN_398, F(13)=>ImgReg1IN_397, F(12)=>
      ImgReg1IN_396, F(11)=>ImgReg1IN_395, F(10)=>ImgReg1IN_394, F(9)=>
      ImgReg1IN_393, F(8)=>ImgReg1IN_392, F(7)=>ImgReg1IN_391, F(6)=>
      ImgReg1IN_390, F(5)=>ImgReg1IN_389, F(4)=>ImgReg1IN_388, F(3)=>
      ImgReg1IN_387, F(2)=>ImgReg1IN_386, F(1)=>ImgReg1IN_385, F(0)=>
      ImgReg1IN_384);
   loop3_24_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_399_EXMPLR, D(14)=>OutputImg3_398_EXMPLR, D(13)=>
      OutputImg3_397_EXMPLR, D(12)=>OutputImg3_396_EXMPLR, D(11)=>
      OutputImg3_395_EXMPLR, D(10)=>OutputImg3_394_EXMPLR, D(9)=>
      OutputImg3_393_EXMPLR, D(8)=>OutputImg3_392_EXMPLR, D(7)=>
      OutputImg3_391_EXMPLR, D(6)=>OutputImg3_390_EXMPLR, D(5)=>
      OutputImg3_389_EXMPLR, D(4)=>OutputImg3_388_EXMPLR, D(3)=>
      OutputImg3_387_EXMPLR, D(2)=>OutputImg3_386_EXMPLR, D(1)=>
      OutputImg3_385_EXMPLR, D(0)=>OutputImg3_384_EXMPLR, EN=>nx23820, F(15)
      =>ImgReg2IN_399, F(14)=>ImgReg2IN_398, F(13)=>ImgReg2IN_397, F(12)=>
      ImgReg2IN_396, F(11)=>ImgReg2IN_395, F(10)=>ImgReg2IN_394, F(9)=>
      ImgReg2IN_393, F(8)=>ImgReg2IN_392, F(7)=>ImgReg2IN_391, F(6)=>
      ImgReg2IN_390, F(5)=>ImgReg2IN_389, F(4)=>ImgReg2IN_388, F(3)=>
      ImgReg2IN_387, F(2)=>ImgReg2IN_386, F(1)=>ImgReg2IN_385, F(0)=>
      ImgReg2IN_384);
   loop3_24_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_399_EXMPLR, D(14)=>OutputImg4_398_EXMPLR, D(13)=>
      OutputImg4_397_EXMPLR, D(12)=>OutputImg4_396_EXMPLR, D(11)=>
      OutputImg4_395_EXMPLR, D(10)=>OutputImg4_394_EXMPLR, D(9)=>
      OutputImg4_393_EXMPLR, D(8)=>OutputImg4_392_EXMPLR, D(7)=>
      OutputImg4_391_EXMPLR, D(6)=>OutputImg4_390_EXMPLR, D(5)=>
      OutputImg4_389_EXMPLR, D(4)=>OutputImg4_388_EXMPLR, D(3)=>
      OutputImg4_387_EXMPLR, D(2)=>OutputImg4_386_EXMPLR, D(1)=>
      OutputImg4_385_EXMPLR, D(0)=>OutputImg4_384_EXMPLR, EN=>nx23820, F(15)
      =>ImgReg3IN_399, F(14)=>ImgReg3IN_398, F(13)=>ImgReg3IN_397, F(12)=>
      ImgReg3IN_396, F(11)=>ImgReg3IN_395, F(10)=>ImgReg3IN_394, F(9)=>
      ImgReg3IN_393, F(8)=>ImgReg3IN_392, F(7)=>ImgReg3IN_391, F(6)=>
      ImgReg3IN_390, F(5)=>ImgReg3IN_389, F(4)=>ImgReg3IN_388, F(3)=>
      ImgReg3IN_387, F(2)=>ImgReg3IN_386, F(1)=>ImgReg3IN_385, F(0)=>
      ImgReg3IN_384);
   loop3_24_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_399_EXMPLR, D(14)=>OutputImg5_398_EXMPLR, D(13)=>
      OutputImg5_397_EXMPLR, D(12)=>OutputImg5_396_EXMPLR, D(11)=>
      OutputImg5_395_EXMPLR, D(10)=>OutputImg5_394_EXMPLR, D(9)=>
      OutputImg5_393_EXMPLR, D(8)=>OutputImg5_392_EXMPLR, D(7)=>
      OutputImg5_391_EXMPLR, D(6)=>OutputImg5_390_EXMPLR, D(5)=>
      OutputImg5_389_EXMPLR, D(4)=>OutputImg5_388_EXMPLR, D(3)=>
      OutputImg5_387_EXMPLR, D(2)=>OutputImg5_386_EXMPLR, D(1)=>
      OutputImg5_385_EXMPLR, D(0)=>OutputImg5_384_EXMPLR, EN=>nx23820, F(15)
      =>ImgReg4IN_399, F(14)=>ImgReg4IN_398, F(13)=>ImgReg4IN_397, F(12)=>
      ImgReg4IN_396, F(11)=>ImgReg4IN_395, F(10)=>ImgReg4IN_394, F(9)=>
      ImgReg4IN_393, F(8)=>ImgReg4IN_392, F(7)=>ImgReg4IN_391, F(6)=>
      ImgReg4IN_390, F(5)=>ImgReg4IN_389, F(4)=>ImgReg4IN_388, F(3)=>
      ImgReg4IN_387, F(2)=>ImgReg4IN_386, F(1)=>ImgReg4IN_385, F(0)=>
      ImgReg4IN_384);
   loop3_24_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_399, D(14)=>
      ImgReg0IN_398, D(13)=>ImgReg0IN_397, D(12)=>ImgReg0IN_396, D(11)=>
      ImgReg0IN_395, D(10)=>ImgReg0IN_394, D(9)=>ImgReg0IN_393, D(8)=>
      ImgReg0IN_392, D(7)=>ImgReg0IN_391, D(6)=>ImgReg0IN_390, D(5)=>
      ImgReg0IN_389, D(4)=>ImgReg0IN_388, D(3)=>ImgReg0IN_387, D(2)=>
      ImgReg0IN_386, D(1)=>ImgReg0IN_385, D(0)=>ImgReg0IN_384, CLK=>nx23972, 
      RST=>RST, EN=>nx23724, Q(15)=>OutputImg0_399_EXMPLR, Q(14)=>
      OutputImg0_398_EXMPLR, Q(13)=>OutputImg0_397_EXMPLR, Q(12)=>
      OutputImg0_396_EXMPLR, Q(11)=>OutputImg0_395_EXMPLR, Q(10)=>
      OutputImg0_394_EXMPLR, Q(9)=>OutputImg0_393_EXMPLR, Q(8)=>
      OutputImg0_392_EXMPLR, Q(7)=>OutputImg0_391_EXMPLR, Q(6)=>
      OutputImg0_390_EXMPLR, Q(5)=>OutputImg0_389_EXMPLR, Q(4)=>
      OutputImg0_388_EXMPLR, Q(3)=>OutputImg0_387_EXMPLR, Q(2)=>
      OutputImg0_386_EXMPLR, Q(1)=>OutputImg0_385_EXMPLR, Q(0)=>
      OutputImg0_384_EXMPLR);
   loop3_24_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_399, D(14)=>
      ImgReg1IN_398, D(13)=>ImgReg1IN_397, D(12)=>ImgReg1IN_396, D(11)=>
      ImgReg1IN_395, D(10)=>ImgReg1IN_394, D(9)=>ImgReg1IN_393, D(8)=>
      ImgReg1IN_392, D(7)=>ImgReg1IN_391, D(6)=>ImgReg1IN_390, D(5)=>
      ImgReg1IN_389, D(4)=>ImgReg1IN_388, D(3)=>ImgReg1IN_387, D(2)=>
      ImgReg1IN_386, D(1)=>ImgReg1IN_385, D(0)=>ImgReg1IN_384, CLK=>nx23974, 
      RST=>RST, EN=>nx23734, Q(15)=>OutputImg1_399_EXMPLR, Q(14)=>
      OutputImg1_398_EXMPLR, Q(13)=>OutputImg1_397_EXMPLR, Q(12)=>
      OutputImg1_396_EXMPLR, Q(11)=>OutputImg1_395_EXMPLR, Q(10)=>
      OutputImg1_394_EXMPLR, Q(9)=>OutputImg1_393_EXMPLR, Q(8)=>
      OutputImg1_392_EXMPLR, Q(7)=>OutputImg1_391_EXMPLR, Q(6)=>
      OutputImg1_390_EXMPLR, Q(5)=>OutputImg1_389_EXMPLR, Q(4)=>
      OutputImg1_388_EXMPLR, Q(3)=>OutputImg1_387_EXMPLR, Q(2)=>
      OutputImg1_386_EXMPLR, Q(1)=>OutputImg1_385_EXMPLR, Q(0)=>
      OutputImg1_384_EXMPLR);
   loop3_24_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_399, D(14)=>
      ImgReg2IN_398, D(13)=>ImgReg2IN_397, D(12)=>ImgReg2IN_396, D(11)=>
      ImgReg2IN_395, D(10)=>ImgReg2IN_394, D(9)=>ImgReg2IN_393, D(8)=>
      ImgReg2IN_392, D(7)=>ImgReg2IN_391, D(6)=>ImgReg2IN_390, D(5)=>
      ImgReg2IN_389, D(4)=>ImgReg2IN_388, D(3)=>ImgReg2IN_387, D(2)=>
      ImgReg2IN_386, D(1)=>ImgReg2IN_385, D(0)=>ImgReg2IN_384, CLK=>nx23974, 
      RST=>RST, EN=>nx23744, Q(15)=>OutputImg2_399_EXMPLR, Q(14)=>
      OutputImg2_398_EXMPLR, Q(13)=>OutputImg2_397_EXMPLR, Q(12)=>
      OutputImg2_396_EXMPLR, Q(11)=>OutputImg2_395_EXMPLR, Q(10)=>
      OutputImg2_394_EXMPLR, Q(9)=>OutputImg2_393_EXMPLR, Q(8)=>
      OutputImg2_392_EXMPLR, Q(7)=>OutputImg2_391_EXMPLR, Q(6)=>
      OutputImg2_390_EXMPLR, Q(5)=>OutputImg2_389_EXMPLR, Q(4)=>
      OutputImg2_388_EXMPLR, Q(3)=>OutputImg2_387_EXMPLR, Q(2)=>
      OutputImg2_386_EXMPLR, Q(1)=>OutputImg2_385_EXMPLR, Q(0)=>
      OutputImg2_384_EXMPLR);
   loop3_24_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_399, D(14)=>
      ImgReg3IN_398, D(13)=>ImgReg3IN_397, D(12)=>ImgReg3IN_396, D(11)=>
      ImgReg3IN_395, D(10)=>ImgReg3IN_394, D(9)=>ImgReg3IN_393, D(8)=>
      ImgReg3IN_392, D(7)=>ImgReg3IN_391, D(6)=>ImgReg3IN_390, D(5)=>
      ImgReg3IN_389, D(4)=>ImgReg3IN_388, D(3)=>ImgReg3IN_387, D(2)=>
      ImgReg3IN_386, D(1)=>ImgReg3IN_385, D(0)=>ImgReg3IN_384, CLK=>nx23976, 
      RST=>RST, EN=>nx23754, Q(15)=>OutputImg3_399_EXMPLR, Q(14)=>
      OutputImg3_398_EXMPLR, Q(13)=>OutputImg3_397_EXMPLR, Q(12)=>
      OutputImg3_396_EXMPLR, Q(11)=>OutputImg3_395_EXMPLR, Q(10)=>
      OutputImg3_394_EXMPLR, Q(9)=>OutputImg3_393_EXMPLR, Q(8)=>
      OutputImg3_392_EXMPLR, Q(7)=>OutputImg3_391_EXMPLR, Q(6)=>
      OutputImg3_390_EXMPLR, Q(5)=>OutputImg3_389_EXMPLR, Q(4)=>
      OutputImg3_388_EXMPLR, Q(3)=>OutputImg3_387_EXMPLR, Q(2)=>
      OutputImg3_386_EXMPLR, Q(1)=>OutputImg3_385_EXMPLR, Q(0)=>
      OutputImg3_384_EXMPLR);
   loop3_24_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_399, D(14)=>
      ImgReg4IN_398, D(13)=>ImgReg4IN_397, D(12)=>ImgReg4IN_396, D(11)=>
      ImgReg4IN_395, D(10)=>ImgReg4IN_394, D(9)=>ImgReg4IN_393, D(8)=>
      ImgReg4IN_392, D(7)=>ImgReg4IN_391, D(6)=>ImgReg4IN_390, D(5)=>
      ImgReg4IN_389, D(4)=>ImgReg4IN_388, D(3)=>ImgReg4IN_387, D(2)=>
      ImgReg4IN_386, D(1)=>ImgReg4IN_385, D(0)=>ImgReg4IN_384, CLK=>nx23976, 
      RST=>RST, EN=>nx23764, Q(15)=>OutputImg4_399_EXMPLR, Q(14)=>
      OutputImg4_398_EXMPLR, Q(13)=>OutputImg4_397_EXMPLR, Q(12)=>
      OutputImg4_396_EXMPLR, Q(11)=>OutputImg4_395_EXMPLR, Q(10)=>
      OutputImg4_394_EXMPLR, Q(9)=>OutputImg4_393_EXMPLR, Q(8)=>
      OutputImg4_392_EXMPLR, Q(7)=>OutputImg4_391_EXMPLR, Q(6)=>
      OutputImg4_390_EXMPLR, Q(5)=>OutputImg4_389_EXMPLR, Q(4)=>
      OutputImg4_388_EXMPLR, Q(3)=>OutputImg4_387_EXMPLR, Q(2)=>
      OutputImg4_386_EXMPLR, Q(1)=>OutputImg4_385_EXMPLR, Q(0)=>
      OutputImg4_384_EXMPLR);
   loop3_24_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_399, D(14)=>
      ImgReg5IN_398, D(13)=>ImgReg5IN_397, D(12)=>ImgReg5IN_396, D(11)=>
      ImgReg5IN_395, D(10)=>ImgReg5IN_394, D(9)=>ImgReg5IN_393, D(8)=>
      ImgReg5IN_392, D(7)=>ImgReg5IN_391, D(6)=>ImgReg5IN_390, D(5)=>
      ImgReg5IN_389, D(4)=>ImgReg5IN_388, D(3)=>ImgReg5IN_387, D(2)=>
      ImgReg5IN_386, D(1)=>ImgReg5IN_385, D(0)=>ImgReg5IN_384, CLK=>nx23978, 
      RST=>RST, EN=>nx23774, Q(15)=>OutputImg5_399_EXMPLR, Q(14)=>
      OutputImg5_398_EXMPLR, Q(13)=>OutputImg5_397_EXMPLR, Q(12)=>
      OutputImg5_396_EXMPLR, Q(11)=>OutputImg5_395_EXMPLR, Q(10)=>
      OutputImg5_394_EXMPLR, Q(9)=>OutputImg5_393_EXMPLR, Q(8)=>
      OutputImg5_392_EXMPLR, Q(7)=>OutputImg5_391_EXMPLR, Q(6)=>
      OutputImg5_390_EXMPLR, Q(5)=>OutputImg5_389_EXMPLR, Q(4)=>
      OutputImg5_388_EXMPLR, Q(3)=>OutputImg5_387_EXMPLR, Q(2)=>
      OutputImg5_386_EXMPLR, Q(1)=>OutputImg5_385_EXMPLR, Q(0)=>
      OutputImg5_384_EXMPLR);
   loop3_25_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_431_EXMPLR, D(14)=>OutputImg0_430_EXMPLR, D(13)=>
      OutputImg0_429_EXMPLR, D(12)=>OutputImg0_428_EXMPLR, D(11)=>
      OutputImg0_427_EXMPLR, D(10)=>OutputImg0_426_EXMPLR, D(9)=>
      OutputImg0_425_EXMPLR, D(8)=>OutputImg0_424_EXMPLR, D(7)=>
      OutputImg0_423_EXMPLR, D(6)=>OutputImg0_422_EXMPLR, D(5)=>
      OutputImg0_421_EXMPLR, D(4)=>OutputImg0_420_EXMPLR, D(3)=>
      OutputImg0_419_EXMPLR, D(2)=>OutputImg0_418_EXMPLR, D(1)=>
      OutputImg0_417_EXMPLR, D(0)=>OutputImg0_416_EXMPLR, EN=>nx23708, F(15)
      =>ImgReg0IN_415, F(14)=>ImgReg0IN_414, F(13)=>ImgReg0IN_413, F(12)=>
      ImgReg0IN_412, F(11)=>ImgReg0IN_411, F(10)=>ImgReg0IN_410, F(9)=>
      ImgReg0IN_409, F(8)=>ImgReg0IN_408, F(7)=>ImgReg0IN_407, F(6)=>
      ImgReg0IN_406, F(5)=>ImgReg0IN_405, F(4)=>ImgReg0IN_404, F(3)=>
      ImgReg0IN_403, F(2)=>ImgReg0IN_402, F(1)=>ImgReg0IN_401, F(0)=>
      ImgReg0IN_400);
   loop3_25_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_431_EXMPLR, D(14)=>OutputImg1_430_EXMPLR, D(13)=>
      OutputImg1_429_EXMPLR, D(12)=>OutputImg1_428_EXMPLR, D(11)=>
      OutputImg1_427_EXMPLR, D(10)=>OutputImg1_426_EXMPLR, D(9)=>
      OutputImg1_425_EXMPLR, D(8)=>OutputImg1_424_EXMPLR, D(7)=>
      OutputImg1_423_EXMPLR, D(6)=>OutputImg1_422_EXMPLR, D(5)=>
      OutputImg1_421_EXMPLR, D(4)=>OutputImg1_420_EXMPLR, D(3)=>
      OutputImg1_419_EXMPLR, D(2)=>OutputImg1_418_EXMPLR, D(1)=>
      OutputImg1_417_EXMPLR, D(0)=>OutputImg1_416_EXMPLR, EN=>nx23708, F(15)
      =>ImgReg1IN_415, F(14)=>ImgReg1IN_414, F(13)=>ImgReg1IN_413, F(12)=>
      ImgReg1IN_412, F(11)=>ImgReg1IN_411, F(10)=>ImgReg1IN_410, F(9)=>
      ImgReg1IN_409, F(8)=>ImgReg1IN_408, F(7)=>ImgReg1IN_407, F(6)=>
      ImgReg1IN_406, F(5)=>ImgReg1IN_405, F(4)=>ImgReg1IN_404, F(3)=>
      ImgReg1IN_403, F(2)=>ImgReg1IN_402, F(1)=>ImgReg1IN_401, F(0)=>
      ImgReg1IN_400);
   loop3_25_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_431_EXMPLR, D(14)=>OutputImg2_430_EXMPLR, D(13)=>
      OutputImg2_429_EXMPLR, D(12)=>OutputImg2_428_EXMPLR, D(11)=>
      OutputImg2_427_EXMPLR, D(10)=>OutputImg2_426_EXMPLR, D(9)=>
      OutputImg2_425_EXMPLR, D(8)=>OutputImg2_424_EXMPLR, D(7)=>
      OutputImg2_423_EXMPLR, D(6)=>OutputImg2_422_EXMPLR, D(5)=>
      OutputImg2_421_EXMPLR, D(4)=>OutputImg2_420_EXMPLR, D(3)=>
      OutputImg2_419_EXMPLR, D(2)=>OutputImg2_418_EXMPLR, D(1)=>
      OutputImg2_417_EXMPLR, D(0)=>OutputImg2_416_EXMPLR, EN=>nx23708, F(15)
      =>ImgReg2IN_415, F(14)=>ImgReg2IN_414, F(13)=>ImgReg2IN_413, F(12)=>
      ImgReg2IN_412, F(11)=>ImgReg2IN_411, F(10)=>ImgReg2IN_410, F(9)=>
      ImgReg2IN_409, F(8)=>ImgReg2IN_408, F(7)=>ImgReg2IN_407, F(6)=>
      ImgReg2IN_406, F(5)=>ImgReg2IN_405, F(4)=>ImgReg2IN_404, F(3)=>
      ImgReg2IN_403, F(2)=>ImgReg2IN_402, F(1)=>ImgReg2IN_401, F(0)=>
      ImgReg2IN_400);
   loop3_25_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_431_EXMPLR, D(14)=>OutputImg3_430_EXMPLR, D(13)=>
      OutputImg3_429_EXMPLR, D(12)=>OutputImg3_428_EXMPLR, D(11)=>
      OutputImg3_427_EXMPLR, D(10)=>OutputImg3_426_EXMPLR, D(9)=>
      OutputImg3_425_EXMPLR, D(8)=>OutputImg3_424_EXMPLR, D(7)=>
      OutputImg3_423_EXMPLR, D(6)=>OutputImg3_422_EXMPLR, D(5)=>
      OutputImg3_421_EXMPLR, D(4)=>OutputImg3_420_EXMPLR, D(3)=>
      OutputImg3_419_EXMPLR, D(2)=>OutputImg3_418_EXMPLR, D(1)=>
      OutputImg3_417_EXMPLR, D(0)=>OutputImg3_416_EXMPLR, EN=>nx23708, F(15)
      =>ImgReg3IN_415, F(14)=>ImgReg3IN_414, F(13)=>ImgReg3IN_413, F(12)=>
      ImgReg3IN_412, F(11)=>ImgReg3IN_411, F(10)=>ImgReg3IN_410, F(9)=>
      ImgReg3IN_409, F(8)=>ImgReg3IN_408, F(7)=>ImgReg3IN_407, F(6)=>
      ImgReg3IN_406, F(5)=>ImgReg3IN_405, F(4)=>ImgReg3IN_404, F(3)=>
      ImgReg3IN_403, F(2)=>ImgReg3IN_402, F(1)=>ImgReg3IN_401, F(0)=>
      ImgReg3IN_400);
   loop3_25_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_431_EXMPLR, D(14)=>OutputImg4_430_EXMPLR, D(13)=>
      OutputImg4_429_EXMPLR, D(12)=>OutputImg4_428_EXMPLR, D(11)=>
      OutputImg4_427_EXMPLR, D(10)=>OutputImg4_426_EXMPLR, D(9)=>
      OutputImg4_425_EXMPLR, D(8)=>OutputImg4_424_EXMPLR, D(7)=>
      OutputImg4_423_EXMPLR, D(6)=>OutputImg4_422_EXMPLR, D(5)=>
      OutputImg4_421_EXMPLR, D(4)=>OutputImg4_420_EXMPLR, D(3)=>
      OutputImg4_419_EXMPLR, D(2)=>OutputImg4_418_EXMPLR, D(1)=>
      OutputImg4_417_EXMPLR, D(0)=>OutputImg4_416_EXMPLR, EN=>nx23710, F(15)
      =>ImgReg4IN_415, F(14)=>ImgReg4IN_414, F(13)=>ImgReg4IN_413, F(12)=>
      ImgReg4IN_412, F(11)=>ImgReg4IN_411, F(10)=>ImgReg4IN_410, F(9)=>
      ImgReg4IN_409, F(8)=>ImgReg4IN_408, F(7)=>ImgReg4IN_407, F(6)=>
      ImgReg4IN_406, F(5)=>ImgReg4IN_405, F(4)=>ImgReg4IN_404, F(3)=>
      ImgReg4IN_403, F(2)=>ImgReg4IN_402, F(1)=>ImgReg4IN_401, F(0)=>
      ImgReg4IN_400);
   loop3_25_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_431_EXMPLR, D(14)=>OutputImg5_430_EXMPLR, D(13)=>
      OutputImg5_429_EXMPLR, D(12)=>OutputImg5_428_EXMPLR, D(11)=>
      OutputImg5_427_EXMPLR, D(10)=>OutputImg5_426_EXMPLR, D(9)=>
      OutputImg5_425_EXMPLR, D(8)=>OutputImg5_424_EXMPLR, D(7)=>
      OutputImg5_423_EXMPLR, D(6)=>OutputImg5_422_EXMPLR, D(5)=>
      OutputImg5_421_EXMPLR, D(4)=>OutputImg5_420_EXMPLR, D(3)=>
      OutputImg5_419_EXMPLR, D(2)=>OutputImg5_418_EXMPLR, D(1)=>
      OutputImg5_417_EXMPLR, D(0)=>OutputImg5_416_EXMPLR, EN=>nx23710, F(15)
      =>ImgReg5IN_415, F(14)=>ImgReg5IN_414, F(13)=>ImgReg5IN_413, F(12)=>
      ImgReg5IN_412, F(11)=>ImgReg5IN_411, F(10)=>ImgReg5IN_410, F(9)=>
      ImgReg5IN_409, F(8)=>ImgReg5IN_408, F(7)=>ImgReg5IN_407, F(6)=>
      ImgReg5IN_406, F(5)=>ImgReg5IN_405, F(4)=>ImgReg5IN_404, F(3)=>
      ImgReg5IN_403, F(2)=>ImgReg5IN_402, F(1)=>ImgReg5IN_401, F(0)=>
      ImgReg5IN_400);
   loop3_25_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(415), 
      D(14)=>DATA(414), D(13)=>DATA(413), D(12)=>DATA(412), D(11)=>DATA(411), 
      D(10)=>DATA(410), D(9)=>DATA(409), D(8)=>DATA(408), D(7)=>DATA(407), 
      D(6)=>DATA(406), D(5)=>DATA(405), D(4)=>DATA(404), D(3)=>DATA(403), 
      D(2)=>DATA(402), D(1)=>DATA(401), D(0)=>DATA(400), EN=>nx23660, F(15)
      =>ImgReg0IN_415, F(14)=>ImgReg0IN_414, F(13)=>ImgReg0IN_413, F(12)=>
      ImgReg0IN_412, F(11)=>ImgReg0IN_411, F(10)=>ImgReg0IN_410, F(9)=>
      ImgReg0IN_409, F(8)=>ImgReg0IN_408, F(7)=>ImgReg0IN_407, F(6)=>
      ImgReg0IN_406, F(5)=>ImgReg0IN_405, F(4)=>ImgReg0IN_404, F(3)=>
      ImgReg0IN_403, F(2)=>ImgReg0IN_402, F(1)=>ImgReg0IN_401, F(0)=>
      ImgReg0IN_400);
   loop3_25_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(415), 
      D(14)=>DATA(414), D(13)=>DATA(413), D(12)=>DATA(412), D(11)=>DATA(411), 
      D(10)=>DATA(410), D(9)=>DATA(409), D(8)=>DATA(408), D(7)=>DATA(407), 
      D(6)=>DATA(406), D(5)=>DATA(405), D(4)=>DATA(404), D(3)=>DATA(403), 
      D(2)=>DATA(402), D(1)=>DATA(401), D(0)=>DATA(400), EN=>nx23648, F(15)
      =>ImgReg1IN_415, F(14)=>ImgReg1IN_414, F(13)=>ImgReg1IN_413, F(12)=>
      ImgReg1IN_412, F(11)=>ImgReg1IN_411, F(10)=>ImgReg1IN_410, F(9)=>
      ImgReg1IN_409, F(8)=>ImgReg1IN_408, F(7)=>ImgReg1IN_407, F(6)=>
      ImgReg1IN_406, F(5)=>ImgReg1IN_405, F(4)=>ImgReg1IN_404, F(3)=>
      ImgReg1IN_403, F(2)=>ImgReg1IN_402, F(1)=>ImgReg1IN_401, F(0)=>
      ImgReg1IN_400);
   loop3_25_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(415), 
      D(14)=>DATA(414), D(13)=>DATA(413), D(12)=>DATA(412), D(11)=>DATA(411), 
      D(10)=>DATA(410), D(9)=>DATA(409), D(8)=>DATA(408), D(7)=>DATA(407), 
      D(6)=>DATA(406), D(5)=>DATA(405), D(4)=>DATA(404), D(3)=>DATA(403), 
      D(2)=>DATA(402), D(1)=>DATA(401), D(0)=>DATA(400), EN=>nx23636, F(15)
      =>ImgReg2IN_415, F(14)=>ImgReg2IN_414, F(13)=>ImgReg2IN_413, F(12)=>
      ImgReg2IN_412, F(11)=>ImgReg2IN_411, F(10)=>ImgReg2IN_410, F(9)=>
      ImgReg2IN_409, F(8)=>ImgReg2IN_408, F(7)=>ImgReg2IN_407, F(6)=>
      ImgReg2IN_406, F(5)=>ImgReg2IN_405, F(4)=>ImgReg2IN_404, F(3)=>
      ImgReg2IN_403, F(2)=>ImgReg2IN_402, F(1)=>ImgReg2IN_401, F(0)=>
      ImgReg2IN_400);
   loop3_25_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(415), 
      D(14)=>DATA(414), D(13)=>DATA(413), D(12)=>DATA(412), D(11)=>DATA(411), 
      D(10)=>DATA(410), D(9)=>DATA(409), D(8)=>DATA(408), D(7)=>DATA(407), 
      D(6)=>DATA(406), D(5)=>DATA(405), D(4)=>DATA(404), D(3)=>DATA(403), 
      D(2)=>DATA(402), D(1)=>DATA(401), D(0)=>DATA(400), EN=>nx23624, F(15)
      =>ImgReg3IN_415, F(14)=>ImgReg3IN_414, F(13)=>ImgReg3IN_413, F(12)=>
      ImgReg3IN_412, F(11)=>ImgReg3IN_411, F(10)=>ImgReg3IN_410, F(9)=>
      ImgReg3IN_409, F(8)=>ImgReg3IN_408, F(7)=>ImgReg3IN_407, F(6)=>
      ImgReg3IN_406, F(5)=>ImgReg3IN_405, F(4)=>ImgReg3IN_404, F(3)=>
      ImgReg3IN_403, F(2)=>ImgReg3IN_402, F(1)=>ImgReg3IN_401, F(0)=>
      ImgReg3IN_400);
   loop3_25_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(415), 
      D(14)=>DATA(414), D(13)=>DATA(413), D(12)=>DATA(412), D(11)=>DATA(411), 
      D(10)=>DATA(410), D(9)=>DATA(409), D(8)=>DATA(408), D(7)=>DATA(407), 
      D(6)=>DATA(406), D(5)=>DATA(405), D(4)=>DATA(404), D(3)=>DATA(403), 
      D(2)=>DATA(402), D(1)=>DATA(401), D(0)=>DATA(400), EN=>nx23612, F(15)
      =>ImgReg4IN_415, F(14)=>ImgReg4IN_414, F(13)=>ImgReg4IN_413, F(12)=>
      ImgReg4IN_412, F(11)=>ImgReg4IN_411, F(10)=>ImgReg4IN_410, F(9)=>
      ImgReg4IN_409, F(8)=>ImgReg4IN_408, F(7)=>ImgReg4IN_407, F(6)=>
      ImgReg4IN_406, F(5)=>ImgReg4IN_405, F(4)=>ImgReg4IN_404, F(3)=>
      ImgReg4IN_403, F(2)=>ImgReg4IN_402, F(1)=>ImgReg4IN_401, F(0)=>
      ImgReg4IN_400);
   loop3_25_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(415), 
      D(14)=>DATA(414), D(13)=>DATA(413), D(12)=>DATA(412), D(11)=>DATA(411), 
      D(10)=>DATA(410), D(9)=>DATA(409), D(8)=>DATA(408), D(7)=>DATA(407), 
      D(6)=>DATA(406), D(5)=>DATA(405), D(4)=>DATA(404), D(3)=>DATA(403), 
      D(2)=>DATA(402), D(1)=>DATA(401), D(0)=>DATA(400), EN=>nx23600, F(15)
      =>ImgReg5IN_415, F(14)=>ImgReg5IN_414, F(13)=>ImgReg5IN_413, F(12)=>
      ImgReg5IN_412, F(11)=>ImgReg5IN_411, F(10)=>ImgReg5IN_410, F(9)=>
      ImgReg5IN_409, F(8)=>ImgReg5IN_408, F(7)=>ImgReg5IN_407, F(6)=>
      ImgReg5IN_406, F(5)=>ImgReg5IN_405, F(4)=>ImgReg5IN_404, F(3)=>
      ImgReg5IN_403, F(2)=>ImgReg5IN_402, F(1)=>ImgReg5IN_401, F(0)=>
      ImgReg5IN_400);
   loop3_25_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_415_EXMPLR, D(14)=>OutputImg1_414_EXMPLR, D(13)=>
      OutputImg1_413_EXMPLR, D(12)=>OutputImg1_412_EXMPLR, D(11)=>
      OutputImg1_411_EXMPLR, D(10)=>OutputImg1_410_EXMPLR, D(9)=>
      OutputImg1_409_EXMPLR, D(8)=>OutputImg1_408_EXMPLR, D(7)=>
      OutputImg1_407_EXMPLR, D(6)=>OutputImg1_406_EXMPLR, D(5)=>
      OutputImg1_405_EXMPLR, D(4)=>OutputImg1_404_EXMPLR, D(3)=>
      OutputImg1_403_EXMPLR, D(2)=>OutputImg1_402_EXMPLR, D(1)=>
      OutputImg1_401_EXMPLR, D(0)=>OutputImg1_400_EXMPLR, EN=>nx23820, F(15)
      =>ImgReg0IN_415, F(14)=>ImgReg0IN_414, F(13)=>ImgReg0IN_413, F(12)=>
      ImgReg0IN_412, F(11)=>ImgReg0IN_411, F(10)=>ImgReg0IN_410, F(9)=>
      ImgReg0IN_409, F(8)=>ImgReg0IN_408, F(7)=>ImgReg0IN_407, F(6)=>
      ImgReg0IN_406, F(5)=>ImgReg0IN_405, F(4)=>ImgReg0IN_404, F(3)=>
      ImgReg0IN_403, F(2)=>ImgReg0IN_402, F(1)=>ImgReg0IN_401, F(0)=>
      ImgReg0IN_400);
   loop3_25_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_415_EXMPLR, D(14)=>OutputImg2_414_EXMPLR, D(13)=>
      OutputImg2_413_EXMPLR, D(12)=>OutputImg2_412_EXMPLR, D(11)=>
      OutputImg2_411_EXMPLR, D(10)=>OutputImg2_410_EXMPLR, D(9)=>
      OutputImg2_409_EXMPLR, D(8)=>OutputImg2_408_EXMPLR, D(7)=>
      OutputImg2_407_EXMPLR, D(6)=>OutputImg2_406_EXMPLR, D(5)=>
      OutputImg2_405_EXMPLR, D(4)=>OutputImg2_404_EXMPLR, D(3)=>
      OutputImg2_403_EXMPLR, D(2)=>OutputImg2_402_EXMPLR, D(1)=>
      OutputImg2_401_EXMPLR, D(0)=>OutputImg2_400_EXMPLR, EN=>nx23822, F(15)
      =>ImgReg1IN_415, F(14)=>ImgReg1IN_414, F(13)=>ImgReg1IN_413, F(12)=>
      ImgReg1IN_412, F(11)=>ImgReg1IN_411, F(10)=>ImgReg1IN_410, F(9)=>
      ImgReg1IN_409, F(8)=>ImgReg1IN_408, F(7)=>ImgReg1IN_407, F(6)=>
      ImgReg1IN_406, F(5)=>ImgReg1IN_405, F(4)=>ImgReg1IN_404, F(3)=>
      ImgReg1IN_403, F(2)=>ImgReg1IN_402, F(1)=>ImgReg1IN_401, F(0)=>
      ImgReg1IN_400);
   loop3_25_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_415_EXMPLR, D(14)=>OutputImg3_414_EXMPLR, D(13)=>
      OutputImg3_413_EXMPLR, D(12)=>OutputImg3_412_EXMPLR, D(11)=>
      OutputImg3_411_EXMPLR, D(10)=>OutputImg3_410_EXMPLR, D(9)=>
      OutputImg3_409_EXMPLR, D(8)=>OutputImg3_408_EXMPLR, D(7)=>
      OutputImg3_407_EXMPLR, D(6)=>OutputImg3_406_EXMPLR, D(5)=>
      OutputImg3_405_EXMPLR, D(4)=>OutputImg3_404_EXMPLR, D(3)=>
      OutputImg3_403_EXMPLR, D(2)=>OutputImg3_402_EXMPLR, D(1)=>
      OutputImg3_401_EXMPLR, D(0)=>OutputImg3_400_EXMPLR, EN=>nx23822, F(15)
      =>ImgReg2IN_415, F(14)=>ImgReg2IN_414, F(13)=>ImgReg2IN_413, F(12)=>
      ImgReg2IN_412, F(11)=>ImgReg2IN_411, F(10)=>ImgReg2IN_410, F(9)=>
      ImgReg2IN_409, F(8)=>ImgReg2IN_408, F(7)=>ImgReg2IN_407, F(6)=>
      ImgReg2IN_406, F(5)=>ImgReg2IN_405, F(4)=>ImgReg2IN_404, F(3)=>
      ImgReg2IN_403, F(2)=>ImgReg2IN_402, F(1)=>ImgReg2IN_401, F(0)=>
      ImgReg2IN_400);
   loop3_25_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_415_EXMPLR, D(14)=>OutputImg4_414_EXMPLR, D(13)=>
      OutputImg4_413_EXMPLR, D(12)=>OutputImg4_412_EXMPLR, D(11)=>
      OutputImg4_411_EXMPLR, D(10)=>OutputImg4_410_EXMPLR, D(9)=>
      OutputImg4_409_EXMPLR, D(8)=>OutputImg4_408_EXMPLR, D(7)=>
      OutputImg4_407_EXMPLR, D(6)=>OutputImg4_406_EXMPLR, D(5)=>
      OutputImg4_405_EXMPLR, D(4)=>OutputImg4_404_EXMPLR, D(3)=>
      OutputImg4_403_EXMPLR, D(2)=>OutputImg4_402_EXMPLR, D(1)=>
      OutputImg4_401_EXMPLR, D(0)=>OutputImg4_400_EXMPLR, EN=>nx23822, F(15)
      =>ImgReg3IN_415, F(14)=>ImgReg3IN_414, F(13)=>ImgReg3IN_413, F(12)=>
      ImgReg3IN_412, F(11)=>ImgReg3IN_411, F(10)=>ImgReg3IN_410, F(9)=>
      ImgReg3IN_409, F(8)=>ImgReg3IN_408, F(7)=>ImgReg3IN_407, F(6)=>
      ImgReg3IN_406, F(5)=>ImgReg3IN_405, F(4)=>ImgReg3IN_404, F(3)=>
      ImgReg3IN_403, F(2)=>ImgReg3IN_402, F(1)=>ImgReg3IN_401, F(0)=>
      ImgReg3IN_400);
   loop3_25_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_415_EXMPLR, D(14)=>OutputImg5_414_EXMPLR, D(13)=>
      OutputImg5_413_EXMPLR, D(12)=>OutputImg5_412_EXMPLR, D(11)=>
      OutputImg5_411_EXMPLR, D(10)=>OutputImg5_410_EXMPLR, D(9)=>
      OutputImg5_409_EXMPLR, D(8)=>OutputImg5_408_EXMPLR, D(7)=>
      OutputImg5_407_EXMPLR, D(6)=>OutputImg5_406_EXMPLR, D(5)=>
      OutputImg5_405_EXMPLR, D(4)=>OutputImg5_404_EXMPLR, D(3)=>
      OutputImg5_403_EXMPLR, D(2)=>OutputImg5_402_EXMPLR, D(1)=>
      OutputImg5_401_EXMPLR, D(0)=>OutputImg5_400_EXMPLR, EN=>nx23822, F(15)
      =>ImgReg4IN_415, F(14)=>ImgReg4IN_414, F(13)=>ImgReg4IN_413, F(12)=>
      ImgReg4IN_412, F(11)=>ImgReg4IN_411, F(10)=>ImgReg4IN_410, F(9)=>
      ImgReg4IN_409, F(8)=>ImgReg4IN_408, F(7)=>ImgReg4IN_407, F(6)=>
      ImgReg4IN_406, F(5)=>ImgReg4IN_405, F(4)=>ImgReg4IN_404, F(3)=>
      ImgReg4IN_403, F(2)=>ImgReg4IN_402, F(1)=>ImgReg4IN_401, F(0)=>
      ImgReg4IN_400);
   loop3_25_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_415, D(14)=>
      ImgReg0IN_414, D(13)=>ImgReg0IN_413, D(12)=>ImgReg0IN_412, D(11)=>
      ImgReg0IN_411, D(10)=>ImgReg0IN_410, D(9)=>ImgReg0IN_409, D(8)=>
      ImgReg0IN_408, D(7)=>ImgReg0IN_407, D(6)=>ImgReg0IN_406, D(5)=>
      ImgReg0IN_405, D(4)=>ImgReg0IN_404, D(3)=>ImgReg0IN_403, D(2)=>
      ImgReg0IN_402, D(1)=>ImgReg0IN_401, D(0)=>ImgReg0IN_400, CLK=>nx23978, 
      RST=>RST, EN=>nx23724, Q(15)=>OutputImg0_415_EXMPLR, Q(14)=>
      OutputImg0_414_EXMPLR, Q(13)=>OutputImg0_413_EXMPLR, Q(12)=>
      OutputImg0_412_EXMPLR, Q(11)=>OutputImg0_411_EXMPLR, Q(10)=>
      OutputImg0_410_EXMPLR, Q(9)=>OutputImg0_409_EXMPLR, Q(8)=>
      OutputImg0_408_EXMPLR, Q(7)=>OutputImg0_407_EXMPLR, Q(6)=>
      OutputImg0_406_EXMPLR, Q(5)=>OutputImg0_405_EXMPLR, Q(4)=>
      OutputImg0_404_EXMPLR, Q(3)=>OutputImg0_403_EXMPLR, Q(2)=>
      OutputImg0_402_EXMPLR, Q(1)=>OutputImg0_401_EXMPLR, Q(0)=>
      OutputImg0_400_EXMPLR);
   loop3_25_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_415, D(14)=>
      ImgReg1IN_414, D(13)=>ImgReg1IN_413, D(12)=>ImgReg1IN_412, D(11)=>
      ImgReg1IN_411, D(10)=>ImgReg1IN_410, D(9)=>ImgReg1IN_409, D(8)=>
      ImgReg1IN_408, D(7)=>ImgReg1IN_407, D(6)=>ImgReg1IN_406, D(5)=>
      ImgReg1IN_405, D(4)=>ImgReg1IN_404, D(3)=>ImgReg1IN_403, D(2)=>
      ImgReg1IN_402, D(1)=>ImgReg1IN_401, D(0)=>ImgReg1IN_400, CLK=>nx23980, 
      RST=>RST, EN=>nx23734, Q(15)=>OutputImg1_415_EXMPLR, Q(14)=>
      OutputImg1_414_EXMPLR, Q(13)=>OutputImg1_413_EXMPLR, Q(12)=>
      OutputImg1_412_EXMPLR, Q(11)=>OutputImg1_411_EXMPLR, Q(10)=>
      OutputImg1_410_EXMPLR, Q(9)=>OutputImg1_409_EXMPLR, Q(8)=>
      OutputImg1_408_EXMPLR, Q(7)=>OutputImg1_407_EXMPLR, Q(6)=>
      OutputImg1_406_EXMPLR, Q(5)=>OutputImg1_405_EXMPLR, Q(4)=>
      OutputImg1_404_EXMPLR, Q(3)=>OutputImg1_403_EXMPLR, Q(2)=>
      OutputImg1_402_EXMPLR, Q(1)=>OutputImg1_401_EXMPLR, Q(0)=>
      OutputImg1_400_EXMPLR);
   loop3_25_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_415, D(14)=>
      ImgReg2IN_414, D(13)=>ImgReg2IN_413, D(12)=>ImgReg2IN_412, D(11)=>
      ImgReg2IN_411, D(10)=>ImgReg2IN_410, D(9)=>ImgReg2IN_409, D(8)=>
      ImgReg2IN_408, D(7)=>ImgReg2IN_407, D(6)=>ImgReg2IN_406, D(5)=>
      ImgReg2IN_405, D(4)=>ImgReg2IN_404, D(3)=>ImgReg2IN_403, D(2)=>
      ImgReg2IN_402, D(1)=>ImgReg2IN_401, D(0)=>ImgReg2IN_400, CLK=>nx23980, 
      RST=>RST, EN=>nx23744, Q(15)=>OutputImg2_415_EXMPLR, Q(14)=>
      OutputImg2_414_EXMPLR, Q(13)=>OutputImg2_413_EXMPLR, Q(12)=>
      OutputImg2_412_EXMPLR, Q(11)=>OutputImg2_411_EXMPLR, Q(10)=>
      OutputImg2_410_EXMPLR, Q(9)=>OutputImg2_409_EXMPLR, Q(8)=>
      OutputImg2_408_EXMPLR, Q(7)=>OutputImg2_407_EXMPLR, Q(6)=>
      OutputImg2_406_EXMPLR, Q(5)=>OutputImg2_405_EXMPLR, Q(4)=>
      OutputImg2_404_EXMPLR, Q(3)=>OutputImg2_403_EXMPLR, Q(2)=>
      OutputImg2_402_EXMPLR, Q(1)=>OutputImg2_401_EXMPLR, Q(0)=>
      OutputImg2_400_EXMPLR);
   loop3_25_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_415, D(14)=>
      ImgReg3IN_414, D(13)=>ImgReg3IN_413, D(12)=>ImgReg3IN_412, D(11)=>
      ImgReg3IN_411, D(10)=>ImgReg3IN_410, D(9)=>ImgReg3IN_409, D(8)=>
      ImgReg3IN_408, D(7)=>ImgReg3IN_407, D(6)=>ImgReg3IN_406, D(5)=>
      ImgReg3IN_405, D(4)=>ImgReg3IN_404, D(3)=>ImgReg3IN_403, D(2)=>
      ImgReg3IN_402, D(1)=>ImgReg3IN_401, D(0)=>ImgReg3IN_400, CLK=>nx23982, 
      RST=>RST, EN=>nx23754, Q(15)=>OutputImg3_415_EXMPLR, Q(14)=>
      OutputImg3_414_EXMPLR, Q(13)=>OutputImg3_413_EXMPLR, Q(12)=>
      OutputImg3_412_EXMPLR, Q(11)=>OutputImg3_411_EXMPLR, Q(10)=>
      OutputImg3_410_EXMPLR, Q(9)=>OutputImg3_409_EXMPLR, Q(8)=>
      OutputImg3_408_EXMPLR, Q(7)=>OutputImg3_407_EXMPLR, Q(6)=>
      OutputImg3_406_EXMPLR, Q(5)=>OutputImg3_405_EXMPLR, Q(4)=>
      OutputImg3_404_EXMPLR, Q(3)=>OutputImg3_403_EXMPLR, Q(2)=>
      OutputImg3_402_EXMPLR, Q(1)=>OutputImg3_401_EXMPLR, Q(0)=>
      OutputImg3_400_EXMPLR);
   loop3_25_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_415, D(14)=>
      ImgReg4IN_414, D(13)=>ImgReg4IN_413, D(12)=>ImgReg4IN_412, D(11)=>
      ImgReg4IN_411, D(10)=>ImgReg4IN_410, D(9)=>ImgReg4IN_409, D(8)=>
      ImgReg4IN_408, D(7)=>ImgReg4IN_407, D(6)=>ImgReg4IN_406, D(5)=>
      ImgReg4IN_405, D(4)=>ImgReg4IN_404, D(3)=>ImgReg4IN_403, D(2)=>
      ImgReg4IN_402, D(1)=>ImgReg4IN_401, D(0)=>ImgReg4IN_400, CLK=>nx23982, 
      RST=>RST, EN=>nx23764, Q(15)=>OutputImg4_415_EXMPLR, Q(14)=>
      OutputImg4_414_EXMPLR, Q(13)=>OutputImg4_413_EXMPLR, Q(12)=>
      OutputImg4_412_EXMPLR, Q(11)=>OutputImg4_411_EXMPLR, Q(10)=>
      OutputImg4_410_EXMPLR, Q(9)=>OutputImg4_409_EXMPLR, Q(8)=>
      OutputImg4_408_EXMPLR, Q(7)=>OutputImg4_407_EXMPLR, Q(6)=>
      OutputImg4_406_EXMPLR, Q(5)=>OutputImg4_405_EXMPLR, Q(4)=>
      OutputImg4_404_EXMPLR, Q(3)=>OutputImg4_403_EXMPLR, Q(2)=>
      OutputImg4_402_EXMPLR, Q(1)=>OutputImg4_401_EXMPLR, Q(0)=>
      OutputImg4_400_EXMPLR);
   loop3_25_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_415, D(14)=>
      ImgReg5IN_414, D(13)=>ImgReg5IN_413, D(12)=>ImgReg5IN_412, D(11)=>
      ImgReg5IN_411, D(10)=>ImgReg5IN_410, D(9)=>ImgReg5IN_409, D(8)=>
      ImgReg5IN_408, D(7)=>ImgReg5IN_407, D(6)=>ImgReg5IN_406, D(5)=>
      ImgReg5IN_405, D(4)=>ImgReg5IN_404, D(3)=>ImgReg5IN_403, D(2)=>
      ImgReg5IN_402, D(1)=>ImgReg5IN_401, D(0)=>ImgReg5IN_400, CLK=>nx23984, 
      RST=>RST, EN=>nx23774, Q(15)=>OutputImg5_415_EXMPLR, Q(14)=>
      OutputImg5_414_EXMPLR, Q(13)=>OutputImg5_413_EXMPLR, Q(12)=>
      OutputImg5_412_EXMPLR, Q(11)=>OutputImg5_411_EXMPLR, Q(10)=>
      OutputImg5_410_EXMPLR, Q(9)=>OutputImg5_409_EXMPLR, Q(8)=>
      OutputImg5_408_EXMPLR, Q(7)=>OutputImg5_407_EXMPLR, Q(6)=>
      OutputImg5_406_EXMPLR, Q(5)=>OutputImg5_405_EXMPLR, Q(4)=>
      OutputImg5_404_EXMPLR, Q(3)=>OutputImg5_403_EXMPLR, Q(2)=>
      OutputImg5_402_EXMPLR, Q(1)=>OutputImg5_401_EXMPLR, Q(0)=>
      OutputImg5_400_EXMPLR);
   loop3_26_TriState0L : triStateBuffer_16 port map ( D(15)=>
      OutputImg0_447_EXMPLR, D(14)=>OutputImg0_446_EXMPLR, D(13)=>
      OutputImg0_445_EXMPLR, D(12)=>OutputImg0_444_EXMPLR, D(11)=>
      OutputImg0_443_EXMPLR, D(10)=>OutputImg0_442_EXMPLR, D(9)=>
      OutputImg0_441_EXMPLR, D(8)=>OutputImg0_440_EXMPLR, D(7)=>
      OutputImg0_439_EXMPLR, D(6)=>OutputImg0_438_EXMPLR, D(5)=>
      OutputImg0_437_EXMPLR, D(4)=>OutputImg0_436_EXMPLR, D(3)=>
      OutputImg0_435_EXMPLR, D(2)=>OutputImg0_434_EXMPLR, D(1)=>
      OutputImg0_433_EXMPLR, D(0)=>OutputImg0_432_EXMPLR, EN=>nx23710, F(15)
      =>ImgReg0IN_431, F(14)=>ImgReg0IN_430, F(13)=>ImgReg0IN_429, F(12)=>
      ImgReg0IN_428, F(11)=>ImgReg0IN_427, F(10)=>ImgReg0IN_426, F(9)=>
      ImgReg0IN_425, F(8)=>ImgReg0IN_424, F(7)=>ImgReg0IN_423, F(6)=>
      ImgReg0IN_422, F(5)=>ImgReg0IN_421, F(4)=>ImgReg0IN_420, F(3)=>
      ImgReg0IN_419, F(2)=>ImgReg0IN_418, F(1)=>ImgReg0IN_417, F(0)=>
      ImgReg0IN_416);
   loop3_26_TriState1L : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_447_EXMPLR, D(14)=>OutputImg1_446_EXMPLR, D(13)=>
      OutputImg1_445_EXMPLR, D(12)=>OutputImg1_444_EXMPLR, D(11)=>
      OutputImg1_443_EXMPLR, D(10)=>OutputImg1_442_EXMPLR, D(9)=>
      OutputImg1_441_EXMPLR, D(8)=>OutputImg1_440_EXMPLR, D(7)=>
      OutputImg1_439_EXMPLR, D(6)=>OutputImg1_438_EXMPLR, D(5)=>
      OutputImg1_437_EXMPLR, D(4)=>OutputImg1_436_EXMPLR, D(3)=>
      OutputImg1_435_EXMPLR, D(2)=>OutputImg1_434_EXMPLR, D(1)=>
      OutputImg1_433_EXMPLR, D(0)=>OutputImg1_432_EXMPLR, EN=>nx23710, F(15)
      =>ImgReg1IN_431, F(14)=>ImgReg1IN_430, F(13)=>ImgReg1IN_429, F(12)=>
      ImgReg1IN_428, F(11)=>ImgReg1IN_427, F(10)=>ImgReg1IN_426, F(9)=>
      ImgReg1IN_425, F(8)=>ImgReg1IN_424, F(7)=>ImgReg1IN_423, F(6)=>
      ImgReg1IN_422, F(5)=>ImgReg1IN_421, F(4)=>ImgReg1IN_420, F(3)=>
      ImgReg1IN_419, F(2)=>ImgReg1IN_418, F(1)=>ImgReg1IN_417, F(0)=>
      ImgReg1IN_416);
   loop3_26_TriState2L : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_447_EXMPLR, D(14)=>OutputImg2_446_EXMPLR, D(13)=>
      OutputImg2_445_EXMPLR, D(12)=>OutputImg2_444_EXMPLR, D(11)=>
      OutputImg2_443_EXMPLR, D(10)=>OutputImg2_442_EXMPLR, D(9)=>
      OutputImg2_441_EXMPLR, D(8)=>OutputImg2_440_EXMPLR, D(7)=>
      OutputImg2_439_EXMPLR, D(6)=>OutputImg2_438_EXMPLR, D(5)=>
      OutputImg2_437_EXMPLR, D(4)=>OutputImg2_436_EXMPLR, D(3)=>
      OutputImg2_435_EXMPLR, D(2)=>OutputImg2_434_EXMPLR, D(1)=>
      OutputImg2_433_EXMPLR, D(0)=>OutputImg2_432_EXMPLR, EN=>nx23710, F(15)
      =>ImgReg2IN_431, F(14)=>ImgReg2IN_430, F(13)=>ImgReg2IN_429, F(12)=>
      ImgReg2IN_428, F(11)=>ImgReg2IN_427, F(10)=>ImgReg2IN_426, F(9)=>
      ImgReg2IN_425, F(8)=>ImgReg2IN_424, F(7)=>ImgReg2IN_423, F(6)=>
      ImgReg2IN_422, F(5)=>ImgReg2IN_421, F(4)=>ImgReg2IN_420, F(3)=>
      ImgReg2IN_419, F(2)=>ImgReg2IN_418, F(1)=>ImgReg2IN_417, F(0)=>
      ImgReg2IN_416);
   loop3_26_TriState3L : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_447_EXMPLR, D(14)=>OutputImg3_446_EXMPLR, D(13)=>
      OutputImg3_445_EXMPLR, D(12)=>OutputImg3_444_EXMPLR, D(11)=>
      OutputImg3_443_EXMPLR, D(10)=>OutputImg3_442_EXMPLR, D(9)=>
      OutputImg3_441_EXMPLR, D(8)=>OutputImg3_440_EXMPLR, D(7)=>
      OutputImg3_439_EXMPLR, D(6)=>OutputImg3_438_EXMPLR, D(5)=>
      OutputImg3_437_EXMPLR, D(4)=>OutputImg3_436_EXMPLR, D(3)=>
      OutputImg3_435_EXMPLR, D(2)=>OutputImg3_434_EXMPLR, D(1)=>
      OutputImg3_433_EXMPLR, D(0)=>OutputImg3_432_EXMPLR, EN=>nx23710, F(15)
      =>ImgReg3IN_431, F(14)=>ImgReg3IN_430, F(13)=>ImgReg3IN_429, F(12)=>
      ImgReg3IN_428, F(11)=>ImgReg3IN_427, F(10)=>ImgReg3IN_426, F(9)=>
      ImgReg3IN_425, F(8)=>ImgReg3IN_424, F(7)=>ImgReg3IN_423, F(6)=>
      ImgReg3IN_422, F(5)=>ImgReg3IN_421, F(4)=>ImgReg3IN_420, F(3)=>
      ImgReg3IN_419, F(2)=>ImgReg3IN_418, F(1)=>ImgReg3IN_417, F(0)=>
      ImgReg3IN_416);
   loop3_26_TriState4L : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_447_EXMPLR, D(14)=>OutputImg4_446_EXMPLR, D(13)=>
      OutputImg4_445_EXMPLR, D(12)=>OutputImg4_444_EXMPLR, D(11)=>
      OutputImg4_443_EXMPLR, D(10)=>OutputImg4_442_EXMPLR, D(9)=>
      OutputImg4_441_EXMPLR, D(8)=>OutputImg4_440_EXMPLR, D(7)=>
      OutputImg4_439_EXMPLR, D(6)=>OutputImg4_438_EXMPLR, D(5)=>
      OutputImg4_437_EXMPLR, D(4)=>OutputImg4_436_EXMPLR, D(3)=>
      OutputImg4_435_EXMPLR, D(2)=>OutputImg4_434_EXMPLR, D(1)=>
      OutputImg4_433_EXMPLR, D(0)=>OutputImg4_432_EXMPLR, EN=>nx23710, F(15)
      =>ImgReg4IN_431, F(14)=>ImgReg4IN_430, F(13)=>ImgReg4IN_429, F(12)=>
      ImgReg4IN_428, F(11)=>ImgReg4IN_427, F(10)=>ImgReg4IN_426, F(9)=>
      ImgReg4IN_425, F(8)=>ImgReg4IN_424, F(7)=>ImgReg4IN_423, F(6)=>
      ImgReg4IN_422, F(5)=>ImgReg4IN_421, F(4)=>ImgReg4IN_420, F(3)=>
      ImgReg4IN_419, F(2)=>ImgReg4IN_418, F(1)=>ImgReg4IN_417, F(0)=>
      ImgReg4IN_416);
   loop3_26_TriState5L : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_447_EXMPLR, D(14)=>OutputImg5_446_EXMPLR, D(13)=>
      OutputImg5_445_EXMPLR, D(12)=>OutputImg5_444_EXMPLR, D(11)=>
      OutputImg5_443_EXMPLR, D(10)=>OutputImg5_442_EXMPLR, D(9)=>
      OutputImg5_441_EXMPLR, D(8)=>OutputImg5_440_EXMPLR, D(7)=>
      OutputImg5_439_EXMPLR, D(6)=>OutputImg5_438_EXMPLR, D(5)=>
      OutputImg5_437_EXMPLR, D(4)=>OutputImg5_436_EXMPLR, D(3)=>
      OutputImg5_435_EXMPLR, D(2)=>OutputImg5_434_EXMPLR, D(1)=>
      OutputImg5_433_EXMPLR, D(0)=>OutputImg5_432_EXMPLR, EN=>nx23712, F(15)
      =>ImgReg5IN_431, F(14)=>ImgReg5IN_430, F(13)=>ImgReg5IN_429, F(12)=>
      ImgReg5IN_428, F(11)=>ImgReg5IN_427, F(10)=>ImgReg5IN_426, F(9)=>
      ImgReg5IN_425, F(8)=>ImgReg5IN_424, F(7)=>ImgReg5IN_423, F(6)=>
      ImgReg5IN_422, F(5)=>ImgReg5IN_421, F(4)=>ImgReg5IN_420, F(3)=>
      ImgReg5IN_419, F(2)=>ImgReg5IN_418, F(1)=>ImgReg5IN_417, F(0)=>
      ImgReg5IN_416);
   loop3_26_TriState0N : triStateBuffer_16 port map ( D(15)=>DATA(431), 
      D(14)=>DATA(430), D(13)=>DATA(429), D(12)=>DATA(428), D(11)=>DATA(427), 
      D(10)=>DATA(426), D(9)=>DATA(425), D(8)=>DATA(424), D(7)=>DATA(423), 
      D(6)=>DATA(422), D(5)=>DATA(421), D(4)=>DATA(420), D(3)=>DATA(419), 
      D(2)=>DATA(418), D(1)=>DATA(417), D(0)=>DATA(416), EN=>nx23660, F(15)
      =>ImgReg0IN_431, F(14)=>ImgReg0IN_430, F(13)=>ImgReg0IN_429, F(12)=>
      ImgReg0IN_428, F(11)=>ImgReg0IN_427, F(10)=>ImgReg0IN_426, F(9)=>
      ImgReg0IN_425, F(8)=>ImgReg0IN_424, F(7)=>ImgReg0IN_423, F(6)=>
      ImgReg0IN_422, F(5)=>ImgReg0IN_421, F(4)=>ImgReg0IN_420, F(3)=>
      ImgReg0IN_419, F(2)=>ImgReg0IN_418, F(1)=>ImgReg0IN_417, F(0)=>
      ImgReg0IN_416);
   loop3_26_TriState1N : triStateBuffer_16 port map ( D(15)=>DATA(431), 
      D(14)=>DATA(430), D(13)=>DATA(429), D(12)=>DATA(428), D(11)=>DATA(427), 
      D(10)=>DATA(426), D(9)=>DATA(425), D(8)=>DATA(424), D(7)=>DATA(423), 
      D(6)=>DATA(422), D(5)=>DATA(421), D(4)=>DATA(420), D(3)=>DATA(419), 
      D(2)=>DATA(418), D(1)=>DATA(417), D(0)=>DATA(416), EN=>nx23648, F(15)
      =>ImgReg1IN_431, F(14)=>ImgReg1IN_430, F(13)=>ImgReg1IN_429, F(12)=>
      ImgReg1IN_428, F(11)=>ImgReg1IN_427, F(10)=>ImgReg1IN_426, F(9)=>
      ImgReg1IN_425, F(8)=>ImgReg1IN_424, F(7)=>ImgReg1IN_423, F(6)=>
      ImgReg1IN_422, F(5)=>ImgReg1IN_421, F(4)=>ImgReg1IN_420, F(3)=>
      ImgReg1IN_419, F(2)=>ImgReg1IN_418, F(1)=>ImgReg1IN_417, F(0)=>
      ImgReg1IN_416);
   loop3_26_TriState2N : triStateBuffer_16 port map ( D(15)=>DATA(431), 
      D(14)=>DATA(430), D(13)=>DATA(429), D(12)=>DATA(428), D(11)=>DATA(427), 
      D(10)=>DATA(426), D(9)=>DATA(425), D(8)=>DATA(424), D(7)=>DATA(423), 
      D(6)=>DATA(422), D(5)=>DATA(421), D(4)=>DATA(420), D(3)=>DATA(419), 
      D(2)=>DATA(418), D(1)=>DATA(417), D(0)=>DATA(416), EN=>nx23636, F(15)
      =>ImgReg2IN_431, F(14)=>ImgReg2IN_430, F(13)=>ImgReg2IN_429, F(12)=>
      ImgReg2IN_428, F(11)=>ImgReg2IN_427, F(10)=>ImgReg2IN_426, F(9)=>
      ImgReg2IN_425, F(8)=>ImgReg2IN_424, F(7)=>ImgReg2IN_423, F(6)=>
      ImgReg2IN_422, F(5)=>ImgReg2IN_421, F(4)=>ImgReg2IN_420, F(3)=>
      ImgReg2IN_419, F(2)=>ImgReg2IN_418, F(1)=>ImgReg2IN_417, F(0)=>
      ImgReg2IN_416);
   loop3_26_TriState3N : triStateBuffer_16 port map ( D(15)=>DATA(431), 
      D(14)=>DATA(430), D(13)=>DATA(429), D(12)=>DATA(428), D(11)=>DATA(427), 
      D(10)=>DATA(426), D(9)=>DATA(425), D(8)=>DATA(424), D(7)=>DATA(423), 
      D(6)=>DATA(422), D(5)=>DATA(421), D(4)=>DATA(420), D(3)=>DATA(419), 
      D(2)=>DATA(418), D(1)=>DATA(417), D(0)=>DATA(416), EN=>nx23624, F(15)
      =>ImgReg3IN_431, F(14)=>ImgReg3IN_430, F(13)=>ImgReg3IN_429, F(12)=>
      ImgReg3IN_428, F(11)=>ImgReg3IN_427, F(10)=>ImgReg3IN_426, F(9)=>
      ImgReg3IN_425, F(8)=>ImgReg3IN_424, F(7)=>ImgReg3IN_423, F(6)=>
      ImgReg3IN_422, F(5)=>ImgReg3IN_421, F(4)=>ImgReg3IN_420, F(3)=>
      ImgReg3IN_419, F(2)=>ImgReg3IN_418, F(1)=>ImgReg3IN_417, F(0)=>
      ImgReg3IN_416);
   loop3_26_TriState4N : triStateBuffer_16 port map ( D(15)=>DATA(431), 
      D(14)=>DATA(430), D(13)=>DATA(429), D(12)=>DATA(428), D(11)=>DATA(427), 
      D(10)=>DATA(426), D(9)=>DATA(425), D(8)=>DATA(424), D(7)=>DATA(423), 
      D(6)=>DATA(422), D(5)=>DATA(421), D(4)=>DATA(420), D(3)=>DATA(419), 
      D(2)=>DATA(418), D(1)=>DATA(417), D(0)=>DATA(416), EN=>nx23612, F(15)
      =>ImgReg4IN_431, F(14)=>ImgReg4IN_430, F(13)=>ImgReg4IN_429, F(12)=>
      ImgReg4IN_428, F(11)=>ImgReg4IN_427, F(10)=>ImgReg4IN_426, F(9)=>
      ImgReg4IN_425, F(8)=>ImgReg4IN_424, F(7)=>ImgReg4IN_423, F(6)=>
      ImgReg4IN_422, F(5)=>ImgReg4IN_421, F(4)=>ImgReg4IN_420, F(3)=>
      ImgReg4IN_419, F(2)=>ImgReg4IN_418, F(1)=>ImgReg4IN_417, F(0)=>
      ImgReg4IN_416);
   loop3_26_TriState5N : triStateBuffer_16 port map ( D(15)=>DATA(431), 
      D(14)=>DATA(430), D(13)=>DATA(429), D(12)=>DATA(428), D(11)=>DATA(427), 
      D(10)=>DATA(426), D(9)=>DATA(425), D(8)=>DATA(424), D(7)=>DATA(423), 
      D(6)=>DATA(422), D(5)=>DATA(421), D(4)=>DATA(420), D(3)=>DATA(419), 
      D(2)=>DATA(418), D(1)=>DATA(417), D(0)=>DATA(416), EN=>nx23600, F(15)
      =>ImgReg5IN_431, F(14)=>ImgReg5IN_430, F(13)=>ImgReg5IN_429, F(12)=>
      ImgReg5IN_428, F(11)=>ImgReg5IN_427, F(10)=>ImgReg5IN_426, F(9)=>
      ImgReg5IN_425, F(8)=>ImgReg5IN_424, F(7)=>ImgReg5IN_423, F(6)=>
      ImgReg5IN_422, F(5)=>ImgReg5IN_421, F(4)=>ImgReg5IN_420, F(3)=>
      ImgReg5IN_419, F(2)=>ImgReg5IN_418, F(1)=>ImgReg5IN_417, F(0)=>
      ImgReg5IN_416);
   loop3_26_TriState0U : triStateBuffer_16 port map ( D(15)=>
      OutputImg1_431_EXMPLR, D(14)=>OutputImg1_430_EXMPLR, D(13)=>
      OutputImg1_429_EXMPLR, D(12)=>OutputImg1_428_EXMPLR, D(11)=>
      OutputImg1_427_EXMPLR, D(10)=>OutputImg1_426_EXMPLR, D(9)=>
      OutputImg1_425_EXMPLR, D(8)=>OutputImg1_424_EXMPLR, D(7)=>
      OutputImg1_423_EXMPLR, D(6)=>OutputImg1_422_EXMPLR, D(5)=>
      OutputImg1_421_EXMPLR, D(4)=>OutputImg1_420_EXMPLR, D(3)=>
      OutputImg1_419_EXMPLR, D(2)=>OutputImg1_418_EXMPLR, D(1)=>
      OutputImg1_417_EXMPLR, D(0)=>OutputImg1_416_EXMPLR, EN=>nx23822, F(15)
      =>ImgReg0IN_431, F(14)=>ImgReg0IN_430, F(13)=>ImgReg0IN_429, F(12)=>
      ImgReg0IN_428, F(11)=>ImgReg0IN_427, F(10)=>ImgReg0IN_426, F(9)=>
      ImgReg0IN_425, F(8)=>ImgReg0IN_424, F(7)=>ImgReg0IN_423, F(6)=>
      ImgReg0IN_422, F(5)=>ImgReg0IN_421, F(4)=>ImgReg0IN_420, F(3)=>
      ImgReg0IN_419, F(2)=>ImgReg0IN_418, F(1)=>ImgReg0IN_417, F(0)=>
      ImgReg0IN_416);
   loop3_26_TriState1U : triStateBuffer_16 port map ( D(15)=>
      OutputImg2_431_EXMPLR, D(14)=>OutputImg2_430_EXMPLR, D(13)=>
      OutputImg2_429_EXMPLR, D(12)=>OutputImg2_428_EXMPLR, D(11)=>
      OutputImg2_427_EXMPLR, D(10)=>OutputImg2_426_EXMPLR, D(9)=>
      OutputImg2_425_EXMPLR, D(8)=>OutputImg2_424_EXMPLR, D(7)=>
      OutputImg2_423_EXMPLR, D(6)=>OutputImg2_422_EXMPLR, D(5)=>
      OutputImg2_421_EXMPLR, D(4)=>OutputImg2_420_EXMPLR, D(3)=>
      OutputImg2_419_EXMPLR, D(2)=>OutputImg2_418_EXMPLR, D(1)=>
      OutputImg2_417_EXMPLR, D(0)=>OutputImg2_416_EXMPLR, EN=>nx23822, F(15)
      =>ImgReg1IN_431, F(14)=>ImgReg1IN_430, F(13)=>ImgReg1IN_429, F(12)=>
      ImgReg1IN_428, F(11)=>ImgReg1IN_427, F(10)=>ImgReg1IN_426, F(9)=>
      ImgReg1IN_425, F(8)=>ImgReg1IN_424, F(7)=>ImgReg1IN_423, F(6)=>
      ImgReg1IN_422, F(5)=>ImgReg1IN_421, F(4)=>ImgReg1IN_420, F(3)=>
      ImgReg1IN_419, F(2)=>ImgReg1IN_418, F(1)=>ImgReg1IN_417, F(0)=>
      ImgReg1IN_416);
   loop3_26_TriState2U : triStateBuffer_16 port map ( D(15)=>
      OutputImg3_431_EXMPLR, D(14)=>OutputImg3_430_EXMPLR, D(13)=>
      OutputImg3_429_EXMPLR, D(12)=>OutputImg3_428_EXMPLR, D(11)=>
      OutputImg3_427_EXMPLR, D(10)=>OutputImg3_426_EXMPLR, D(9)=>
      OutputImg3_425_EXMPLR, D(8)=>OutputImg3_424_EXMPLR, D(7)=>
      OutputImg3_423_EXMPLR, D(6)=>OutputImg3_422_EXMPLR, D(5)=>
      OutputImg3_421_EXMPLR, D(4)=>OutputImg3_420_EXMPLR, D(3)=>
      OutputImg3_419_EXMPLR, D(2)=>OutputImg3_418_EXMPLR, D(1)=>
      OutputImg3_417_EXMPLR, D(0)=>OutputImg3_416_EXMPLR, EN=>nx23822, F(15)
      =>ImgReg2IN_431, F(14)=>ImgReg2IN_430, F(13)=>ImgReg2IN_429, F(12)=>
      ImgReg2IN_428, F(11)=>ImgReg2IN_427, F(10)=>ImgReg2IN_426, F(9)=>
      ImgReg2IN_425, F(8)=>ImgReg2IN_424, F(7)=>ImgReg2IN_423, F(6)=>
      ImgReg2IN_422, F(5)=>ImgReg2IN_421, F(4)=>ImgReg2IN_420, F(3)=>
      ImgReg2IN_419, F(2)=>ImgReg2IN_418, F(1)=>ImgReg2IN_417, F(0)=>
      ImgReg2IN_416);
   loop3_26_TriState3U : triStateBuffer_16 port map ( D(15)=>
      OutputImg4_431_EXMPLR, D(14)=>OutputImg4_430_EXMPLR, D(13)=>
      OutputImg4_429_EXMPLR, D(12)=>OutputImg4_428_EXMPLR, D(11)=>
      OutputImg4_427_EXMPLR, D(10)=>OutputImg4_426_EXMPLR, D(9)=>
      OutputImg4_425_EXMPLR, D(8)=>OutputImg4_424_EXMPLR, D(7)=>
      OutputImg4_423_EXMPLR, D(6)=>OutputImg4_422_EXMPLR, D(5)=>
      OutputImg4_421_EXMPLR, D(4)=>OutputImg4_420_EXMPLR, D(3)=>
      OutputImg4_419_EXMPLR, D(2)=>OutputImg4_418_EXMPLR, D(1)=>
      OutputImg4_417_EXMPLR, D(0)=>OutputImg4_416_EXMPLR, EN=>nx23824, F(15)
      =>ImgReg3IN_431, F(14)=>ImgReg3IN_430, F(13)=>ImgReg3IN_429, F(12)=>
      ImgReg3IN_428, F(11)=>ImgReg3IN_427, F(10)=>ImgReg3IN_426, F(9)=>
      ImgReg3IN_425, F(8)=>ImgReg3IN_424, F(7)=>ImgReg3IN_423, F(6)=>
      ImgReg3IN_422, F(5)=>ImgReg3IN_421, F(4)=>ImgReg3IN_420, F(3)=>
      ImgReg3IN_419, F(2)=>ImgReg3IN_418, F(1)=>ImgReg3IN_417, F(0)=>
      ImgReg3IN_416);
   loop3_26_TriState4U : triStateBuffer_16 port map ( D(15)=>
      OutputImg5_431_EXMPLR, D(14)=>OutputImg5_430_EXMPLR, D(13)=>
      OutputImg5_429_EXMPLR, D(12)=>OutputImg5_428_EXMPLR, D(11)=>
      OutputImg5_427_EXMPLR, D(10)=>OutputImg5_426_EXMPLR, D(9)=>
      OutputImg5_425_EXMPLR, D(8)=>OutputImg5_424_EXMPLR, D(7)=>
      OutputImg5_423_EXMPLR, D(6)=>OutputImg5_422_EXMPLR, D(5)=>
      OutputImg5_421_EXMPLR, D(4)=>OutputImg5_420_EXMPLR, D(3)=>
      OutputImg5_419_EXMPLR, D(2)=>OutputImg5_418_EXMPLR, D(1)=>
      OutputImg5_417_EXMPLR, D(0)=>OutputImg5_416_EXMPLR, EN=>nx23824, F(15)
      =>ImgReg4IN_431, F(14)=>ImgReg4IN_430, F(13)=>ImgReg4IN_429, F(12)=>
      ImgReg4IN_428, F(11)=>ImgReg4IN_427, F(10)=>ImgReg4IN_426, F(9)=>
      ImgReg4IN_425, F(8)=>ImgReg4IN_424, F(7)=>ImgReg4IN_423, F(6)=>
      ImgReg4IN_422, F(5)=>ImgReg4IN_421, F(4)=>ImgReg4IN_420, F(3)=>
      ImgReg4IN_419, F(2)=>ImgReg4IN_418, F(1)=>ImgReg4IN_417, F(0)=>
      ImgReg4IN_416);
   loop3_26_reg1 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_431, D(14)=>
      ImgReg0IN_430, D(13)=>ImgReg0IN_429, D(12)=>ImgReg0IN_428, D(11)=>
      ImgReg0IN_427, D(10)=>ImgReg0IN_426, D(9)=>ImgReg0IN_425, D(8)=>
      ImgReg0IN_424, D(7)=>ImgReg0IN_423, D(6)=>ImgReg0IN_422, D(5)=>
      ImgReg0IN_421, D(4)=>ImgReg0IN_420, D(3)=>ImgReg0IN_419, D(2)=>
      ImgReg0IN_418, D(1)=>ImgReg0IN_417, D(0)=>ImgReg0IN_416, CLK=>nx23984, 
      RST=>RST, EN=>nx23724, Q(15)=>OutputImg0_431_EXMPLR, Q(14)=>
      OutputImg0_430_EXMPLR, Q(13)=>OutputImg0_429_EXMPLR, Q(12)=>
      OutputImg0_428_EXMPLR, Q(11)=>OutputImg0_427_EXMPLR, Q(10)=>
      OutputImg0_426_EXMPLR, Q(9)=>OutputImg0_425_EXMPLR, Q(8)=>
      OutputImg0_424_EXMPLR, Q(7)=>OutputImg0_423_EXMPLR, Q(6)=>
      OutputImg0_422_EXMPLR, Q(5)=>OutputImg0_421_EXMPLR, Q(4)=>
      OutputImg0_420_EXMPLR, Q(3)=>OutputImg0_419_EXMPLR, Q(2)=>
      OutputImg0_418_EXMPLR, Q(1)=>OutputImg0_417_EXMPLR, Q(0)=>
      OutputImg0_416_EXMPLR);
   loop3_26_reg2 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_431, D(14)=>
      ImgReg1IN_430, D(13)=>ImgReg1IN_429, D(12)=>ImgReg1IN_428, D(11)=>
      ImgReg1IN_427, D(10)=>ImgReg1IN_426, D(9)=>ImgReg1IN_425, D(8)=>
      ImgReg1IN_424, D(7)=>ImgReg1IN_423, D(6)=>ImgReg1IN_422, D(5)=>
      ImgReg1IN_421, D(4)=>ImgReg1IN_420, D(3)=>ImgReg1IN_419, D(2)=>
      ImgReg1IN_418, D(1)=>ImgReg1IN_417, D(0)=>ImgReg1IN_416, CLK=>nx23986, 
      RST=>RST, EN=>nx23734, Q(15)=>OutputImg1_431_EXMPLR, Q(14)=>
      OutputImg1_430_EXMPLR, Q(13)=>OutputImg1_429_EXMPLR, Q(12)=>
      OutputImg1_428_EXMPLR, Q(11)=>OutputImg1_427_EXMPLR, Q(10)=>
      OutputImg1_426_EXMPLR, Q(9)=>OutputImg1_425_EXMPLR, Q(8)=>
      OutputImg1_424_EXMPLR, Q(7)=>OutputImg1_423_EXMPLR, Q(6)=>
      OutputImg1_422_EXMPLR, Q(5)=>OutputImg1_421_EXMPLR, Q(4)=>
      OutputImg1_420_EXMPLR, Q(3)=>OutputImg1_419_EXMPLR, Q(2)=>
      OutputImg1_418_EXMPLR, Q(1)=>OutputImg1_417_EXMPLR, Q(0)=>
      OutputImg1_416_EXMPLR);
   loop3_26_reg3 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_431, D(14)=>
      ImgReg2IN_430, D(13)=>ImgReg2IN_429, D(12)=>ImgReg2IN_428, D(11)=>
      ImgReg2IN_427, D(10)=>ImgReg2IN_426, D(9)=>ImgReg2IN_425, D(8)=>
      ImgReg2IN_424, D(7)=>ImgReg2IN_423, D(6)=>ImgReg2IN_422, D(5)=>
      ImgReg2IN_421, D(4)=>ImgReg2IN_420, D(3)=>ImgReg2IN_419, D(2)=>
      ImgReg2IN_418, D(1)=>ImgReg2IN_417, D(0)=>ImgReg2IN_416, CLK=>nx23986, 
      RST=>RST, EN=>nx23744, Q(15)=>OutputImg2_431_EXMPLR, Q(14)=>
      OutputImg2_430_EXMPLR, Q(13)=>OutputImg2_429_EXMPLR, Q(12)=>
      OutputImg2_428_EXMPLR, Q(11)=>OutputImg2_427_EXMPLR, Q(10)=>
      OutputImg2_426_EXMPLR, Q(9)=>OutputImg2_425_EXMPLR, Q(8)=>
      OutputImg2_424_EXMPLR, Q(7)=>OutputImg2_423_EXMPLR, Q(6)=>
      OutputImg2_422_EXMPLR, Q(5)=>OutputImg2_421_EXMPLR, Q(4)=>
      OutputImg2_420_EXMPLR, Q(3)=>OutputImg2_419_EXMPLR, Q(2)=>
      OutputImg2_418_EXMPLR, Q(1)=>OutputImg2_417_EXMPLR, Q(0)=>
      OutputImg2_416_EXMPLR);
   loop3_26_reg4 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_431, D(14)=>
      ImgReg3IN_430, D(13)=>ImgReg3IN_429, D(12)=>ImgReg3IN_428, D(11)=>
      ImgReg3IN_427, D(10)=>ImgReg3IN_426, D(9)=>ImgReg3IN_425, D(8)=>
      ImgReg3IN_424, D(7)=>ImgReg3IN_423, D(6)=>ImgReg3IN_422, D(5)=>
      ImgReg3IN_421, D(4)=>ImgReg3IN_420, D(3)=>ImgReg3IN_419, D(2)=>
      ImgReg3IN_418, D(1)=>ImgReg3IN_417, D(0)=>ImgReg3IN_416, CLK=>nx23988, 
      RST=>RST, EN=>nx23754, Q(15)=>OutputImg3_431_EXMPLR, Q(14)=>
      OutputImg3_430_EXMPLR, Q(13)=>OutputImg3_429_EXMPLR, Q(12)=>
      OutputImg3_428_EXMPLR, Q(11)=>OutputImg3_427_EXMPLR, Q(10)=>
      OutputImg3_426_EXMPLR, Q(9)=>OutputImg3_425_EXMPLR, Q(8)=>
      OutputImg3_424_EXMPLR, Q(7)=>OutputImg3_423_EXMPLR, Q(6)=>
      OutputImg3_422_EXMPLR, Q(5)=>OutputImg3_421_EXMPLR, Q(4)=>
      OutputImg3_420_EXMPLR, Q(3)=>OutputImg3_419_EXMPLR, Q(2)=>
      OutputImg3_418_EXMPLR, Q(1)=>OutputImg3_417_EXMPLR, Q(0)=>
      OutputImg3_416_EXMPLR);
   loop3_26_reg5 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_431, D(14)=>
      ImgReg4IN_430, D(13)=>ImgReg4IN_429, D(12)=>ImgReg4IN_428, D(11)=>
      ImgReg4IN_427, D(10)=>ImgReg4IN_426, D(9)=>ImgReg4IN_425, D(8)=>
      ImgReg4IN_424, D(7)=>ImgReg4IN_423, D(6)=>ImgReg4IN_422, D(5)=>
      ImgReg4IN_421, D(4)=>ImgReg4IN_420, D(3)=>ImgReg4IN_419, D(2)=>
      ImgReg4IN_418, D(1)=>ImgReg4IN_417, D(0)=>ImgReg4IN_416, CLK=>nx23988, 
      RST=>RST, EN=>nx23764, Q(15)=>OutputImg4_431_EXMPLR, Q(14)=>
      OutputImg4_430_EXMPLR, Q(13)=>OutputImg4_429_EXMPLR, Q(12)=>
      OutputImg4_428_EXMPLR, Q(11)=>OutputImg4_427_EXMPLR, Q(10)=>
      OutputImg4_426_EXMPLR, Q(9)=>OutputImg4_425_EXMPLR, Q(8)=>
      OutputImg4_424_EXMPLR, Q(7)=>OutputImg4_423_EXMPLR, Q(6)=>
      OutputImg4_422_EXMPLR, Q(5)=>OutputImg4_421_EXMPLR, Q(4)=>
      OutputImg4_420_EXMPLR, Q(3)=>OutputImg4_419_EXMPLR, Q(2)=>
      OutputImg4_418_EXMPLR, Q(1)=>OutputImg4_417_EXMPLR, Q(0)=>
      OutputImg4_416_EXMPLR);
   loop3_26_reg6 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_431, D(14)=>
      ImgReg5IN_430, D(13)=>ImgReg5IN_429, D(12)=>ImgReg5IN_428, D(11)=>
      ImgReg5IN_427, D(10)=>ImgReg5IN_426, D(9)=>ImgReg5IN_425, D(8)=>
      ImgReg5IN_424, D(7)=>ImgReg5IN_423, D(6)=>ImgReg5IN_422, D(5)=>
      ImgReg5IN_421, D(4)=>ImgReg5IN_420, D(3)=>ImgReg5IN_419, D(2)=>
      ImgReg5IN_418, D(1)=>ImgReg5IN_417, D(0)=>ImgReg5IN_416, CLK=>nx23990, 
      RST=>RST, EN=>nx23774, Q(15)=>OutputImg5_431_EXMPLR, Q(14)=>
      OutputImg5_430_EXMPLR, Q(13)=>OutputImg5_429_EXMPLR, Q(12)=>
      OutputImg5_428_EXMPLR, Q(11)=>OutputImg5_427_EXMPLR, Q(10)=>
      OutputImg5_426_EXMPLR, Q(9)=>OutputImg5_425_EXMPLR, Q(8)=>
      OutputImg5_424_EXMPLR, Q(7)=>OutputImg5_423_EXMPLR, Q(6)=>
      OutputImg5_422_EXMPLR, Q(5)=>OutputImg5_421_EXMPLR, Q(4)=>
      OutputImg5_420_EXMPLR, Q(3)=>OutputImg5_419_EXMPLR, Q(2)=>
      OutputImg5_418_EXMPLR, Q(1)=>OutputImg5_417_EXMPLR, Q(0)=>
      OutputImg5_416_EXMPLR);
   TriState00L : triStateBuffer_16 port map ( D(15)=>OutputImg0_15_EXMPLR, 
      D(14)=>OutputImg0_14_EXMPLR, D(13)=>OutputImg0_13_EXMPLR, D(12)=>
      OutputImg0_12_EXMPLR, D(11)=>OutputImg0_11_EXMPLR, D(10)=>
      OutputImg0_10_EXMPLR, D(9)=>OutputImg0_9_EXMPLR, D(8)=>
      OutputImg0_8_EXMPLR, D(7)=>OutputImg0_7_EXMPLR, D(6)=>
      OutputImg0_6_EXMPLR, D(5)=>OutputImg0_5_EXMPLR, D(4)=>
      OutputImg0_4_EXMPLR, D(3)=>OutputImg0_3_EXMPLR, D(2)=>
      OutputImg0_2_EXMPLR, D(1)=>OutputImg0_1_EXMPLR, D(0)=>
      OutputImg0_0_EXMPLR, EN=>nx23712, F(15)=>ImgReg0IN_447, F(14)=>
      ImgReg0IN_446, F(13)=>ImgReg0IN_445, F(12)=>ImgReg0IN_444, F(11)=>
      ImgReg0IN_443, F(10)=>ImgReg0IN_442, F(9)=>ImgReg0IN_441, F(8)=>
      ImgReg0IN_440, F(7)=>ImgReg0IN_439, F(6)=>ImgReg0IN_438, F(5)=>
      ImgReg0IN_437, F(4)=>ImgReg0IN_436, F(3)=>ImgReg0IN_435, F(2)=>
      ImgReg0IN_434, F(1)=>ImgReg0IN_433, F(0)=>ImgReg0IN_432);
   TriState11L : triStateBuffer_16 port map ( D(15)=>OutputImg1_15_EXMPLR, 
      D(14)=>OutputImg1_14_EXMPLR, D(13)=>OutputImg1_13_EXMPLR, D(12)=>
      OutputImg1_12_EXMPLR, D(11)=>OutputImg1_11_EXMPLR, D(10)=>
      OutputImg1_10_EXMPLR, D(9)=>OutputImg1_9_EXMPLR, D(8)=>
      OutputImg1_8_EXMPLR, D(7)=>OutputImg1_7_EXMPLR, D(6)=>
      OutputImg1_6_EXMPLR, D(5)=>OutputImg1_5_EXMPLR, D(4)=>
      OutputImg1_4_EXMPLR, D(3)=>OutputImg1_3_EXMPLR, D(2)=>
      OutputImg1_2_EXMPLR, D(1)=>OutputImg1_1_EXMPLR, D(0)=>
      OutputImg1_0_EXMPLR, EN=>nx23712, F(15)=>ImgReg1IN_447, F(14)=>
      ImgReg1IN_446, F(13)=>ImgReg1IN_445, F(12)=>ImgReg1IN_444, F(11)=>
      ImgReg1IN_443, F(10)=>ImgReg1IN_442, F(9)=>ImgReg1IN_441, F(8)=>
      ImgReg1IN_440, F(7)=>ImgReg1IN_439, F(6)=>ImgReg1IN_438, F(5)=>
      ImgReg1IN_437, F(4)=>ImgReg1IN_436, F(3)=>ImgReg1IN_435, F(2)=>
      ImgReg1IN_434, F(1)=>ImgReg1IN_433, F(0)=>ImgReg1IN_432);
   TriState22L : triStateBuffer_16 port map ( D(15)=>OutputImg2_15_EXMPLR, 
      D(14)=>OutputImg2_14_EXMPLR, D(13)=>OutputImg2_13_EXMPLR, D(12)=>
      OutputImg2_12_EXMPLR, D(11)=>OutputImg2_11_EXMPLR, D(10)=>
      OutputImg2_10_EXMPLR, D(9)=>OutputImg2_9_EXMPLR, D(8)=>
      OutputImg2_8_EXMPLR, D(7)=>OutputImg2_7_EXMPLR, D(6)=>
      OutputImg2_6_EXMPLR, D(5)=>OutputImg2_5_EXMPLR, D(4)=>
      OutputImg2_4_EXMPLR, D(3)=>OutputImg2_3_EXMPLR, D(2)=>
      OutputImg2_2_EXMPLR, D(1)=>OutputImg2_1_EXMPLR, D(0)=>
      OutputImg2_0_EXMPLR, EN=>nx23712, F(15)=>ImgReg2IN_447, F(14)=>
      ImgReg2IN_446, F(13)=>ImgReg2IN_445, F(12)=>ImgReg2IN_444, F(11)=>
      ImgReg2IN_443, F(10)=>ImgReg2IN_442, F(9)=>ImgReg2IN_441, F(8)=>
      ImgReg2IN_440, F(7)=>ImgReg2IN_439, F(6)=>ImgReg2IN_438, F(5)=>
      ImgReg2IN_437, F(4)=>ImgReg2IN_436, F(3)=>ImgReg2IN_435, F(2)=>
      ImgReg2IN_434, F(1)=>ImgReg2IN_433, F(0)=>ImgReg2IN_432);
   TriState33L : triStateBuffer_16 port map ( D(15)=>OutputImg3_15_EXMPLR, 
      D(14)=>OutputImg3_14_EXMPLR, D(13)=>OutputImg3_13_EXMPLR, D(12)=>
      OutputImg3_12_EXMPLR, D(11)=>OutputImg3_11_EXMPLR, D(10)=>
      OutputImg3_10_EXMPLR, D(9)=>OutputImg3_9_EXMPLR, D(8)=>
      OutputImg3_8_EXMPLR, D(7)=>OutputImg3_7_EXMPLR, D(6)=>
      OutputImg3_6_EXMPLR, D(5)=>OutputImg3_5_EXMPLR, D(4)=>
      OutputImg3_4_EXMPLR, D(3)=>OutputImg3_3_EXMPLR, D(2)=>
      OutputImg3_2_EXMPLR, D(1)=>OutputImg3_1_EXMPLR, D(0)=>
      OutputImg3_0_EXMPLR, EN=>nx23712, F(15)=>ImgReg3IN_447, F(14)=>
      ImgReg3IN_446, F(13)=>ImgReg3IN_445, F(12)=>ImgReg3IN_444, F(11)=>
      ImgReg3IN_443, F(10)=>ImgReg3IN_442, F(9)=>ImgReg3IN_441, F(8)=>
      ImgReg3IN_440, F(7)=>ImgReg3IN_439, F(6)=>ImgReg3IN_438, F(5)=>
      ImgReg3IN_437, F(4)=>ImgReg3IN_436, F(3)=>ImgReg3IN_435, F(2)=>
      ImgReg3IN_434, F(1)=>ImgReg3IN_433, F(0)=>ImgReg3IN_432);
   TriState44L : triStateBuffer_16 port map ( D(15)=>OutputImg4_15_EXMPLR, 
      D(14)=>OutputImg4_14_EXMPLR, D(13)=>OutputImg4_13_EXMPLR, D(12)=>
      OutputImg4_12_EXMPLR, D(11)=>OutputImg4_11_EXMPLR, D(10)=>
      OutputImg4_10_EXMPLR, D(9)=>OutputImg4_9_EXMPLR, D(8)=>
      OutputImg4_8_EXMPLR, D(7)=>OutputImg4_7_EXMPLR, D(6)=>
      OutputImg4_6_EXMPLR, D(5)=>OutputImg4_5_EXMPLR, D(4)=>
      OutputImg4_4_EXMPLR, D(3)=>OutputImg4_3_EXMPLR, D(2)=>
      OutputImg4_2_EXMPLR, D(1)=>OutputImg4_1_EXMPLR, D(0)=>
      OutputImg4_0_EXMPLR, EN=>nx23712, F(15)=>ImgReg4IN_447, F(14)=>
      ImgReg4IN_446, F(13)=>ImgReg4IN_445, F(12)=>ImgReg4IN_444, F(11)=>
      ImgReg4IN_443, F(10)=>ImgReg4IN_442, F(9)=>ImgReg4IN_441, F(8)=>
      ImgReg4IN_440, F(7)=>ImgReg4IN_439, F(6)=>ImgReg4IN_438, F(5)=>
      ImgReg4IN_437, F(4)=>ImgReg4IN_436, F(3)=>ImgReg4IN_435, F(2)=>
      ImgReg4IN_434, F(1)=>ImgReg4IN_433, F(0)=>ImgReg4IN_432);
   TriState55L : triStateBuffer_16 port map ( D(15)=>OutputImg5_15_EXMPLR, 
      D(14)=>OutputImg5_14_EXMPLR, D(13)=>OutputImg5_13_EXMPLR, D(12)=>
      OutputImg5_12_EXMPLR, D(11)=>OutputImg5_11_EXMPLR, D(10)=>
      OutputImg5_10_EXMPLR, D(9)=>OutputImg5_9_EXMPLR, D(8)=>
      OutputImg5_8_EXMPLR, D(7)=>OutputImg5_7_EXMPLR, D(6)=>
      OutputImg5_6_EXMPLR, D(5)=>OutputImg5_5_EXMPLR, D(4)=>
      OutputImg5_4_EXMPLR, D(3)=>OutputImg5_3_EXMPLR, D(2)=>
      OutputImg5_2_EXMPLR, D(1)=>OutputImg5_1_EXMPLR, D(0)=>
      OutputImg5_0_EXMPLR, EN=>nx23712, F(15)=>ImgReg5IN_447, F(14)=>
      ImgReg5IN_446, F(13)=>ImgReg5IN_445, F(12)=>ImgReg5IN_444, F(11)=>
      ImgReg5IN_443, F(10)=>ImgReg5IN_442, F(9)=>ImgReg5IN_441, F(8)=>
      ImgReg5IN_440, F(7)=>ImgReg5IN_439, F(6)=>ImgReg5IN_438, F(5)=>
      ImgReg5IN_437, F(4)=>ImgReg5IN_436, F(3)=>ImgReg5IN_435, F(2)=>
      ImgReg5IN_434, F(1)=>ImgReg5IN_433, F(0)=>ImgReg5IN_432);
   TriState00N : triStateBuffer_16 port map ( D(15)=>DATA(447), D(14)=>
      DATA(446), D(13)=>DATA(445), D(12)=>DATA(444), D(11)=>DATA(443), D(10)
      =>DATA(442), D(9)=>DATA(441), D(8)=>DATA(440), D(7)=>DATA(439), D(6)=>
      DATA(438), D(5)=>DATA(437), D(4)=>DATA(436), D(3)=>DATA(435), D(2)=>
      DATA(434), D(1)=>DATA(433), D(0)=>DATA(432), EN=>nx23660, F(15)=>
      ImgReg0IN_447, F(14)=>ImgReg0IN_446, F(13)=>ImgReg0IN_445, F(12)=>
      ImgReg0IN_444, F(11)=>ImgReg0IN_443, F(10)=>ImgReg0IN_442, F(9)=>
      ImgReg0IN_441, F(8)=>ImgReg0IN_440, F(7)=>ImgReg0IN_439, F(6)=>
      ImgReg0IN_438, F(5)=>ImgReg0IN_437, F(4)=>ImgReg0IN_436, F(3)=>
      ImgReg0IN_435, F(2)=>ImgReg0IN_434, F(1)=>ImgReg0IN_433, F(0)=>
      ImgReg0IN_432);
   TriState11N : triStateBuffer_16 port map ( D(15)=>DATA(447), D(14)=>
      DATA(446), D(13)=>DATA(445), D(12)=>DATA(444), D(11)=>DATA(443), D(10)
      =>DATA(442), D(9)=>DATA(441), D(8)=>DATA(440), D(7)=>DATA(439), D(6)=>
      DATA(438), D(5)=>DATA(437), D(4)=>DATA(436), D(3)=>DATA(435), D(2)=>
      DATA(434), D(1)=>DATA(433), D(0)=>DATA(432), EN=>nx23648, F(15)=>
      ImgReg1IN_447, F(14)=>ImgReg1IN_446, F(13)=>ImgReg1IN_445, F(12)=>
      ImgReg1IN_444, F(11)=>ImgReg1IN_443, F(10)=>ImgReg1IN_442, F(9)=>
      ImgReg1IN_441, F(8)=>ImgReg1IN_440, F(7)=>ImgReg1IN_439, F(6)=>
      ImgReg1IN_438, F(5)=>ImgReg1IN_437, F(4)=>ImgReg1IN_436, F(3)=>
      ImgReg1IN_435, F(2)=>ImgReg1IN_434, F(1)=>ImgReg1IN_433, F(0)=>
      ImgReg1IN_432);
   TriState22N : triStateBuffer_16 port map ( D(15)=>DATA(447), D(14)=>
      DATA(446), D(13)=>DATA(445), D(12)=>DATA(444), D(11)=>DATA(443), D(10)
      =>DATA(442), D(9)=>DATA(441), D(8)=>DATA(440), D(7)=>DATA(439), D(6)=>
      DATA(438), D(5)=>DATA(437), D(4)=>DATA(436), D(3)=>DATA(435), D(2)=>
      DATA(434), D(1)=>DATA(433), D(0)=>DATA(432), EN=>nx23636, F(15)=>
      ImgReg2IN_447, F(14)=>ImgReg2IN_446, F(13)=>ImgReg2IN_445, F(12)=>
      ImgReg2IN_444, F(11)=>ImgReg2IN_443, F(10)=>ImgReg2IN_442, F(9)=>
      ImgReg2IN_441, F(8)=>ImgReg2IN_440, F(7)=>ImgReg2IN_439, F(6)=>
      ImgReg2IN_438, F(5)=>ImgReg2IN_437, F(4)=>ImgReg2IN_436, F(3)=>
      ImgReg2IN_435, F(2)=>ImgReg2IN_434, F(1)=>ImgReg2IN_433, F(0)=>
      ImgReg2IN_432);
   TriState33N : triStateBuffer_16 port map ( D(15)=>DATA(447), D(14)=>
      DATA(446), D(13)=>DATA(445), D(12)=>DATA(444), D(11)=>DATA(443), D(10)
      =>DATA(442), D(9)=>DATA(441), D(8)=>DATA(440), D(7)=>DATA(439), D(6)=>
      DATA(438), D(5)=>DATA(437), D(4)=>DATA(436), D(3)=>DATA(435), D(2)=>
      DATA(434), D(1)=>DATA(433), D(0)=>DATA(432), EN=>nx23624, F(15)=>
      ImgReg3IN_447, F(14)=>ImgReg3IN_446, F(13)=>ImgReg3IN_445, F(12)=>
      ImgReg3IN_444, F(11)=>ImgReg3IN_443, F(10)=>ImgReg3IN_442, F(9)=>
      ImgReg3IN_441, F(8)=>ImgReg3IN_440, F(7)=>ImgReg3IN_439, F(6)=>
      ImgReg3IN_438, F(5)=>ImgReg3IN_437, F(4)=>ImgReg3IN_436, F(3)=>
      ImgReg3IN_435, F(2)=>ImgReg3IN_434, F(1)=>ImgReg3IN_433, F(0)=>
      ImgReg3IN_432);
   TriState44N : triStateBuffer_16 port map ( D(15)=>DATA(447), D(14)=>
      DATA(446), D(13)=>DATA(445), D(12)=>DATA(444), D(11)=>DATA(443), D(10)
      =>DATA(442), D(9)=>DATA(441), D(8)=>DATA(440), D(7)=>DATA(439), D(6)=>
      DATA(438), D(5)=>DATA(437), D(4)=>DATA(436), D(3)=>DATA(435), D(2)=>
      DATA(434), D(1)=>DATA(433), D(0)=>DATA(432), EN=>nx23612, F(15)=>
      ImgReg4IN_447, F(14)=>ImgReg4IN_446, F(13)=>ImgReg4IN_445, F(12)=>
      ImgReg4IN_444, F(11)=>ImgReg4IN_443, F(10)=>ImgReg4IN_442, F(9)=>
      ImgReg4IN_441, F(8)=>ImgReg4IN_440, F(7)=>ImgReg4IN_439, F(6)=>
      ImgReg4IN_438, F(5)=>ImgReg4IN_437, F(4)=>ImgReg4IN_436, F(3)=>
      ImgReg4IN_435, F(2)=>ImgReg4IN_434, F(1)=>ImgReg4IN_433, F(0)=>
      ImgReg4IN_432);
   TriState55N : triStateBuffer_16 port map ( D(15)=>DATA(447), D(14)=>
      DATA(446), D(13)=>DATA(445), D(12)=>DATA(444), D(11)=>DATA(443), D(10)
      =>DATA(442), D(9)=>DATA(441), D(8)=>DATA(440), D(7)=>DATA(439), D(6)=>
      DATA(438), D(5)=>DATA(437), D(4)=>DATA(436), D(3)=>DATA(435), D(2)=>
      DATA(434), D(1)=>DATA(433), D(0)=>DATA(432), EN=>nx23600, F(15)=>
      ImgReg5IN_447, F(14)=>ImgReg5IN_446, F(13)=>ImgReg5IN_445, F(12)=>
      ImgReg5IN_444, F(11)=>ImgReg5IN_443, F(10)=>ImgReg5IN_442, F(9)=>
      ImgReg5IN_441, F(8)=>ImgReg5IN_440, F(7)=>ImgReg5IN_439, F(6)=>
      ImgReg5IN_438, F(5)=>ImgReg5IN_437, F(4)=>ImgReg5IN_436, F(3)=>
      ImgReg5IN_435, F(2)=>ImgReg5IN_434, F(1)=>ImgReg5IN_433, F(0)=>
      ImgReg5IN_432);
   TriState00U : triStateBuffer_16 port map ( D(15)=>OutputImg1_447_EXMPLR, 
      D(14)=>OutputImg1_446_EXMPLR, D(13)=>OutputImg1_445_EXMPLR, D(12)=>
      OutputImg1_444_EXMPLR, D(11)=>OutputImg1_443_EXMPLR, D(10)=>
      OutputImg1_442_EXMPLR, D(9)=>OutputImg1_441_EXMPLR, D(8)=>
      OutputImg1_440_EXMPLR, D(7)=>OutputImg1_439_EXMPLR, D(6)=>
      OutputImg1_438_EXMPLR, D(5)=>OutputImg1_437_EXMPLR, D(4)=>
      OutputImg1_436_EXMPLR, D(3)=>OutputImg1_435_EXMPLR, D(2)=>
      OutputImg1_434_EXMPLR, D(1)=>OutputImg1_433_EXMPLR, D(0)=>
      OutputImg1_432_EXMPLR, EN=>nx23824, F(15)=>ImgReg0IN_447, F(14)=>
      ImgReg0IN_446, F(13)=>ImgReg0IN_445, F(12)=>ImgReg0IN_444, F(11)=>
      ImgReg0IN_443, F(10)=>ImgReg0IN_442, F(9)=>ImgReg0IN_441, F(8)=>
      ImgReg0IN_440, F(7)=>ImgReg0IN_439, F(6)=>ImgReg0IN_438, F(5)=>
      ImgReg0IN_437, F(4)=>ImgReg0IN_436, F(3)=>ImgReg0IN_435, F(2)=>
      ImgReg0IN_434, F(1)=>ImgReg0IN_433, F(0)=>ImgReg0IN_432);
   TriState11U : triStateBuffer_16 port map ( D(15)=>OutputImg2_447_EXMPLR, 
      D(14)=>OutputImg2_446_EXMPLR, D(13)=>OutputImg2_445_EXMPLR, D(12)=>
      OutputImg2_444_EXMPLR, D(11)=>OutputImg2_443_EXMPLR, D(10)=>
      OutputImg2_442_EXMPLR, D(9)=>OutputImg2_441_EXMPLR, D(8)=>
      OutputImg2_440_EXMPLR, D(7)=>OutputImg2_439_EXMPLR, D(6)=>
      OutputImg2_438_EXMPLR, D(5)=>OutputImg2_437_EXMPLR, D(4)=>
      OutputImg2_436_EXMPLR, D(3)=>OutputImg2_435_EXMPLR, D(2)=>
      OutputImg2_434_EXMPLR, D(1)=>OutputImg2_433_EXMPLR, D(0)=>
      OutputImg2_432_EXMPLR, EN=>nx23824, F(15)=>ImgReg1IN_447, F(14)=>
      ImgReg1IN_446, F(13)=>ImgReg1IN_445, F(12)=>ImgReg1IN_444, F(11)=>
      ImgReg1IN_443, F(10)=>ImgReg1IN_442, F(9)=>ImgReg1IN_441, F(8)=>
      ImgReg1IN_440, F(7)=>ImgReg1IN_439, F(6)=>ImgReg1IN_438, F(5)=>
      ImgReg1IN_437, F(4)=>ImgReg1IN_436, F(3)=>ImgReg1IN_435, F(2)=>
      ImgReg1IN_434, F(1)=>ImgReg1IN_433, F(0)=>ImgReg1IN_432);
   TriState22U : triStateBuffer_16 port map ( D(15)=>OutputImg3_447_EXMPLR, 
      D(14)=>OutputImg3_446_EXMPLR, D(13)=>OutputImg3_445_EXMPLR, D(12)=>
      OutputImg3_444_EXMPLR, D(11)=>OutputImg3_443_EXMPLR, D(10)=>
      OutputImg3_442_EXMPLR, D(9)=>OutputImg3_441_EXMPLR, D(8)=>
      OutputImg3_440_EXMPLR, D(7)=>OutputImg3_439_EXMPLR, D(6)=>
      OutputImg3_438_EXMPLR, D(5)=>OutputImg3_437_EXMPLR, D(4)=>
      OutputImg3_436_EXMPLR, D(3)=>OutputImg3_435_EXMPLR, D(2)=>
      OutputImg3_434_EXMPLR, D(1)=>OutputImg3_433_EXMPLR, D(0)=>
      OutputImg3_432_EXMPLR, EN=>nx23824, F(15)=>ImgReg2IN_447, F(14)=>
      ImgReg2IN_446, F(13)=>ImgReg2IN_445, F(12)=>ImgReg2IN_444, F(11)=>
      ImgReg2IN_443, F(10)=>ImgReg2IN_442, F(9)=>ImgReg2IN_441, F(8)=>
      ImgReg2IN_440, F(7)=>ImgReg2IN_439, F(6)=>ImgReg2IN_438, F(5)=>
      ImgReg2IN_437, F(4)=>ImgReg2IN_436, F(3)=>ImgReg2IN_435, F(2)=>
      ImgReg2IN_434, F(1)=>ImgReg2IN_433, F(0)=>ImgReg2IN_432);
   TriState33U : triStateBuffer_16 port map ( D(15)=>OutputImg4_447_EXMPLR, 
      D(14)=>OutputImg4_446_EXMPLR, D(13)=>OutputImg4_445_EXMPLR, D(12)=>
      OutputImg4_444_EXMPLR, D(11)=>OutputImg4_443_EXMPLR, D(10)=>
      OutputImg4_442_EXMPLR, D(9)=>OutputImg4_441_EXMPLR, D(8)=>
      OutputImg4_440_EXMPLR, D(7)=>OutputImg4_439_EXMPLR, D(6)=>
      OutputImg4_438_EXMPLR, D(5)=>OutputImg4_437_EXMPLR, D(4)=>
      OutputImg4_436_EXMPLR, D(3)=>OutputImg4_435_EXMPLR, D(2)=>
      OutputImg4_434_EXMPLR, D(1)=>OutputImg4_433_EXMPLR, D(0)=>
      OutputImg4_432_EXMPLR, EN=>nx23824, F(15)=>ImgReg3IN_447, F(14)=>
      ImgReg3IN_446, F(13)=>ImgReg3IN_445, F(12)=>ImgReg3IN_444, F(11)=>
      ImgReg3IN_443, F(10)=>ImgReg3IN_442, F(9)=>ImgReg3IN_441, F(8)=>
      ImgReg3IN_440, F(7)=>ImgReg3IN_439, F(6)=>ImgReg3IN_438, F(5)=>
      ImgReg3IN_437, F(4)=>ImgReg3IN_436, F(3)=>ImgReg3IN_435, F(2)=>
      ImgReg3IN_434, F(1)=>ImgReg3IN_433, F(0)=>ImgReg3IN_432);
   TriState44U : triStateBuffer_16 port map ( D(15)=>OutputImg5_447_EXMPLR, 
      D(14)=>OutputImg5_446_EXMPLR, D(13)=>OutputImg5_445_EXMPLR, D(12)=>
      OutputImg5_444_EXMPLR, D(11)=>OutputImg5_443_EXMPLR, D(10)=>
      OutputImg5_442_EXMPLR, D(9)=>OutputImg5_441_EXMPLR, D(8)=>
      OutputImg5_440_EXMPLR, D(7)=>OutputImg5_439_EXMPLR, D(6)=>
      OutputImg5_438_EXMPLR, D(5)=>OutputImg5_437_EXMPLR, D(4)=>
      OutputImg5_436_EXMPLR, D(3)=>OutputImg5_435_EXMPLR, D(2)=>
      OutputImg5_434_EXMPLR, D(1)=>OutputImg5_433_EXMPLR, D(0)=>
      OutputImg5_432_EXMPLR, EN=>nx23824, F(15)=>ImgReg4IN_447, F(14)=>
      ImgReg4IN_446, F(13)=>ImgReg4IN_445, F(12)=>ImgReg4IN_444, F(11)=>
      ImgReg4IN_443, F(10)=>ImgReg4IN_442, F(9)=>ImgReg4IN_441, F(8)=>
      ImgReg4IN_440, F(7)=>ImgReg4IN_439, F(6)=>ImgReg4IN_438, F(5)=>
      ImgReg4IN_437, F(4)=>ImgReg4IN_436, F(3)=>ImgReg4IN_435, F(2)=>
      ImgReg4IN_434, F(1)=>ImgReg4IN_433, F(0)=>ImgReg4IN_432);
   reg11 : nBitRegister_16 port map ( D(15)=>ImgReg0IN_447, D(14)=>
      ImgReg0IN_446, D(13)=>ImgReg0IN_445, D(12)=>ImgReg0IN_444, D(11)=>
      ImgReg0IN_443, D(10)=>ImgReg0IN_442, D(9)=>ImgReg0IN_441, D(8)=>
      ImgReg0IN_440, D(7)=>ImgReg0IN_439, D(6)=>ImgReg0IN_438, D(5)=>
      ImgReg0IN_437, D(4)=>ImgReg0IN_436, D(3)=>ImgReg0IN_435, D(2)=>
      ImgReg0IN_434, D(1)=>ImgReg0IN_433, D(0)=>ImgReg0IN_432, CLK=>nx23990, 
      RST=>RST, EN=>nx23724, Q(15)=>OutputImg0_447_EXMPLR, Q(14)=>
      OutputImg0_446_EXMPLR, Q(13)=>OutputImg0_445_EXMPLR, Q(12)=>
      OutputImg0_444_EXMPLR, Q(11)=>OutputImg0_443_EXMPLR, Q(10)=>
      OutputImg0_442_EXMPLR, Q(9)=>OutputImg0_441_EXMPLR, Q(8)=>
      OutputImg0_440_EXMPLR, Q(7)=>OutputImg0_439_EXMPLR, Q(6)=>
      OutputImg0_438_EXMPLR, Q(5)=>OutputImg0_437_EXMPLR, Q(4)=>
      OutputImg0_436_EXMPLR, Q(3)=>OutputImg0_435_EXMPLR, Q(2)=>
      OutputImg0_434_EXMPLR, Q(1)=>OutputImg0_433_EXMPLR, Q(0)=>
      OutputImg0_432_EXMPLR);
   reg22 : nBitRegister_16 port map ( D(15)=>ImgReg1IN_447, D(14)=>
      ImgReg1IN_446, D(13)=>ImgReg1IN_445, D(12)=>ImgReg1IN_444, D(11)=>
      ImgReg1IN_443, D(10)=>ImgReg1IN_442, D(9)=>ImgReg1IN_441, D(8)=>
      ImgReg1IN_440, D(7)=>ImgReg1IN_439, D(6)=>ImgReg1IN_438, D(5)=>
      ImgReg1IN_437, D(4)=>ImgReg1IN_436, D(3)=>ImgReg1IN_435, D(2)=>
      ImgReg1IN_434, D(1)=>ImgReg1IN_433, D(0)=>ImgReg1IN_432, CLK=>nx23992, 
      RST=>RST, EN=>nx23734, Q(15)=>OutputImg1_447_EXMPLR, Q(14)=>
      OutputImg1_446_EXMPLR, Q(13)=>OutputImg1_445_EXMPLR, Q(12)=>
      OutputImg1_444_EXMPLR, Q(11)=>OutputImg1_443_EXMPLR, Q(10)=>
      OutputImg1_442_EXMPLR, Q(9)=>OutputImg1_441_EXMPLR, Q(8)=>
      OutputImg1_440_EXMPLR, Q(7)=>OutputImg1_439_EXMPLR, Q(6)=>
      OutputImg1_438_EXMPLR, Q(5)=>OutputImg1_437_EXMPLR, Q(4)=>
      OutputImg1_436_EXMPLR, Q(3)=>OutputImg1_435_EXMPLR, Q(2)=>
      OutputImg1_434_EXMPLR, Q(1)=>OutputImg1_433_EXMPLR, Q(0)=>
      OutputImg1_432_EXMPLR);
   reg33 : nBitRegister_16 port map ( D(15)=>ImgReg2IN_447, D(14)=>
      ImgReg2IN_446, D(13)=>ImgReg2IN_445, D(12)=>ImgReg2IN_444, D(11)=>
      ImgReg2IN_443, D(10)=>ImgReg2IN_442, D(9)=>ImgReg2IN_441, D(8)=>
      ImgReg2IN_440, D(7)=>ImgReg2IN_439, D(6)=>ImgReg2IN_438, D(5)=>
      ImgReg2IN_437, D(4)=>ImgReg2IN_436, D(3)=>ImgReg2IN_435, D(2)=>
      ImgReg2IN_434, D(1)=>ImgReg2IN_433, D(0)=>ImgReg2IN_432, CLK=>nx23992, 
      RST=>RST, EN=>nx23744, Q(15)=>OutputImg2_447_EXMPLR, Q(14)=>
      OutputImg2_446_EXMPLR, Q(13)=>OutputImg2_445_EXMPLR, Q(12)=>
      OutputImg2_444_EXMPLR, Q(11)=>OutputImg2_443_EXMPLR, Q(10)=>
      OutputImg2_442_EXMPLR, Q(9)=>OutputImg2_441_EXMPLR, Q(8)=>
      OutputImg2_440_EXMPLR, Q(7)=>OutputImg2_439_EXMPLR, Q(6)=>
      OutputImg2_438_EXMPLR, Q(5)=>OutputImg2_437_EXMPLR, Q(4)=>
      OutputImg2_436_EXMPLR, Q(3)=>OutputImg2_435_EXMPLR, Q(2)=>
      OutputImg2_434_EXMPLR, Q(1)=>OutputImg2_433_EXMPLR, Q(0)=>
      OutputImg2_432_EXMPLR);
   reg44 : nBitRegister_16 port map ( D(15)=>ImgReg3IN_447, D(14)=>
      ImgReg3IN_446, D(13)=>ImgReg3IN_445, D(12)=>ImgReg3IN_444, D(11)=>
      ImgReg3IN_443, D(10)=>ImgReg3IN_442, D(9)=>ImgReg3IN_441, D(8)=>
      ImgReg3IN_440, D(7)=>ImgReg3IN_439, D(6)=>ImgReg3IN_438, D(5)=>
      ImgReg3IN_437, D(4)=>ImgReg3IN_436, D(3)=>ImgReg3IN_435, D(2)=>
      ImgReg3IN_434, D(1)=>ImgReg3IN_433, D(0)=>ImgReg3IN_432, CLK=>nx23994, 
      RST=>RST, EN=>nx23754, Q(15)=>OutputImg3_447_EXMPLR, Q(14)=>
      OutputImg3_446_EXMPLR, Q(13)=>OutputImg3_445_EXMPLR, Q(12)=>
      OutputImg3_444_EXMPLR, Q(11)=>OutputImg3_443_EXMPLR, Q(10)=>
      OutputImg3_442_EXMPLR, Q(9)=>OutputImg3_441_EXMPLR, Q(8)=>
      OutputImg3_440_EXMPLR, Q(7)=>OutputImg3_439_EXMPLR, Q(6)=>
      OutputImg3_438_EXMPLR, Q(5)=>OutputImg3_437_EXMPLR, Q(4)=>
      OutputImg3_436_EXMPLR, Q(3)=>OutputImg3_435_EXMPLR, Q(2)=>
      OutputImg3_434_EXMPLR, Q(1)=>OutputImg3_433_EXMPLR, Q(0)=>
      OutputImg3_432_EXMPLR);
   reg55 : nBitRegister_16 port map ( D(15)=>ImgReg4IN_447, D(14)=>
      ImgReg4IN_446, D(13)=>ImgReg4IN_445, D(12)=>ImgReg4IN_444, D(11)=>
      ImgReg4IN_443, D(10)=>ImgReg4IN_442, D(9)=>ImgReg4IN_441, D(8)=>
      ImgReg4IN_440, D(7)=>ImgReg4IN_439, D(6)=>ImgReg4IN_438, D(5)=>
      ImgReg4IN_437, D(4)=>ImgReg4IN_436, D(3)=>ImgReg4IN_435, D(2)=>
      ImgReg4IN_434, D(1)=>ImgReg4IN_433, D(0)=>ImgReg4IN_432, CLK=>nx23994, 
      RST=>RST, EN=>nx23764, Q(15)=>OutputImg4_447_EXMPLR, Q(14)=>
      OutputImg4_446_EXMPLR, Q(13)=>OutputImg4_445_EXMPLR, Q(12)=>
      OutputImg4_444_EXMPLR, Q(11)=>OutputImg4_443_EXMPLR, Q(10)=>
      OutputImg4_442_EXMPLR, Q(9)=>OutputImg4_441_EXMPLR, Q(8)=>
      OutputImg4_440_EXMPLR, Q(7)=>OutputImg4_439_EXMPLR, Q(6)=>
      OutputImg4_438_EXMPLR, Q(5)=>OutputImg4_437_EXMPLR, Q(4)=>
      OutputImg4_436_EXMPLR, Q(3)=>OutputImg4_435_EXMPLR, Q(2)=>
      OutputImg4_434_EXMPLR, Q(1)=>OutputImg4_433_EXMPLR, Q(0)=>
      OutputImg4_432_EXMPLR);
   reg66 : nBitRegister_16 port map ( D(15)=>ImgReg5IN_447, D(14)=>
      ImgReg5IN_446, D(13)=>ImgReg5IN_445, D(12)=>ImgReg5IN_444, D(11)=>
      ImgReg5IN_443, D(10)=>ImgReg5IN_442, D(9)=>ImgReg5IN_441, D(8)=>
      ImgReg5IN_440, D(7)=>ImgReg5IN_439, D(6)=>ImgReg5IN_438, D(5)=>
      ImgReg5IN_437, D(4)=>ImgReg5IN_436, D(3)=>ImgReg5IN_435, D(2)=>
      ImgReg5IN_434, D(1)=>ImgReg5IN_433, D(0)=>ImgReg5IN_432, CLK=>nx23996, 
      RST=>RST, EN=>nx23774, Q(15)=>OutputImg5_447_EXMPLR, Q(14)=>
      OutputImg5_446_EXMPLR, Q(13)=>OutputImg5_445_EXMPLR, Q(12)=>
      OutputImg5_444_EXMPLR, Q(11)=>OutputImg5_443_EXMPLR, Q(10)=>
      OutputImg5_442_EXMPLR, Q(9)=>OutputImg5_441_EXMPLR, Q(8)=>
      OutputImg5_440_EXMPLR, Q(7)=>OutputImg5_439_EXMPLR, Q(6)=>
      OutputImg5_438_EXMPLR, Q(5)=>OutputImg5_437_EXMPLR, Q(4)=>
      OutputImg5_436_EXMPLR, Q(3)=>OutputImg5_435_EXMPLR, Q(2)=>
      OutputImg5_434_EXMPLR, Q(1)=>OutputImg5_433_EXMPLR, Q(0)=>
      OutputImg5_432_EXMPLR);
   ix23555 : inv01 port map ( Y=>NOT_ImgIndic_0, A=>ImgIndic_0_EXMPLR);
   ix23530 : fake_gnd port map ( Y=>firstOperand_15);
   ix23528 : fake_vcc port map ( Y=>PWR);
   ix5 : or02 port map ( Y=>TriImgLeftEn, A0=>nx2, A1=>current_state(10));
   ix3 : and03 port map ( Y=>nx2, A0=>ACK, A1=>WI, A2=>current_state(8));
   ix43 : oai21 port map ( Y=>TriImgRegEn, A0=>ImgIndic_0_EXMPLR, A1=>nx34, 
      B0=>nx23568);
   ix35 : nand02 port map ( Y=>nx34, A0=>current_state(7), A1=>ACK);
   ix29 : nor02ii port map ( Y=>cEnable, A0=>nx23573, A1=>ACK);
   ix23574 : nor04 port map ( Y=>nx23573, A0=>current_state(2), A1=>
      current_state(3), A2=>nx20, A3=>current_state(4));
   ix21 : or02 port map ( Y=>nx20, A0=>current_state(5), A1=>
      current_state(6));
   ix45 : or02 port map ( Y=>cReset, A0=>RST, A1=>current_state(12));
   ix51 : oai21 port map ( Y=>IndRst, A0=>nx23998, A1=>dontTrust, B0=>
      nx23580);
   ix23581 : inv01 port map ( Y=>nx23580, A=>RST);
   ix63 : oai21 port map ( Y=>TriAddEn, A0=>nx23583, A1=>ImgIndic_0_EXMPLR, 
      B0=>nx23573);
   ix23584 : inv01 port map ( Y=>nx23583, A=>current_state(7));
   reg_DFFCLK_dup_0 : dffr port map ( Q=>DFFCLK, QB=>OPEN, D=>PWR, CLK=>
      nx23830, R=>nx34);
   ix23569 : inv01 port map ( Y=>nx23568, A=>cEnable);
   ix23591 : inv01 port map ( Y=>nx23592, A=>ImgEn_5_EXMPLR);
   ix23593 : inv01 port map ( Y=>nx23594, A=>nx23592);
   ix23595 : inv01 port map ( Y=>nx23596, A=>nx23592);
   ix23597 : inv01 port map ( Y=>nx23598, A=>nx23592);
   ix23599 : inv01 port map ( Y=>nx23600, A=>nx23592);
   ix23603 : inv01 port map ( Y=>nx23604, A=>ImgEn_4_EXMPLR);
   ix23605 : inv01 port map ( Y=>nx23606, A=>nx23604);
   ix23607 : inv01 port map ( Y=>nx23608, A=>nx23604);
   ix23609 : inv01 port map ( Y=>nx23610, A=>nx23604);
   ix23611 : inv01 port map ( Y=>nx23612, A=>nx23604);
   ix23615 : inv01 port map ( Y=>nx23616, A=>ImgEn_3_EXMPLR);
   ix23617 : inv01 port map ( Y=>nx23618, A=>nx23616);
   ix23619 : inv01 port map ( Y=>nx23620, A=>nx23616);
   ix23621 : inv01 port map ( Y=>nx23622, A=>nx23616);
   ix23623 : inv01 port map ( Y=>nx23624, A=>nx23616);
   ix23627 : inv01 port map ( Y=>nx23628, A=>ImgEn_2_EXMPLR);
   ix23629 : inv01 port map ( Y=>nx23630, A=>nx23628);
   ix23631 : inv01 port map ( Y=>nx23632, A=>nx23628);
   ix23633 : inv01 port map ( Y=>nx23634, A=>nx23628);
   ix23635 : inv01 port map ( Y=>nx23636, A=>nx23628);
   ix23639 : inv01 port map ( Y=>nx23640, A=>ImgEn_1_EXMPLR);
   ix23641 : inv01 port map ( Y=>nx23642, A=>nx23640);
   ix23643 : inv01 port map ( Y=>nx23644, A=>nx23640);
   ix23645 : inv01 port map ( Y=>nx23646, A=>nx23640);
   ix23647 : inv01 port map ( Y=>nx23648, A=>nx23640);
   ix23651 : inv01 port map ( Y=>nx23652, A=>ImgEn_0_EXMPLR);
   ix23653 : inv01 port map ( Y=>nx23654, A=>nx23652);
   ix23655 : inv01 port map ( Y=>nx23656, A=>nx23652);
   ix23657 : inv01 port map ( Y=>nx23658, A=>nx23652);
   ix23659 : inv01 port map ( Y=>nx23660, A=>nx23652);
   ix23663 : inv01 port map ( Y=>nx23664, A=>TriImgLeftEn);
   ix23665 : inv01 port map ( Y=>nx23666, A=>nx23776);
   ix23667 : inv01 port map ( Y=>nx23668, A=>nx23776);
   ix23669 : inv01 port map ( Y=>nx23670, A=>nx23776);
   ix23671 : inv01 port map ( Y=>nx23672, A=>nx23776);
   ix23673 : inv01 port map ( Y=>nx23674, A=>nx23776);
   ix23675 : inv01 port map ( Y=>nx23676, A=>nx23776);
   ix23677 : inv01 port map ( Y=>nx23678, A=>nx23776);
   ix23679 : inv01 port map ( Y=>nx23680, A=>nx23778);
   ix23681 : inv01 port map ( Y=>nx23682, A=>nx23778);
   ix23683 : inv01 port map ( Y=>nx23684, A=>nx23778);
   ix23685 : inv01 port map ( Y=>nx23686, A=>nx23778);
   ix23687 : inv01 port map ( Y=>nx23688, A=>nx23778);
   ix23689 : inv01 port map ( Y=>nx23690, A=>nx23778);
   ix23691 : inv01 port map ( Y=>nx23692, A=>nx23778);
   ix23693 : inv01 port map ( Y=>nx23694, A=>nx23780);
   ix23695 : inv01 port map ( Y=>nx23696, A=>nx23780);
   ix23697 : inv01 port map ( Y=>nx23698, A=>nx23780);
   ix23699 : inv01 port map ( Y=>nx23700, A=>nx23780);
   ix23701 : inv01 port map ( Y=>nx23702, A=>nx23780);
   ix23703 : inv01 port map ( Y=>nx23704, A=>nx23780);
   ix23705 : inv01 port map ( Y=>nx23706, A=>nx23780);
   ix23707 : inv01 port map ( Y=>nx23708, A=>nx24006);
   ix23709 : inv01 port map ( Y=>nx23710, A=>nx24006);
   ix23711 : inv01 port map ( Y=>nx23712, A=>nx24006);
   ix23717 : inv01 port map ( Y=>nx23718, A=>nx23716);
   ix23719 : inv01 port map ( Y=>nx23720, A=>nx23716);
   ix23721 : inv01 port map ( Y=>nx23722, A=>nx23716);
   ix23723 : inv01 port map ( Y=>nx23724, A=>nx23716);
   ix23727 : inv01 port map ( Y=>nx23728, A=>nx23726);
   ix23729 : inv01 port map ( Y=>nx23730, A=>nx23726);
   ix23731 : inv01 port map ( Y=>nx23732, A=>nx23726);
   ix23733 : inv01 port map ( Y=>nx23734, A=>nx23726);
   ix23737 : inv01 port map ( Y=>nx23738, A=>nx23736);
   ix23739 : inv01 port map ( Y=>nx23740, A=>nx23736);
   ix23741 : inv01 port map ( Y=>nx23742, A=>nx23736);
   ix23743 : inv01 port map ( Y=>nx23744, A=>nx23736);
   ix23747 : inv01 port map ( Y=>nx23748, A=>nx23746);
   ix23749 : inv01 port map ( Y=>nx23750, A=>nx23746);
   ix23751 : inv01 port map ( Y=>nx23752, A=>nx23746);
   ix23753 : inv01 port map ( Y=>nx23754, A=>nx23746);
   ix23757 : inv01 port map ( Y=>nx23758, A=>nx23756);
   ix23759 : inv01 port map ( Y=>nx23760, A=>nx23756);
   ix23761 : inv01 port map ( Y=>nx23762, A=>nx23756);
   ix23763 : inv01 port map ( Y=>nx23764, A=>nx23756);
   ix23767 : inv01 port map ( Y=>nx23768, A=>nx23766);
   ix23769 : inv01 port map ( Y=>nx23770, A=>nx23766);
   ix23771 : inv01 port map ( Y=>nx23772, A=>nx23766);
   ix23773 : inv01 port map ( Y=>nx23774, A=>nx23766);
   ix23775 : inv01 port map ( Y=>nx23776, A=>TriImgLeftEn);
   ix23777 : inv01 port map ( Y=>nx23778, A=>TriImgLeftEn);
   ix23779 : inv01 port map ( Y=>nx23780, A=>TriImgLeftEn);
   ix7 : and02 port map ( Y=>nx23766, A0=>nx24006, A1=>nx23592);
   ix11 : and03 port map ( Y=>nx23756, A0=>nx24006, A1=>nx23998, A2=>nx23604
   );
   ix13 : and03 port map ( Y=>nx23746, A0=>nx24006, A1=>nx23998, A2=>nx23616
   );
   ix15 : and03 port map ( Y=>nx23736, A0=>nx24006, A1=>nx23998, A2=>nx23628
   );
   ix17 : and03 port map ( Y=>nx23726, A0=>nx23664, A1=>nx23998, A2=>nx23640
   );
   ix19 : and03 port map ( Y=>nx23716, A0=>nx23664, A1=>nx23998, A2=>nx23652
   );
   ix23785 : inv01 port map ( Y=>nx23786, A=>nx23998);
   ix23787 : inv01 port map ( Y=>nx23788, A=>nx24000);
   ix23789 : inv01 port map ( Y=>nx23790, A=>nx24000);
   ix23791 : inv01 port map ( Y=>nx23792, A=>nx24000);
   ix23793 : inv01 port map ( Y=>nx23794, A=>nx24000);
   ix23795 : inv01 port map ( Y=>nx23796, A=>nx24000);
   ix23797 : inv01 port map ( Y=>nx23798, A=>nx24000);
   ix23799 : inv01 port map ( Y=>nx23800, A=>nx24000);
   ix23801 : inv01 port map ( Y=>nx23802, A=>nx24002);
   ix23803 : inv01 port map ( Y=>nx23804, A=>nx24002);
   ix23805 : inv01 port map ( Y=>nx23806, A=>nx24002);
   ix23807 : inv01 port map ( Y=>nx23808, A=>nx24002);
   ix23809 : inv01 port map ( Y=>nx23810, A=>nx24002);
   ix23811 : inv01 port map ( Y=>nx23812, A=>nx24002);
   ix23813 : inv01 port map ( Y=>nx23814, A=>nx24002);
   ix23815 : inv01 port map ( Y=>nx23816, A=>nx24004);
   ix23817 : inv01 port map ( Y=>nx23818, A=>nx24004);
   ix23819 : inv01 port map ( Y=>nx23820, A=>nx24004);
   ix23821 : inv01 port map ( Y=>nx23822, A=>nx24004);
   ix23823 : inv01 port map ( Y=>nx23824, A=>nx24004);
   ix23827 : inv02 port map ( Y=>nx23828, A=>nx24008);
   ix23829 : inv02 port map ( Y=>nx23830, A=>nx24008);
   ix23831 : inv02 port map ( Y=>nx23832, A=>nx24008);
   ix23833 : inv02 port map ( Y=>nx23834, A=>nx24008);
   ix23835 : inv02 port map ( Y=>nx23836, A=>nx24008);
   ix23837 : inv02 port map ( Y=>nx23838, A=>nx24008);
   ix23839 : inv02 port map ( Y=>nx23840, A=>nx24008);
   ix23841 : inv02 port map ( Y=>nx23842, A=>nx24010);
   ix23843 : inv02 port map ( Y=>nx23844, A=>nx24010);
   ix23845 : inv02 port map ( Y=>nx23846, A=>nx24010);
   ix23847 : inv02 port map ( Y=>nx23848, A=>nx24010);
   ix23849 : inv02 port map ( Y=>nx23850, A=>nx24010);
   ix23851 : inv02 port map ( Y=>nx23852, A=>nx24010);
   ix23853 : inv02 port map ( Y=>nx23854, A=>nx24010);
   ix23855 : inv02 port map ( Y=>nx23856, A=>nx24012);
   ix23857 : inv02 port map ( Y=>nx23858, A=>nx24012);
   ix23859 : inv02 port map ( Y=>nx23860, A=>nx24012);
   ix23861 : inv02 port map ( Y=>nx23862, A=>nx24012);
   ix23863 : inv02 port map ( Y=>nx23864, A=>nx24012);
   ix23865 : inv02 port map ( Y=>nx23866, A=>nx24012);
   ix23867 : inv02 port map ( Y=>nx23868, A=>nx24012);
   ix23869 : inv02 port map ( Y=>nx23870, A=>nx24014);
   ix23871 : inv02 port map ( Y=>nx23872, A=>nx24014);
   ix23873 : inv02 port map ( Y=>nx23874, A=>nx24014);
   ix23875 : inv02 port map ( Y=>nx23876, A=>nx24014);
   ix23877 : inv02 port map ( Y=>nx23878, A=>nx24014);
   ix23879 : inv02 port map ( Y=>nx23880, A=>nx24014);
   ix23881 : inv02 port map ( Y=>nx23882, A=>nx24014);
   ix23883 : inv02 port map ( Y=>nx23884, A=>nx24016);
   ix23885 : inv02 port map ( Y=>nx23886, A=>nx24016);
   ix23887 : inv02 port map ( Y=>nx23888, A=>nx24016);
   ix23889 : inv02 port map ( Y=>nx23890, A=>nx24016);
   ix23891 : inv02 port map ( Y=>nx23892, A=>nx24016);
   ix23893 : inv02 port map ( Y=>nx23894, A=>nx24016);
   ix23895 : inv02 port map ( Y=>nx23896, A=>nx24016);
   ix23897 : inv02 port map ( Y=>nx23898, A=>nx24018);
   ix23899 : inv02 port map ( Y=>nx23900, A=>nx24018);
   ix23901 : inv02 port map ( Y=>nx23902, A=>nx24018);
   ix23903 : inv02 port map ( Y=>nx23904, A=>nx24018);
   ix23905 : inv02 port map ( Y=>nx23906, A=>nx24018);
   ix23907 : inv02 port map ( Y=>nx23908, A=>nx24018);
   ix23909 : inv02 port map ( Y=>nx23910, A=>nx24018);
   ix23911 : inv02 port map ( Y=>nx23912, A=>nx24020);
   ix23913 : inv02 port map ( Y=>nx23914, A=>nx24020);
   ix23915 : inv02 port map ( Y=>nx23916, A=>nx24020);
   ix23917 : inv02 port map ( Y=>nx23918, A=>nx24020);
   ix23919 : inv02 port map ( Y=>nx23920, A=>nx24020);
   ix23921 : inv02 port map ( Y=>nx23922, A=>nx24020);
   ix23923 : inv02 port map ( Y=>nx23924, A=>nx24020);
   ix23925 : inv02 port map ( Y=>nx23926, A=>nx24022);
   ix23927 : inv02 port map ( Y=>nx23928, A=>nx24022);
   ix23929 : inv02 port map ( Y=>nx23930, A=>nx24022);
   ix23931 : inv02 port map ( Y=>nx23932, A=>nx24022);
   ix23933 : inv02 port map ( Y=>nx23934, A=>nx24022);
   ix23935 : inv02 port map ( Y=>nx23936, A=>nx24022);
   ix23937 : inv02 port map ( Y=>nx23938, A=>nx24022);
   ix23939 : inv02 port map ( Y=>nx23940, A=>nx24024);
   ix23941 : inv02 port map ( Y=>nx23942, A=>nx24024);
   ix23943 : inv02 port map ( Y=>nx23944, A=>nx24024);
   ix23945 : inv02 port map ( Y=>nx23946, A=>nx24024);
   ix23947 : inv02 port map ( Y=>nx23948, A=>nx24024);
   ix23949 : inv02 port map ( Y=>nx23950, A=>nx24024);
   ix23951 : inv02 port map ( Y=>nx23952, A=>nx24024);
   ix23953 : inv02 port map ( Y=>nx23954, A=>nx24026);
   ix23955 : inv02 port map ( Y=>nx23956, A=>nx24026);
   ix23957 : inv02 port map ( Y=>nx23958, A=>nx24026);
   ix23959 : inv02 port map ( Y=>nx23960, A=>nx24026);
   ix23961 : inv02 port map ( Y=>nx23962, A=>nx24026);
   ix23963 : inv02 port map ( Y=>nx23964, A=>nx24026);
   ix23965 : inv02 port map ( Y=>nx23966, A=>nx24026);
   ix23967 : inv02 port map ( Y=>nx23968, A=>nx24028);
   ix23969 : inv02 port map ( Y=>nx23970, A=>nx24028);
   ix23971 : inv02 port map ( Y=>nx23972, A=>nx24028);
   ix23973 : inv02 port map ( Y=>nx23974, A=>nx24028);
   ix23975 : inv02 port map ( Y=>nx23976, A=>nx24028);
   ix23977 : inv02 port map ( Y=>nx23978, A=>nx24028);
   ix23979 : inv02 port map ( Y=>nx23980, A=>nx24028);
   ix23981 : inv02 port map ( Y=>nx23982, A=>nx24030);
   ix23983 : inv02 port map ( Y=>nx23984, A=>nx24030);
   ix23985 : inv02 port map ( Y=>nx23986, A=>nx24030);
   ix23987 : inv02 port map ( Y=>nx23988, A=>nx24030);
   ix23989 : inv02 port map ( Y=>nx23990, A=>nx24030);
   ix23991 : inv02 port map ( Y=>nx23992, A=>nx24030);
   ix23993 : inv02 port map ( Y=>nx23994, A=>nx24030);
   ix23995 : inv02 port map ( Y=>nx23996, A=>nx24032);
   ix23997 : inv02 port map ( Y=>nx23998, A=>current_state(11));
   ix23999 : inv02 port map ( Y=>nx24000, A=>current_state(11));
   ix24001 : inv02 port map ( Y=>nx24002, A=>current_state(11));
   ix24003 : inv02 port map ( Y=>nx24004, A=>current_state(11));
   ix24005 : inv01 port map ( Y=>nx24006, A=>TriImgLeftEn);
   ix24007 : inv02 port map ( Y=>nx24008, A=>CLK);
   ix24009 : inv02 port map ( Y=>nx24010, A=>nx24038);
   ix24011 : inv02 port map ( Y=>nx24012, A=>nx24038);
   ix24013 : inv02 port map ( Y=>nx24014, A=>nx24038);
   ix24015 : inv02 port map ( Y=>nx24016, A=>nx24038);
   ix24017 : inv02 port map ( Y=>nx24018, A=>nx24038);
   ix24019 : inv02 port map ( Y=>nx24020, A=>nx24038);
   ix24021 : inv02 port map ( Y=>nx24022, A=>nx24038);
   ix24023 : inv02 port map ( Y=>nx24024, A=>nx24040);
   ix24025 : inv02 port map ( Y=>nx24026, A=>nx24040);
   ix24027 : inv02 port map ( Y=>nx24028, A=>nx24040);
   ix24029 : inv02 port map ( Y=>nx24030, A=>nx24040);
   ix24031 : inv02 port map ( Y=>nx24032, A=>nx24040);
   ix24037 : inv02 port map ( Y=>nx24038, A=>nx24008);
   ix24039 : inv02 port map ( Y=>nx24040, A=>nx24008);
end archRI ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity FC_adder is
   port (
      a : IN std_logic ;
      b : IN std_logic ;
      cin : IN std_logic ;
      f : OUT std_logic ;
      cout : OUT std_logic) ;
end FC_adder ;

architecture a_FC_adder of FC_adder is
   signal nx0, nx69: std_logic ;

begin
   ix7 : ao22 port map ( Y=>cout, A0=>b, A1=>a, B0=>cin, B1=>nx0);
   ix9 : xnor2 port map ( Y=>f, A0=>nx69, A1=>cin);
   ix70 : xnor2 port map ( Y=>nx69, A0=>a, A1=>b);
   ix1 : inv01 port map ( Y=>nx0, A=>nx69);
end a_FC_adder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity FC_nadder_32 is
   port (
      aa : IN std_logic_vector (31 DOWNTO 0) ;
      bb : IN std_logic_vector (31 DOWNTO 0) ;
      c_cin : IN std_logic ;
      ff : OUT std_logic_vector (31 DOWNTO 0)) ;
end FC_nadder_32 ;

architecture a_FC_nadder of FC_nadder_32 is
   component FC_adder
      port (
         a : IN std_logic ;
         b : IN std_logic ;
         cin : IN std_logic ;
         f : OUT std_logic ;
         cout : OUT std_logic) ;
   end component ;
   signal temp_30, temp_29, temp_28, temp_27, temp_26, temp_25, temp_24, 
      temp_23, temp_22, temp_21, temp_20, temp_19, temp_18, temp_17, temp_16, 
      temp_15, temp_14, temp_13, temp_12, temp_11, temp_10, temp_9, temp_8, 
      temp_7, temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   f0 : FC_adder port map ( a=>aa(0), b=>bb(0), cin=>c_cin, f=>ff(0), cout=>
      temp_0);
   loop1_1_fx : FC_adder port map ( a=>aa(1), b=>bb(1), cin=>temp_0, f=>
      ff(1), cout=>temp_1);
   loop1_2_fx : FC_adder port map ( a=>aa(2), b=>bb(2), cin=>temp_1, f=>
      ff(2), cout=>temp_2);
   loop1_3_fx : FC_adder port map ( a=>aa(3), b=>bb(3), cin=>temp_2, f=>
      ff(3), cout=>temp_3);
   loop1_4_fx : FC_adder port map ( a=>aa(4), b=>bb(4), cin=>temp_3, f=>
      ff(4), cout=>temp_4);
   loop1_5_fx : FC_adder port map ( a=>aa(5), b=>bb(5), cin=>temp_4, f=>
      ff(5), cout=>temp_5);
   loop1_6_fx : FC_adder port map ( a=>aa(6), b=>bb(6), cin=>temp_5, f=>
      ff(6), cout=>temp_6);
   loop1_7_fx : FC_adder port map ( a=>aa(7), b=>bb(7), cin=>temp_6, f=>
      ff(7), cout=>temp_7);
   loop1_8_fx : FC_adder port map ( a=>aa(8), b=>bb(8), cin=>temp_7, f=>
      ff(8), cout=>temp_8);
   loop1_9_fx : FC_adder port map ( a=>aa(9), b=>bb(9), cin=>temp_8, f=>
      ff(9), cout=>temp_9);
   loop1_10_fx : FC_adder port map ( a=>aa(10), b=>bb(10), cin=>temp_9, f=>
      ff(10), cout=>temp_10);
   loop1_11_fx : FC_adder port map ( a=>aa(11), b=>bb(11), cin=>temp_10, f=>
      ff(11), cout=>temp_11);
   loop1_12_fx : FC_adder port map ( a=>aa(12), b=>bb(12), cin=>temp_11, f=>
      ff(12), cout=>temp_12);
   loop1_13_fx : FC_adder port map ( a=>aa(13), b=>bb(13), cin=>temp_12, f=>
      ff(13), cout=>temp_13);
   loop1_14_fx : FC_adder port map ( a=>aa(14), b=>bb(14), cin=>temp_13, f=>
      ff(14), cout=>temp_14);
   loop1_15_fx : FC_adder port map ( a=>aa(15), b=>bb(15), cin=>temp_14, f=>
      ff(15), cout=>temp_15);
   loop1_16_fx : FC_adder port map ( a=>aa(16), b=>bb(16), cin=>temp_15, f=>
      ff(16), cout=>temp_16);
   loop1_17_fx : FC_adder port map ( a=>aa(17), b=>bb(17), cin=>temp_16, f=>
      ff(17), cout=>temp_17);
   loop1_18_fx : FC_adder port map ( a=>aa(18), b=>bb(18), cin=>temp_17, f=>
      ff(18), cout=>temp_18);
   loop1_19_fx : FC_adder port map ( a=>aa(19), b=>bb(19), cin=>temp_18, f=>
      ff(19), cout=>temp_19);
   loop1_20_fx : FC_adder port map ( a=>aa(20), b=>bb(20), cin=>temp_19, f=>
      ff(20), cout=>temp_20);
   loop1_21_fx : FC_adder port map ( a=>aa(21), b=>bb(21), cin=>temp_20, f=>
      ff(21), cout=>temp_21);
   loop1_22_fx : FC_adder port map ( a=>aa(22), b=>bb(22), cin=>temp_21, f=>
      ff(22), cout=>temp_22);
   loop1_23_fx : FC_adder port map ( a=>aa(23), b=>bb(23), cin=>temp_22, f=>
      ff(23), cout=>temp_23);
   loop1_24_fx : FC_adder port map ( a=>aa(24), b=>bb(24), cin=>temp_23, f=>
      ff(24), cout=>temp_24);
   loop1_25_fx : FC_adder port map ( a=>aa(25), b=>bb(25), cin=>temp_24, f=>
      ff(25), cout=>temp_25);
   loop1_26_fx : FC_adder port map ( a=>aa(26), b=>bb(26), cin=>temp_25, f=>
      ff(26), cout=>temp_26);
   loop1_27_fx : FC_adder port map ( a=>aa(27), b=>bb(27), cin=>temp_26, f=>
      ff(27), cout=>temp_27);
   loop1_28_fx : FC_adder port map ( a=>aa(28), b=>bb(28), cin=>temp_27, f=>
      ff(28), cout=>temp_28);
   loop1_29_fx : FC_adder port map ( a=>aa(29), b=>bb(29), cin=>temp_28, f=>
      ff(29), cout=>temp_29);
   loop1_30_fx : FC_adder port map ( a=>aa(30), b=>bb(30), cin=>temp_29, f=>
      ff(30), cout=>temp_30);
   loop1_31_fx : FC_adder port map ( a=>aa(31), b=>bb(31), cin=>temp_30, f=>
      ff(31), cout=>DANGLING(0));
end a_FC_nadder ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Multiplier_16 is
   port (
      A : IN std_logic_vector (15 DOWNTO 0) ;
      B : IN std_logic_vector (15 DOWNTO 0) ;
      F : OUT std_logic_vector (31 DOWNTO 0)) ;
end Multiplier_16 ;

architecture Flow of Multiplier_16 is
   component FC_nadder_32
      port (
         aa : IN std_logic_vector (31 DOWNTO 0) ;
         bb : IN std_logic_vector (31 DOWNTO 0) ;
         c_cin : IN std_logic ;
         ff : OUT std_logic_vector (31 DOWNTO 0)) ;
   end component ;
   signal addout_0_31, addout_0_30, addout_0_29, addout_0_28, addout_0_27, 
      addout_0_26, addout_0_25, addout_0_24, addout_0_23, addout_0_22, 
      addout_0_21, addout_0_20, addout_0_19, addout_0_18, addout_0_17, 
      addout_0_16, addout_0_15, addout_0_14, addout_0_13, addout_0_12, 
      addout_0_11, addout_0_10, addout_0_9, addout_0_8, addout_0_7, 
      addout_0_6, addout_0_5, addout_0_4, addout_0_3, addout_0_2, addout_0_1, 
      addout_0_0, addout_1_31, addout_1_30, addout_1_29, addout_1_28, 
      addout_1_27, addout_1_26, addout_1_25, addout_1_24, addout_1_23, 
      addout_1_22, addout_1_21, addout_1_20, addout_1_19, addout_1_18, 
      addout_1_17, addout_1_16, addout_1_15, addout_1_14, addout_1_13, 
      addout_1_12, addout_1_11, addout_1_10, addout_1_9, addout_1_8, 
      addout_1_7, addout_1_6, addout_1_5, addout_1_4, addout_1_3, addout_1_2, 
      addout_1_1, addout_1_0, addout_2_31, addout_2_30, addout_2_29, 
      addout_2_28, addout_2_27, addout_2_26, addout_2_25, addout_2_24, 
      addout_2_23, addout_2_22, addout_2_21, addout_2_20, addout_2_19, 
      addout_2_18, addout_2_17, addout_2_16, addout_2_15, addout_2_14, 
      addout_2_13, addout_2_12, addout_2_11, addout_2_10, addout_2_9, 
      addout_2_8, addout_2_7, addout_2_6, addout_2_5, addout_2_4, addout_2_3, 
      addout_2_2, addout_2_1, addout_2_0, addout_3_31, addout_3_30, 
      addout_3_29, addout_3_28, addout_3_27, addout_3_26, addout_3_25, 
      addout_3_24, addout_3_23, addout_3_22, addout_3_21, addout_3_20, 
      addout_3_19, addout_3_18, addout_3_17, addout_3_16, addout_3_15, 
      addout_3_14, addout_3_13, addout_3_12, addout_3_11, addout_3_10, 
      addout_3_9, addout_3_8, addout_3_7, addout_3_6, addout_3_5, addout_3_4, 
      addout_3_3, addout_3_2, addout_3_1, addout_3_0, addout_4_31, 
      addout_4_30, addout_4_29, addout_4_28, addout_4_27, addout_4_26, 
      addout_4_25, addout_4_24, addout_4_23, addout_4_22, addout_4_21, 
      addout_4_20, addout_4_19, addout_4_18, addout_4_17, addout_4_16, 
      addout_4_15, addout_4_14, addout_4_13, addout_4_12, addout_4_11, 
      addout_4_10, addout_4_9, addout_4_8, addout_4_7, addout_4_6, 
      addout_4_5, addout_4_4, addout_4_3, addout_4_2, addout_4_1, addout_4_0, 
      addout_5_31, addout_5_30, addout_5_29, addout_5_28, addout_5_27, 
      addout_5_26, addout_5_25, addout_5_24, addout_5_23, addout_5_22, 
      addout_5_21, addout_5_20, addout_5_19, addout_5_18, addout_5_17, 
      addout_5_16, addout_5_15, addout_5_14, addout_5_13, addout_5_12, 
      addout_5_11, addout_5_10, addout_5_9, addout_5_8, addout_5_7, 
      addout_5_6, addout_5_5, addout_5_4, addout_5_3, addout_5_2, addout_5_1, 
      addout_5_0, addout_6_31, addout_6_30, addout_6_29, addout_6_28, 
      addout_6_27, addout_6_26, addout_6_25, addout_6_24, addout_6_23, 
      addout_6_22, addout_6_21, addout_6_20, addout_6_19, addout_6_18, 
      addout_6_17, addout_6_16, addout_6_15, addout_6_14, addout_6_13, 
      addout_6_12, addout_6_11, addout_6_10, addout_6_9, addout_6_8, 
      addout_6_7, addout_6_6, addout_6_5, addout_6_4, addout_6_3, addout_6_2, 
      addout_6_1, addout_6_0, addout_7_31, addout_7_30, addout_7_29, 
      addout_7_28, addout_7_27, addout_7_26, addout_7_25, addout_7_24, 
      addout_7_23, addout_7_22, addout_7_21, addout_7_20, addout_7_19, 
      addout_7_18, addout_7_17, addout_7_16, addout_7_15, addout_7_14, 
      addout_7_13, addout_7_12, addout_7_11, addout_7_10, addout_7_9, 
      addout_7_8, addout_7_7, addout_7_6, addout_7_5, addout_7_4, addout_7_3, 
      addout_7_2, addout_7_1, addout_7_0, addout_8_31, addout_8_30, 
      addout_8_29, addout_8_28, addout_8_27, addout_8_26, addout_8_25, 
      addout_8_24, addout_8_23, addout_8_22, addout_8_21, addout_8_20, 
      addout_8_19, addout_8_18, addout_8_17, addout_8_16, addout_8_15, 
      addout_8_14, addout_8_13, addout_8_12, addout_8_11, addout_8_10, 
      addout_8_9, addout_8_8, addout_8_7, addout_8_6, addout_8_5, addout_8_4, 
      addout_8_3, addout_8_2, addout_8_1, addout_8_0, addout_9_31, 
      addout_9_30, addout_9_29, addout_9_28, addout_9_27, addout_9_26, 
      addout_9_25, addout_9_24, addout_9_23, addout_9_22, addout_9_21, 
      addout_9_20, addout_9_19, addout_9_18, addout_9_17, addout_9_16, 
      addout_9_15, addout_9_14, addout_9_13, addout_9_12, addout_9_11, 
      addout_9_10, addout_9_9, addout_9_8, addout_9_7, addout_9_6, 
      addout_9_5, addout_9_4, addout_9_3, addout_9_2, addout_9_1, addout_9_0, 
      addout_10_31, addout_10_30, addout_10_29, addout_10_28, addout_10_27, 
      addout_10_26, addout_10_25, addout_10_24, addout_10_23, addout_10_22, 
      addout_10_21, addout_10_20, addout_10_19, addout_10_18, addout_10_17, 
      addout_10_16, addout_10_15, addout_10_14, addout_10_13, addout_10_12, 
      addout_10_11, addout_10_10, addout_10_9, addout_10_8, addout_10_7, 
      addout_10_6, addout_10_5, addout_10_4, addout_10_3, addout_10_2, 
      addout_10_1, addout_10_0, addout_11_31, addout_11_30, addout_11_29, 
      addout_11_28, addout_11_27, addout_11_26, addout_11_25, addout_11_24, 
      addout_11_23, addout_11_22, addout_11_21, addout_11_20, addout_11_19, 
      addout_11_18, addout_11_17, addout_11_16, addout_11_15, addout_11_14, 
      addout_11_13, addout_11_12, addout_11_11, addout_11_10, addout_11_9, 
      addout_11_8, addout_11_7, addout_11_6, addout_11_5, addout_11_4, 
      addout_11_3, addout_11_2, addout_11_1, addout_11_0, addout_12_31, 
      addout_12_30, addout_12_29, addout_12_28, addout_12_27, addout_12_26, 
      addout_12_25, addout_12_24, addout_12_23, addout_12_22, addout_12_21, 
      addout_12_20, addout_12_19, addout_12_18, addout_12_17, addout_12_16, 
      addout_12_15, addout_12_14, addout_12_13, addout_12_12, addout_12_11, 
      addout_12_10, addout_12_9, addout_12_8, addout_12_7, addout_12_6, 
      addout_12_5, addout_12_4, addout_12_3, addout_12_2, addout_12_1, 
      addout_12_0, addout_13_31, addout_13_30, addout_13_29, addout_13_28, 
      addout_13_27, addout_13_26, addout_13_25, addout_13_24, addout_13_23, 
      addout_13_22, addout_13_21, addout_13_20, addout_13_19, addout_13_18, 
      addout_13_17, addout_13_16, addout_13_15, addout_13_14, addout_13_13, 
      addout_13_12, addout_13_11, addout_13_10, addout_13_9, addout_13_8, 
      addout_13_7, addout_13_6, addout_13_5, addout_13_4, addout_13_3, 
      addout_13_2, addout_13_1, addout_13_0, addout_14_31, addout_14_30, 
      addout_14_29, addout_14_28, addout_14_27, addout_14_26, addout_14_25, 
      addout_14_24, addout_14_23, addout_14_22, addout_14_21, addout_14_20, 
      addout_14_19, addout_14_18, addout_14_17, addout_14_16, addout_14_15, 
      addout_14_14, addout_14_13, addout_14_12, addout_14_11, addout_14_10, 
      addout_14_9, addout_14_8, addout_14_7, addout_14_6, addout_14_5, 
      addout_14_4, addout_14_3, addout_14_2, addout_14_1, addout_14_0, 
      addout_15_31, addout_15_30, addout_15_29, addout_15_28, addout_15_27, 
      addout_15_26, addout_15_25, addout_15_24, addout_15_23, addout_15_22, 
      addout_15_21, addout_15_20, addout_15_19, addout_15_18, addout_15_17, 
      addout_15_16, addout_15_15, addout_15_14, addout_15_13, addout_15_12, 
      addout_15_11, addout_15_10, addout_15_9, addout_15_8, addout_15_7, 
      addout_15_6, addout_15_5, addout_15_4, addout_15_3, addout_15_2, 
      addout_15_1, addout_15_0, addout_16_31, addout_16_30, addout_16_29, 
      addout_16_28, addout_16_27, addout_16_26, addout_16_25, addout_16_24, 
      addout_16_23, addout_16_22, addout_16_21, addout_16_20, addout_16_19, 
      addout_16_18, addout_16_17, addout_16_16, addout_16_15, addout_16_14, 
      addout_16_13, addout_16_12, addout_16_11, addout_16_10, addout_16_9, 
      addout_16_8, addout_16_7, addout_16_6, addout_16_5, addout_16_4, 
      addout_16_3, addout_16_2, addout_16_1, addout_16_0, addout_17_31, 
      addout_17_30, addout_17_29, addout_17_28, addout_17_27, addout_17_26, 
      addout_17_25, addout_17_24, addout_17_23, addout_17_22, addout_17_21, 
      addout_17_20, addout_17_19, addout_17_18, addout_17_17, addout_17_16, 
      addout_17_15, addout_17_14, addout_17_13, addout_17_12, addout_17_11, 
      addout_17_10, addout_17_9, addout_17_8, addout_17_7, addout_17_6, 
      addout_17_5, addout_17_4, addout_17_3, addout_17_2, addout_17_1, 
      addout_17_0, addout_18_31, addout_18_30, addout_18_29, addout_18_28, 
      addout_18_27, addout_18_26, addout_18_25, addout_18_24, addout_18_23, 
      addout_18_22, addout_18_21, addout_18_20, addout_18_19, addout_18_18, 
      addout_18_17, addout_18_16, addout_18_15, addout_18_14, addout_18_13, 
      addout_18_12, addout_18_11, addout_18_10, addout_18_9, addout_18_8, 
      addout_18_7, addout_18_6, addout_18_5, addout_18_4, addout_18_3, 
      addout_18_2, addout_18_1, addout_18_0, addout_19_31, addout_19_30, 
      addout_19_29, addout_19_28, addout_19_27, addout_19_26, addout_19_25, 
      addout_19_24, addout_19_23, addout_19_22, addout_19_21, addout_19_20, 
      addout_19_19, addout_19_18, addout_19_17, addout_19_16, addout_19_15, 
      addout_19_14, addout_19_13, addout_19_12, addout_19_11, addout_19_10, 
      addout_19_9, addout_19_8, addout_19_7, addout_19_6, addout_19_5, 
      addout_19_4, addout_19_3, addout_19_2, addout_19_1, addout_19_0, 
      addout_20_31, addout_20_30, addout_20_29, addout_20_28, addout_20_27, 
      addout_20_26, addout_20_25, addout_20_24, addout_20_23, addout_20_22, 
      addout_20_21, addout_20_20, addout_20_19, addout_20_18, addout_20_17, 
      addout_20_16, addout_20_15, addout_20_14, addout_20_13, addout_20_12, 
      addout_20_11, addout_20_10, addout_20_9, addout_20_8, addout_20_7, 
      addout_20_6, addout_20_5, addout_20_4, addout_20_3, addout_20_2, 
      addout_20_1, addout_20_0, addout_21_31, addout_21_30, addout_21_29, 
      addout_21_28, addout_21_27, addout_21_26, addout_21_25, addout_21_24, 
      addout_21_23, addout_21_22, addout_21_21, addout_21_20, addout_21_19, 
      addout_21_18, addout_21_17, addout_21_16, addout_21_15, addout_21_14, 
      addout_21_13, addout_21_12, addout_21_11, addout_21_10, addout_21_9, 
      addout_21_8, addout_21_7, addout_21_6, addout_21_5, addout_21_4, 
      addout_21_3, addout_21_2, addout_21_1, addout_21_0, addout_22_31, 
      addout_22_30, addout_22_29, addout_22_28, addout_22_27, addout_22_26, 
      addout_22_25, addout_22_24, addout_22_23, addout_22_22, addout_22_21, 
      addout_22_20, addout_22_19, addout_22_18, addout_22_17, addout_22_16, 
      addout_22_15, addout_22_14, addout_22_13, addout_22_12, addout_22_11, 
      addout_22_10, addout_22_9, addout_22_8, addout_22_7, addout_22_6, 
      addout_22_5, addout_22_4, addout_22_3, addout_22_2, addout_22_1, 
      addout_22_0, addout_23_31, addout_23_30, addout_23_29, addout_23_28, 
      addout_23_27, addout_23_26, addout_23_25, addout_23_24, addout_23_23, 
      addout_23_22, addout_23_21, addout_23_20, addout_23_19, addout_23_18, 
      addout_23_17, addout_23_16, addout_23_15, addout_23_14, addout_23_13, 
      addout_23_12, addout_23_11, addout_23_10, addout_23_9, addout_23_8, 
      addout_23_7, addout_23_6, addout_23_5, addout_23_4, addout_23_3, 
      addout_23_2, addout_23_1, addout_23_0, addout_24_31, addout_24_30, 
      addout_24_29, addout_24_28, addout_24_27, addout_24_26, addout_24_25, 
      addout_24_24, addout_24_23, addout_24_22, addout_24_21, addout_24_20, 
      addout_24_19, addout_24_18, addout_24_17, addout_24_16, addout_24_15, 
      addout_24_14, addout_24_13, addout_24_12, addout_24_11, addout_24_10, 
      addout_24_9, addout_24_8, addout_24_7, addout_24_6, addout_24_5, 
      addout_24_4, addout_24_3, addout_24_2, addout_24_1, addout_24_0, 
      addout_25_31, addout_25_30, addout_25_29, addout_25_28, addout_25_27, 
      addout_25_26, addout_25_25, addout_25_24, addout_25_23, addout_25_22, 
      addout_25_21, addout_25_20, addout_25_19, addout_25_18, addout_25_17, 
      addout_25_16, addout_25_15, addout_25_14, addout_25_13, addout_25_12, 
      addout_25_11, addout_25_10, addout_25_9, addout_25_8, addout_25_7, 
      addout_25_6, addout_25_5, addout_25_4, addout_25_3, addout_25_2, 
      addout_25_1, addout_25_0, addout_26_31, addout_26_30, addout_26_29, 
      addout_26_28, addout_26_27, addout_26_26, addout_26_25, addout_26_24, 
      addout_26_23, addout_26_22, addout_26_21, addout_26_20, addout_26_19, 
      addout_26_18, addout_26_17, addout_26_16, addout_26_15, addout_26_14, 
      addout_26_13, addout_26_12, addout_26_11, addout_26_10, addout_26_9, 
      addout_26_8, addout_26_7, addout_26_6, addout_26_5, addout_26_4, 
      addout_26_3, addout_26_2, addout_26_1, addout_26_0, addout_27_31, 
      addout_27_30, addout_27_29, addout_27_28, addout_27_27, addout_27_26, 
      addout_27_25, addout_27_24, addout_27_23, addout_27_22, addout_27_21, 
      addout_27_20, addout_27_19, addout_27_18, addout_27_17, addout_27_16, 
      addout_27_15, addout_27_14, addout_27_13, addout_27_12, addout_27_11, 
      addout_27_10, addout_27_9, addout_27_8, addout_27_7, addout_27_6, 
      addout_27_5, addout_27_4, addout_27_3, addout_27_2, addout_27_1, 
      addout_27_0, addout_28_31, addout_28_30, addout_28_29, addout_28_28, 
      addout_28_27, addout_28_26, addout_28_25, addout_28_24, addout_28_23, 
      addout_28_22, addout_28_21, addout_28_20, addout_28_19, addout_28_18, 
      addout_28_17, addout_28_16, addout_28_15, addout_28_14, addout_28_13, 
      addout_28_12, addout_28_11, addout_28_10, addout_28_9, addout_28_8, 
      addout_28_7, addout_28_6, addout_28_5, addout_28_4, addout_28_3, 
      addout_28_2, addout_28_1, addout_28_0, addout_29_31, addout_29_30, 
      addout_29_29, addout_29_28, addout_29_27, addout_29_26, addout_29_25, 
      addout_29_24, addout_29_23, addout_29_22, addout_29_21, addout_29_20, 
      addout_29_19, addout_29_18, addout_29_17, addout_29_16, addout_29_15, 
      addout_29_14, addout_29_13, addout_29_12, addout_29_11, addout_29_10, 
      addout_29_9, addout_29_8, addout_29_7, addout_29_6, addout_29_5, 
      addout_29_4, addout_29_3, addout_29_2, addout_29_1, addout_29_0, 
      op2_0_15, op2_0_14, op2_0_13, op2_0_12, op2_0_11, op2_0_10, op2_0_9, 
      op2_0_8, op2_0_7, op2_0_6, op2_0_5, op2_0_4, op2_0_3, op2_0_2, op2_0_1, 
      op2_1_16, op2_1_15, op2_1_14, op2_1_13, op2_1_12, op2_1_11, op2_1_10, 
      op2_1_9, op2_1_8, op2_1_7, op2_1_6, op2_1_5, op2_1_4, op2_1_3, op2_1_2, 
      op2_2_17, op2_2_16, op2_2_15, op2_2_14, op2_2_13, op2_2_12, op2_2_11, 
      op2_2_10, op2_2_9, op2_2_8, op2_2_7, op2_2_6, op2_2_5, op2_2_4, 
      op2_2_3, op2_3_18, op2_3_17, op2_3_16, op2_3_15, op2_3_14, op2_3_13, 
      op2_3_12, op2_3_11, op2_3_10, op2_3_9, op2_3_8, op2_3_7, op2_3_6, 
      op2_3_5, op2_3_4, op2_4_19, op2_4_18, op2_4_17, op2_4_16, op2_4_15, 
      op2_4_14, op2_4_13, op2_4_12, op2_4_11, op2_4_10, op2_4_9, op2_4_8, 
      op2_4_7, op2_4_6, op2_4_5, op2_5_20, op2_5_19, op2_5_18, op2_5_17, 
      op2_5_16, op2_5_15, op2_5_14, op2_5_13, op2_5_12, op2_5_11, op2_5_10, 
      op2_5_9, op2_5_8, op2_5_7, op2_5_6, op2_6_21, op2_6_20, op2_6_19, 
      op2_6_18, op2_6_17, op2_6_16, op2_6_15, op2_6_14, op2_6_13, op2_6_12, 
      op2_6_11, op2_6_10, op2_6_9, op2_6_8, op2_6_7, op2_7_22, op2_7_21, 
      op2_7_20, op2_7_19, op2_7_18, op2_7_17, op2_7_16, op2_7_15, op2_7_14, 
      op2_7_13, op2_7_12, op2_7_11, op2_7_10, op2_7_9, op2_7_8, op2_8_23, 
      op2_8_22, op2_8_21, op2_8_20, op2_8_19, op2_8_18, op2_8_17, op2_8_16, 
      op2_8_15, op2_8_14, op2_8_13, op2_8_12, op2_8_11, op2_8_10, op2_8_9, 
      op2_9_24, op2_9_23, op2_9_22, op2_9_21, op2_9_20, op2_9_19, op2_9_18, 
      op2_9_17, op2_9_16, op2_9_15, op2_9_14, op2_9_13, op2_9_12, op2_9_11, 
      op2_9_10, op2_10_26, op2_10_25, op2_10_24, op2_10_23, op2_10_22, 
      op2_10_21, op2_10_20, op2_10_19, op2_10_18, op2_10_17, op2_10_16, 
      op2_10_15, op2_10_14, op2_10_13, op2_10_12, op2_10_11, op2_11_27, 
      op2_11_26, op2_11_25, op2_11_24, op2_11_23, op2_11_22, op2_11_21, 
      op2_11_20, op2_11_19, op2_11_18, op2_11_17, op2_11_16, op2_11_15, 
      op2_11_14, op2_11_13, op2_11_12, op2_12_28, op2_12_27, op2_12_26, 
      op2_12_25, op2_12_24, op2_12_23, op2_12_22, op2_12_21, op2_12_20, 
      op2_12_19, op2_12_18, op2_12_17, op2_12_16, op2_12_15, op2_12_14, 
      op2_12_13, op2_13_29, op2_13_28, op2_13_27, op2_13_26, op2_13_25, 
      op2_13_24, op2_13_23, op2_13_22, op2_13_21, op2_13_20, op2_13_19, 
      op2_13_18, op2_13_17, op2_13_16, op2_13_15, op2_13_14, op2_14_30, 
      op2_14_29, op2_14_28, op2_14_27, op2_14_26, op1_14, op1_13, op1_12, 
      op1_11, op1_10, op1_9, op1_8, op1_7, op1_6, op1_5, op1_4, op1_3, op1_2, 
      op1_1, op1_0, addout_31_31, nx5768, nx5770, nx5772, nx5774, nx5776, 
      nx5778, nx5780, nx5782, nx5784, nx5786, nx5788, nx5790, nx5792, nx5794, 
      nx5796, nx5798, nx5800, nx5802, nx5804, nx5806, nx5808, nx5810, nx5812, 
      nx5814, nx5816, nx5818, nx5820, nx5822, nx5824, nx5826, nx5828, nx5830, 
      nx5832, nx5834, nx5836, nx5838, nx5840, nx5842, nx5844, nx5846, nx5848, 
      nx5850, nx5852, nx5854, nx5856, nx5858, nx5860, nx5862, nx5864, nx5866, 
      nx5868, nx5870, nx5872, nx5874, nx5876, nx5878, nx5880, nx5882, nx5884, 
      nx5886, nx5888, nx5890, nx5892, nx5894, nx5896, nx5898, nx5900, nx5902, 
      nx5904, nx5906, nx5908, nx5910, nx5912, nx5914, nx5916, nx5918, nx5920, 
      nx5922, nx5924, nx5926, nx5928, nx5930, nx5932, nx5934, nx5936, nx5938, 
      nx5940, nx5942, nx5944, nx5946, nx5948, nx5950, nx5952, nx5954, nx5956, 
      nx5958, nx5960, nx5962, nx5964, nx5966, nx5968, nx5970, nx5972, nx5974, 
      nx5976, nx5978, nx5980, nx5982, nx5984, nx5986, nx5988, nx5990, nx5992, 
      nx5994, nx5996, nx5998, nx6000, nx6002, nx6004, nx6006, nx6008, nx6010, 
      nx6012, nx6014, nx6016, nx6018, nx6020, nx6022, nx6024, nx6026, nx6224, 
      nx6226, nx6228, nx6230, nx6232, nx6234, nx6236, nx6238, nx6240, nx6242, 
      nx6244, nx6246, nx6248, nx6250, nx6252, nx6254, nx6256, nx6258, nx6260, 
      nx6262, nx6264, nx6266, nx6268, nx6270, nx6272, nx6274, nx6276, nx6278, 
      nx6280, nx6282, nx6284, nx6286, nx6288, nx6290, nx6292, nx6294, nx6296, 
      nx6298, nx6300, nx6302, nx6304, nx6306, nx6308, nx6310, nx6312, nx6314, 
      nx6316, nx6318, nx6320, nx6322, nx6324, nx6326, nx6328, nx6330, nx6332, 
      nx6334, nx6336, nx6338, nx6340, nx6342, nx6344, nx6346, nx6348, nx6350, 
      nx6352, nx6354, nx6356, nx6358, nx6360, nx6362, nx6364, nx6366, nx6368, 
      nx6370, nx6372, nx6374, nx6376, nx6378, nx6380, nx6382, nx6384, nx6386, 
      nx6388, nx6390, nx6392, nx6394, nx6396, nx6398, nx6400, nx6402, nx6404, 
      nx6406, nx6408, nx6410, nx6412, nx6414, nx6416, nx6418, nx6420, nx6422, 
      nx6424, nx6426, nx6428, nx6430, nx6432, nx6434, nx6436, nx6438, nx6440, 
      nx6442, nx6444, nx6446, nx6448, nx6450, nx6452, nx6454, nx6456, nx6458, 
      nx6460, nx6462, nx6464, nx6466, nx6468, nx6470, nx6472, nx6474, nx6476, 
      nx6478, nx6480, nx6482, nx6484: std_logic ;

begin
   f0 : FC_nadder_32 port map ( aa(31)=>nx6026, aa(30)=>nx6026, aa(29)=>
      nx6024, aa(28)=>nx6024, aa(27)=>nx6024, aa(26)=>nx6022, aa(25)=>nx6022, 
      aa(24)=>nx6022, aa(23)=>nx6020, aa(22)=>nx6020, aa(21)=>nx6020, aa(20)
      =>nx6018, aa(19)=>nx6018, aa(18)=>nx6018, aa(17)=>nx6016, aa(16)=>
      nx6016, aa(15)=>nx6016, aa(14)=>op1_14, aa(13)=>op1_13, aa(12)=>op1_12, 
      aa(11)=>op1_11, aa(10)=>op1_10, aa(9)=>op1_9, aa(8)=>op1_8, aa(7)=>
      op1_7, aa(6)=>op1_6, aa(5)=>op1_5, aa(4)=>op1_4, aa(3)=>op1_3, aa(2)=>
      op1_2, aa(1)=>op1_1, aa(0)=>op1_0, bb(31)=>nx5780, bb(30)=>nx5778, 
      bb(29)=>nx5778, bb(28)=>nx5778, bb(27)=>nx5776, bb(26)=>nx5776, bb(25)
      =>nx5776, bb(24)=>nx5774, bb(23)=>nx5774, bb(22)=>nx5774, bb(21)=>
      nx5772, bb(20)=>nx5772, bb(19)=>nx5772, bb(18)=>nx5770, bb(17)=>nx5770, 
      bb(16)=>nx5770, bb(15)=>op2_0_15, bb(14)=>op2_0_14, bb(13)=>op2_0_13, 
      bb(12)=>op2_0_12, bb(11)=>op2_0_11, bb(10)=>op2_0_10, bb(9)=>op2_0_9, 
      bb(8)=>op2_0_8, bb(7)=>op2_0_7, bb(6)=>op2_0_6, bb(5)=>op2_0_5, bb(4)
      =>op2_0_4, bb(3)=>op2_0_3, bb(2)=>op2_0_2, bb(1)=>op2_0_1, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_0_31, ff(30)=>
      addout_0_30, ff(29)=>addout_0_29, ff(28)=>addout_0_28, ff(27)=>
      addout_0_27, ff(26)=>addout_0_26, ff(25)=>addout_0_25, ff(24)=>
      addout_0_24, ff(23)=>addout_0_23, ff(22)=>addout_0_22, ff(21)=>
      addout_0_21, ff(20)=>addout_0_20, ff(19)=>addout_0_19, ff(18)=>
      addout_0_18, ff(17)=>addout_0_17, ff(16)=>addout_0_16, ff(15)=>
      addout_0_15, ff(14)=>addout_0_14, ff(13)=>addout_0_13, ff(12)=>
      addout_0_12, ff(11)=>addout_0_11, ff(10)=>addout_0_10, ff(9)=>
      addout_0_9, ff(8)=>addout_0_8, ff(7)=>addout_0_7, ff(6)=>addout_0_6, 
      ff(5)=>addout_0_5, ff(4)=>addout_0_4, ff(3)=>addout_0_3, ff(2)=>
      addout_0_2, ff(1)=>addout_0_1, ff(0)=>addout_0_0);
   loop3_1_fx : FC_nadder_32 port map ( aa(31)=>addout_0_31, aa(30)=>
      addout_0_30, aa(29)=>addout_0_29, aa(28)=>addout_0_28, aa(27)=>
      addout_0_27, aa(26)=>addout_0_26, aa(25)=>addout_0_25, aa(24)=>
      addout_0_24, aa(23)=>addout_0_23, aa(22)=>addout_0_22, aa(21)=>
      addout_0_21, aa(20)=>addout_0_20, aa(19)=>addout_0_19, aa(18)=>
      addout_0_18, aa(17)=>addout_0_17, aa(16)=>addout_0_16, aa(15)=>
      addout_0_15, aa(14)=>addout_0_14, aa(13)=>addout_0_13, aa(12)=>
      addout_0_12, aa(11)=>addout_0_11, aa(10)=>addout_0_10, aa(9)=>
      addout_0_9, aa(8)=>addout_0_8, aa(7)=>addout_0_7, aa(6)=>addout_0_6, 
      aa(5)=>addout_0_5, aa(4)=>addout_0_4, aa(3)=>addout_0_3, aa(2)=>
      addout_0_2, aa(1)=>addout_0_1, aa(0)=>addout_0_0, bb(31)=>nx5792, 
      bb(30)=>nx5792, bb(29)=>nx5792, bb(28)=>nx5790, bb(27)=>nx5790, bb(26)
      =>nx5790, bb(25)=>nx5788, bb(24)=>nx5788, bb(23)=>nx5788, bb(22)=>
      nx5786, bb(21)=>nx5786, bb(20)=>nx5786, bb(19)=>nx5784, bb(18)=>nx5784, 
      bb(17)=>nx5784, bb(16)=>op2_1_16, bb(15)=>op2_1_15, bb(14)=>op2_1_14, 
      bb(13)=>op2_1_13, bb(12)=>op2_1_12, bb(11)=>op2_1_11, bb(10)=>op2_1_10, 
      bb(9)=>op2_1_9, bb(8)=>op2_1_8, bb(7)=>op2_1_7, bb(6)=>op2_1_6, bb(5)
      =>op2_1_5, bb(4)=>op2_1_4, bb(3)=>op2_1_3, bb(2)=>op2_1_2, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_1_31, ff(30)=>addout_1_30, ff(29)=>addout_1_29, ff(28)=>
      addout_1_28, ff(27)=>addout_1_27, ff(26)=>addout_1_26, ff(25)=>
      addout_1_25, ff(24)=>addout_1_24, ff(23)=>addout_1_23, ff(22)=>
      addout_1_22, ff(21)=>addout_1_21, ff(20)=>addout_1_20, ff(19)=>
      addout_1_19, ff(18)=>addout_1_18, ff(17)=>addout_1_17, ff(16)=>
      addout_1_16, ff(15)=>addout_1_15, ff(14)=>addout_1_14, ff(13)=>
      addout_1_13, ff(12)=>addout_1_12, ff(11)=>addout_1_11, ff(10)=>
      addout_1_10, ff(9)=>addout_1_9, ff(8)=>addout_1_8, ff(7)=>addout_1_7, 
      ff(6)=>addout_1_6, ff(5)=>addout_1_5, ff(4)=>addout_1_4, ff(3)=>
      addout_1_3, ff(2)=>addout_1_2, ff(1)=>addout_1_1, ff(0)=>addout_1_0);
   loop3_2_fx : FC_nadder_32 port map ( aa(31)=>addout_1_31, aa(30)=>
      addout_1_30, aa(29)=>addout_1_29, aa(28)=>addout_1_28, aa(27)=>
      addout_1_27, aa(26)=>addout_1_26, aa(25)=>addout_1_25, aa(24)=>
      addout_1_24, aa(23)=>addout_1_23, aa(22)=>addout_1_22, aa(21)=>
      addout_1_21, aa(20)=>addout_1_20, aa(19)=>addout_1_19, aa(18)=>
      addout_1_18, aa(17)=>addout_1_17, aa(16)=>addout_1_16, aa(15)=>
      addout_1_15, aa(14)=>addout_1_14, aa(13)=>addout_1_13, aa(12)=>
      addout_1_12, aa(11)=>addout_1_11, aa(10)=>addout_1_10, aa(9)=>
      addout_1_9, aa(8)=>addout_1_8, aa(7)=>addout_1_7, aa(6)=>addout_1_6, 
      aa(5)=>addout_1_5, aa(4)=>addout_1_4, aa(3)=>addout_1_3, aa(2)=>
      addout_1_2, aa(1)=>addout_1_1, aa(0)=>addout_1_0, bb(31)=>nx5804, 
      bb(30)=>nx5804, bb(29)=>nx5802, bb(28)=>nx5802, bb(27)=>nx5802, bb(26)
      =>nx5800, bb(25)=>nx5800, bb(24)=>nx5800, bb(23)=>nx5798, bb(22)=>
      nx5798, bb(21)=>nx5798, bb(20)=>nx5796, bb(19)=>nx5796, bb(18)=>nx5796, 
      bb(17)=>op2_2_17, bb(16)=>op2_2_16, bb(15)=>op2_2_15, bb(14)=>op2_2_14, 
      bb(13)=>op2_2_13, bb(12)=>op2_2_12, bb(11)=>op2_2_11, bb(10)=>op2_2_10, 
      bb(9)=>op2_2_9, bb(8)=>op2_2_8, bb(7)=>op2_2_7, bb(6)=>op2_2_6, bb(5)
      =>op2_2_5, bb(4)=>op2_2_4, bb(3)=>op2_2_3, bb(2)=>addout_31_31, bb(1)
      =>addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_2_31, ff(30)=>addout_2_30, ff(29)=>addout_2_29, ff(28)=>
      addout_2_28, ff(27)=>addout_2_27, ff(26)=>addout_2_26, ff(25)=>
      addout_2_25, ff(24)=>addout_2_24, ff(23)=>addout_2_23, ff(22)=>
      addout_2_22, ff(21)=>addout_2_21, ff(20)=>addout_2_20, ff(19)=>
      addout_2_19, ff(18)=>addout_2_18, ff(17)=>addout_2_17, ff(16)=>
      addout_2_16, ff(15)=>addout_2_15, ff(14)=>addout_2_14, ff(13)=>
      addout_2_13, ff(12)=>addout_2_12, ff(11)=>addout_2_11, ff(10)=>
      addout_2_10, ff(9)=>addout_2_9, ff(8)=>addout_2_8, ff(7)=>addout_2_7, 
      ff(6)=>addout_2_6, ff(5)=>addout_2_5, ff(4)=>addout_2_4, ff(3)=>
      addout_2_3, ff(2)=>addout_2_2, ff(1)=>addout_2_1, ff(0)=>addout_2_0);
   loop3_3_fx : FC_nadder_32 port map ( aa(31)=>addout_2_31, aa(30)=>
      addout_2_30, aa(29)=>addout_2_29, aa(28)=>addout_2_28, aa(27)=>
      addout_2_27, aa(26)=>addout_2_26, aa(25)=>addout_2_25, aa(24)=>
      addout_2_24, aa(23)=>addout_2_23, aa(22)=>addout_2_22, aa(21)=>
      addout_2_21, aa(20)=>addout_2_20, aa(19)=>addout_2_19, aa(18)=>
      addout_2_18, aa(17)=>addout_2_17, aa(16)=>addout_2_16, aa(15)=>
      addout_2_15, aa(14)=>addout_2_14, aa(13)=>addout_2_13, aa(12)=>
      addout_2_12, aa(11)=>addout_2_11, aa(10)=>addout_2_10, aa(9)=>
      addout_2_9, aa(8)=>addout_2_8, aa(7)=>addout_2_7, aa(6)=>addout_2_6, 
      aa(5)=>addout_2_5, aa(4)=>addout_2_4, aa(3)=>addout_2_3, aa(2)=>
      addout_2_2, aa(1)=>addout_2_1, aa(0)=>addout_2_0, bb(31)=>nx5816, 
      bb(30)=>nx5814, bb(29)=>nx5814, bb(28)=>nx5814, bb(27)=>nx5812, bb(26)
      =>nx5812, bb(25)=>nx5812, bb(24)=>nx5810, bb(23)=>nx5810, bb(22)=>
      nx5810, bb(21)=>nx5808, bb(20)=>nx5808, bb(19)=>nx5808, bb(18)=>
      op2_3_18, bb(17)=>op2_3_17, bb(16)=>op2_3_16, bb(15)=>op2_3_15, bb(14)
      =>op2_3_14, bb(13)=>op2_3_13, bb(12)=>op2_3_12, bb(11)=>op2_3_11, 
      bb(10)=>op2_3_10, bb(9)=>op2_3_9, bb(8)=>op2_3_8, bb(7)=>op2_3_7, 
      bb(6)=>op2_3_6, bb(5)=>op2_3_5, bb(4)=>op2_3_4, bb(3)=>addout_31_31, 
      bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>addout_31_31, c_cin=>
      addout_31_31, ff(31)=>addout_3_31, ff(30)=>addout_3_30, ff(29)=>
      addout_3_29, ff(28)=>addout_3_28, ff(27)=>addout_3_27, ff(26)=>
      addout_3_26, ff(25)=>addout_3_25, ff(24)=>addout_3_24, ff(23)=>
      addout_3_23, ff(22)=>addout_3_22, ff(21)=>addout_3_21, ff(20)=>
      addout_3_20, ff(19)=>addout_3_19, ff(18)=>addout_3_18, ff(17)=>
      addout_3_17, ff(16)=>addout_3_16, ff(15)=>addout_3_15, ff(14)=>
      addout_3_14, ff(13)=>addout_3_13, ff(12)=>addout_3_12, ff(11)=>
      addout_3_11, ff(10)=>addout_3_10, ff(9)=>addout_3_9, ff(8)=>addout_3_8, 
      ff(7)=>addout_3_7, ff(6)=>addout_3_6, ff(5)=>addout_3_5, ff(4)=>
      addout_3_4, ff(3)=>addout_3_3, ff(2)=>addout_3_2, ff(1)=>addout_3_1, 
      ff(0)=>addout_3_0);
   loop3_4_fx : FC_nadder_32 port map ( aa(31)=>addout_3_31, aa(30)=>
      addout_3_30, aa(29)=>addout_3_29, aa(28)=>addout_3_28, aa(27)=>
      addout_3_27, aa(26)=>addout_3_26, aa(25)=>addout_3_25, aa(24)=>
      addout_3_24, aa(23)=>addout_3_23, aa(22)=>addout_3_22, aa(21)=>
      addout_3_21, aa(20)=>addout_3_20, aa(19)=>addout_3_19, aa(18)=>
      addout_3_18, aa(17)=>addout_3_17, aa(16)=>addout_3_16, aa(15)=>
      addout_3_15, aa(14)=>addout_3_14, aa(13)=>addout_3_13, aa(12)=>
      addout_3_12, aa(11)=>addout_3_11, aa(10)=>addout_3_10, aa(9)=>
      addout_3_9, aa(8)=>addout_3_8, aa(7)=>addout_3_7, aa(6)=>addout_3_6, 
      aa(5)=>addout_3_5, aa(4)=>addout_3_4, aa(3)=>addout_3_3, aa(2)=>
      addout_3_2, aa(1)=>addout_3_1, aa(0)=>addout_3_0, bb(31)=>nx5826, 
      bb(30)=>nx5826, bb(29)=>nx5826, bb(28)=>nx5824, bb(27)=>nx5824, bb(26)
      =>nx5824, bb(25)=>nx5822, bb(24)=>nx5822, bb(23)=>nx5822, bb(22)=>
      nx5820, bb(21)=>nx5820, bb(20)=>nx5820, bb(19)=>op2_4_19, bb(18)=>
      op2_4_18, bb(17)=>op2_4_17, bb(16)=>op2_4_16, bb(15)=>op2_4_15, bb(14)
      =>op2_4_14, bb(13)=>op2_4_13, bb(12)=>op2_4_12, bb(11)=>op2_4_11, 
      bb(10)=>op2_4_10, bb(9)=>op2_4_9, bb(8)=>op2_4_8, bb(7)=>op2_4_7, 
      bb(6)=>op2_4_6, bb(5)=>op2_4_5, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_4_31, ff(30)=>
      addout_4_30, ff(29)=>addout_4_29, ff(28)=>addout_4_28, ff(27)=>
      addout_4_27, ff(26)=>addout_4_26, ff(25)=>addout_4_25, ff(24)=>
      addout_4_24, ff(23)=>addout_4_23, ff(22)=>addout_4_22, ff(21)=>
      addout_4_21, ff(20)=>addout_4_20, ff(19)=>addout_4_19, ff(18)=>
      addout_4_18, ff(17)=>addout_4_17, ff(16)=>addout_4_16, ff(15)=>
      addout_4_15, ff(14)=>addout_4_14, ff(13)=>addout_4_13, ff(12)=>
      addout_4_12, ff(11)=>addout_4_11, ff(10)=>addout_4_10, ff(9)=>
      addout_4_9, ff(8)=>addout_4_8, ff(7)=>addout_4_7, ff(6)=>addout_4_6, 
      ff(5)=>addout_4_5, ff(4)=>addout_4_4, ff(3)=>addout_4_3, ff(2)=>
      addout_4_2, ff(1)=>addout_4_1, ff(0)=>addout_4_0);
   loop3_5_fx : FC_nadder_32 port map ( aa(31)=>addout_4_31, aa(30)=>
      addout_4_30, aa(29)=>addout_4_29, aa(28)=>addout_4_28, aa(27)=>
      addout_4_27, aa(26)=>addout_4_26, aa(25)=>addout_4_25, aa(24)=>
      addout_4_24, aa(23)=>addout_4_23, aa(22)=>addout_4_22, aa(21)=>
      addout_4_21, aa(20)=>addout_4_20, aa(19)=>addout_4_19, aa(18)=>
      addout_4_18, aa(17)=>addout_4_17, aa(16)=>addout_4_16, aa(15)=>
      addout_4_15, aa(14)=>addout_4_14, aa(13)=>addout_4_13, aa(12)=>
      addout_4_12, aa(11)=>addout_4_11, aa(10)=>addout_4_10, aa(9)=>
      addout_4_9, aa(8)=>addout_4_8, aa(7)=>addout_4_7, aa(6)=>addout_4_6, 
      aa(5)=>addout_4_5, aa(4)=>addout_4_4, aa(3)=>addout_4_3, aa(2)=>
      addout_4_2, aa(1)=>addout_4_1, aa(0)=>addout_4_0, bb(31)=>nx5836, 
      bb(30)=>nx5836, bb(29)=>nx5834, bb(28)=>nx5834, bb(27)=>nx5834, bb(26)
      =>nx5832, bb(25)=>nx5832, bb(24)=>nx5832, bb(23)=>nx5830, bb(22)=>
      nx5830, bb(21)=>nx5830, bb(20)=>op2_5_20, bb(19)=>op2_5_19, bb(18)=>
      op2_5_18, bb(17)=>op2_5_17, bb(16)=>op2_5_16, bb(15)=>op2_5_15, bb(14)
      =>op2_5_14, bb(13)=>op2_5_13, bb(12)=>op2_5_12, bb(11)=>op2_5_11, 
      bb(10)=>op2_5_10, bb(9)=>op2_5_9, bb(8)=>op2_5_8, bb(7)=>op2_5_7, 
      bb(6)=>op2_5_6, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_5_31, ff(30)=>
      addout_5_30, ff(29)=>addout_5_29, ff(28)=>addout_5_28, ff(27)=>
      addout_5_27, ff(26)=>addout_5_26, ff(25)=>addout_5_25, ff(24)=>
      addout_5_24, ff(23)=>addout_5_23, ff(22)=>addout_5_22, ff(21)=>
      addout_5_21, ff(20)=>addout_5_20, ff(19)=>addout_5_19, ff(18)=>
      addout_5_18, ff(17)=>addout_5_17, ff(16)=>addout_5_16, ff(15)=>
      addout_5_15, ff(14)=>addout_5_14, ff(13)=>addout_5_13, ff(12)=>
      addout_5_12, ff(11)=>addout_5_11, ff(10)=>addout_5_10, ff(9)=>
      addout_5_9, ff(8)=>addout_5_8, ff(7)=>addout_5_7, ff(6)=>addout_5_6, 
      ff(5)=>addout_5_5, ff(4)=>addout_5_4, ff(3)=>addout_5_3, ff(2)=>
      addout_5_2, ff(1)=>addout_5_1, ff(0)=>addout_5_0);
   loop3_6_fx : FC_nadder_32 port map ( aa(31)=>addout_5_31, aa(30)=>
      addout_5_30, aa(29)=>addout_5_29, aa(28)=>addout_5_28, aa(27)=>
      addout_5_27, aa(26)=>addout_5_26, aa(25)=>addout_5_25, aa(24)=>
      addout_5_24, aa(23)=>addout_5_23, aa(22)=>addout_5_22, aa(21)=>
      addout_5_21, aa(20)=>addout_5_20, aa(19)=>addout_5_19, aa(18)=>
      addout_5_18, aa(17)=>addout_5_17, aa(16)=>addout_5_16, aa(15)=>
      addout_5_15, aa(14)=>addout_5_14, aa(13)=>addout_5_13, aa(12)=>
      addout_5_12, aa(11)=>addout_5_11, aa(10)=>addout_5_10, aa(9)=>
      addout_5_9, aa(8)=>addout_5_8, aa(7)=>addout_5_7, aa(6)=>addout_5_6, 
      aa(5)=>addout_5_5, aa(4)=>addout_5_4, aa(3)=>addout_5_3, aa(2)=>
      addout_5_2, aa(1)=>addout_5_1, aa(0)=>addout_5_0, bb(31)=>nx5846, 
      bb(30)=>nx5844, bb(29)=>nx5844, bb(28)=>nx5844, bb(27)=>nx5842, bb(26)
      =>nx5842, bb(25)=>nx5842, bb(24)=>nx5840, bb(23)=>nx5840, bb(22)=>
      nx5840, bb(21)=>op2_6_21, bb(20)=>op2_6_20, bb(19)=>op2_6_19, bb(18)=>
      op2_6_18, bb(17)=>op2_6_17, bb(16)=>op2_6_16, bb(15)=>op2_6_15, bb(14)
      =>op2_6_14, bb(13)=>op2_6_13, bb(12)=>op2_6_12, bb(11)=>op2_6_11, 
      bb(10)=>op2_6_10, bb(9)=>op2_6_9, bb(8)=>op2_6_8, bb(7)=>op2_6_7, 
      bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_6_31, ff(30)=>
      addout_6_30, ff(29)=>addout_6_29, ff(28)=>addout_6_28, ff(27)=>
      addout_6_27, ff(26)=>addout_6_26, ff(25)=>addout_6_25, ff(24)=>
      addout_6_24, ff(23)=>addout_6_23, ff(22)=>addout_6_22, ff(21)=>
      addout_6_21, ff(20)=>addout_6_20, ff(19)=>addout_6_19, ff(18)=>
      addout_6_18, ff(17)=>addout_6_17, ff(16)=>addout_6_16, ff(15)=>
      addout_6_15, ff(14)=>addout_6_14, ff(13)=>addout_6_13, ff(12)=>
      addout_6_12, ff(11)=>addout_6_11, ff(10)=>addout_6_10, ff(9)=>
      addout_6_9, ff(8)=>addout_6_8, ff(7)=>addout_6_7, ff(6)=>addout_6_6, 
      ff(5)=>addout_6_5, ff(4)=>addout_6_4, ff(3)=>addout_6_3, ff(2)=>
      addout_6_2, ff(1)=>addout_6_1, ff(0)=>addout_6_0);
   loop3_7_fx : FC_nadder_32 port map ( aa(31)=>addout_6_31, aa(30)=>
      addout_6_30, aa(29)=>addout_6_29, aa(28)=>addout_6_28, aa(27)=>
      addout_6_27, aa(26)=>addout_6_26, aa(25)=>addout_6_25, aa(24)=>
      addout_6_24, aa(23)=>addout_6_23, aa(22)=>addout_6_22, aa(21)=>
      addout_6_21, aa(20)=>addout_6_20, aa(19)=>addout_6_19, aa(18)=>
      addout_6_18, aa(17)=>addout_6_17, aa(16)=>addout_6_16, aa(15)=>
      addout_6_15, aa(14)=>addout_6_14, aa(13)=>addout_6_13, aa(12)=>
      addout_6_12, aa(11)=>addout_6_11, aa(10)=>addout_6_10, aa(9)=>
      addout_6_9, aa(8)=>addout_6_8, aa(7)=>addout_6_7, aa(6)=>addout_6_6, 
      aa(5)=>addout_6_5, aa(4)=>addout_6_4, aa(3)=>addout_6_3, aa(2)=>
      addout_6_2, aa(1)=>addout_6_1, aa(0)=>addout_6_0, bb(31)=>nx5854, 
      bb(30)=>nx5854, bb(29)=>nx5854, bb(28)=>nx5852, bb(27)=>nx5852, bb(26)
      =>nx5852, bb(25)=>nx5850, bb(24)=>nx5850, bb(23)=>nx5850, bb(22)=>
      op2_7_22, bb(21)=>op2_7_21, bb(20)=>op2_7_20, bb(19)=>op2_7_19, bb(18)
      =>op2_7_18, bb(17)=>op2_7_17, bb(16)=>op2_7_16, bb(15)=>op2_7_15, 
      bb(14)=>op2_7_14, bb(13)=>op2_7_13, bb(12)=>op2_7_12, bb(11)=>op2_7_11, 
      bb(10)=>op2_7_10, bb(9)=>op2_7_9, bb(8)=>op2_7_8, bb(7)=>addout_31_31, 
      bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_7_31, ff(30)=>
      addout_7_30, ff(29)=>addout_7_29, ff(28)=>addout_7_28, ff(27)=>
      addout_7_27, ff(26)=>addout_7_26, ff(25)=>addout_7_25, ff(24)=>
      addout_7_24, ff(23)=>addout_7_23, ff(22)=>addout_7_22, ff(21)=>
      addout_7_21, ff(20)=>addout_7_20, ff(19)=>addout_7_19, ff(18)=>
      addout_7_18, ff(17)=>addout_7_17, ff(16)=>addout_7_16, ff(15)=>
      addout_7_15, ff(14)=>addout_7_14, ff(13)=>addout_7_13, ff(12)=>
      addout_7_12, ff(11)=>addout_7_11, ff(10)=>addout_7_10, ff(9)=>
      addout_7_9, ff(8)=>addout_7_8, ff(7)=>addout_7_7, ff(6)=>addout_7_6, 
      ff(5)=>addout_7_5, ff(4)=>addout_7_4, ff(3)=>addout_7_3, ff(2)=>
      addout_7_2, ff(1)=>addout_7_1, ff(0)=>addout_7_0);
   loop3_8_fx : FC_nadder_32 port map ( aa(31)=>addout_7_31, aa(30)=>
      addout_7_30, aa(29)=>addout_7_29, aa(28)=>addout_7_28, aa(27)=>
      addout_7_27, aa(26)=>addout_7_26, aa(25)=>addout_7_25, aa(24)=>
      addout_7_24, aa(23)=>addout_7_23, aa(22)=>addout_7_22, aa(21)=>
      addout_7_21, aa(20)=>addout_7_20, aa(19)=>addout_7_19, aa(18)=>
      addout_7_18, aa(17)=>addout_7_17, aa(16)=>addout_7_16, aa(15)=>
      addout_7_15, aa(14)=>addout_7_14, aa(13)=>addout_7_13, aa(12)=>
      addout_7_12, aa(11)=>addout_7_11, aa(10)=>addout_7_10, aa(9)=>
      addout_7_9, aa(8)=>addout_7_8, aa(7)=>addout_7_7, aa(6)=>addout_7_6, 
      aa(5)=>addout_7_5, aa(4)=>addout_7_4, aa(3)=>addout_7_3, aa(2)=>
      addout_7_2, aa(1)=>addout_7_1, aa(0)=>addout_7_0, bb(31)=>nx5862, 
      bb(30)=>nx5862, bb(29)=>nx5860, bb(28)=>nx5860, bb(27)=>nx5860, bb(26)
      =>nx5858, bb(25)=>nx5858, bb(24)=>nx5858, bb(23)=>op2_8_23, bb(22)=>
      op2_8_22, bb(21)=>op2_8_21, bb(20)=>op2_8_20, bb(19)=>op2_8_19, bb(18)
      =>op2_8_18, bb(17)=>op2_8_17, bb(16)=>op2_8_16, bb(15)=>op2_8_15, 
      bb(14)=>op2_8_14, bb(13)=>op2_8_13, bb(12)=>op2_8_12, bb(11)=>op2_8_11, 
      bb(10)=>op2_8_10, bb(9)=>op2_8_9, bb(8)=>addout_31_31, bb(7)=>
      addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_8_31, ff(30)=>addout_8_30, ff(29)=>addout_8_29, ff(28)=>
      addout_8_28, ff(27)=>addout_8_27, ff(26)=>addout_8_26, ff(25)=>
      addout_8_25, ff(24)=>addout_8_24, ff(23)=>addout_8_23, ff(22)=>
      addout_8_22, ff(21)=>addout_8_21, ff(20)=>addout_8_20, ff(19)=>
      addout_8_19, ff(18)=>addout_8_18, ff(17)=>addout_8_17, ff(16)=>
      addout_8_16, ff(15)=>addout_8_15, ff(14)=>addout_8_14, ff(13)=>
      addout_8_13, ff(12)=>addout_8_12, ff(11)=>addout_8_11, ff(10)=>
      addout_8_10, ff(9)=>addout_8_9, ff(8)=>addout_8_8, ff(7)=>addout_8_7, 
      ff(6)=>addout_8_6, ff(5)=>addout_8_5, ff(4)=>addout_8_4, ff(3)=>
      addout_8_3, ff(2)=>addout_8_2, ff(1)=>addout_8_1, ff(0)=>addout_8_0);
   loop3_9_fx : FC_nadder_32 port map ( aa(31)=>addout_8_31, aa(30)=>
      addout_8_30, aa(29)=>addout_8_29, aa(28)=>addout_8_28, aa(27)=>
      addout_8_27, aa(26)=>addout_8_26, aa(25)=>addout_8_25, aa(24)=>
      addout_8_24, aa(23)=>addout_8_23, aa(22)=>addout_8_22, aa(21)=>
      addout_8_21, aa(20)=>addout_8_20, aa(19)=>addout_8_19, aa(18)=>
      addout_8_18, aa(17)=>addout_8_17, aa(16)=>addout_8_16, aa(15)=>
      addout_8_15, aa(14)=>addout_8_14, aa(13)=>addout_8_13, aa(12)=>
      addout_8_12, aa(11)=>addout_8_11, aa(10)=>addout_8_10, aa(9)=>
      addout_8_9, aa(8)=>addout_8_8, aa(7)=>addout_8_7, aa(6)=>addout_8_6, 
      aa(5)=>addout_8_5, aa(4)=>addout_8_4, aa(3)=>addout_8_3, aa(2)=>
      addout_8_2, aa(1)=>addout_8_1, aa(0)=>addout_8_0, bb(31)=>nx5870, 
      bb(30)=>nx5868, bb(29)=>nx5868, bb(28)=>nx5868, bb(27)=>nx5866, bb(26)
      =>nx5866, bb(25)=>nx5866, bb(24)=>op2_9_24, bb(23)=>op2_9_23, bb(22)=>
      op2_9_22, bb(21)=>op2_9_21, bb(20)=>op2_9_20, bb(19)=>op2_9_19, bb(18)
      =>op2_9_18, bb(17)=>op2_9_17, bb(16)=>op2_9_16, bb(15)=>op2_9_15, 
      bb(14)=>op2_9_14, bb(13)=>op2_9_13, bb(12)=>op2_9_12, bb(11)=>op2_9_11, 
      bb(10)=>op2_9_10, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>
      addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_9_31, ff(30)=>addout_9_30, ff(29)=>addout_9_29, ff(28)=>
      addout_9_28, ff(27)=>addout_9_27, ff(26)=>addout_9_26, ff(25)=>
      addout_9_25, ff(24)=>addout_9_24, ff(23)=>addout_9_23, ff(22)=>
      addout_9_22, ff(21)=>addout_9_21, ff(20)=>addout_9_20, ff(19)=>
      addout_9_19, ff(18)=>addout_9_18, ff(17)=>addout_9_17, ff(16)=>
      addout_9_16, ff(15)=>addout_9_15, ff(14)=>addout_9_14, ff(13)=>
      addout_9_13, ff(12)=>addout_9_12, ff(11)=>addout_9_11, ff(10)=>
      addout_9_10, ff(9)=>addout_9_9, ff(8)=>addout_9_8, ff(7)=>addout_9_7, 
      ff(6)=>addout_9_6, ff(5)=>addout_9_5, ff(4)=>addout_9_4, ff(3)=>
      addout_9_3, ff(2)=>addout_9_2, ff(1)=>addout_9_1, ff(0)=>addout_9_0);
   loop3_10_fx : FC_nadder_32 port map ( aa(31)=>addout_9_31, aa(30)=>
      addout_9_30, aa(29)=>addout_9_29, aa(28)=>addout_9_28, aa(27)=>
      addout_9_27, aa(26)=>addout_9_26, aa(25)=>addout_9_25, aa(24)=>
      addout_9_24, aa(23)=>addout_9_23, aa(22)=>addout_9_22, aa(21)=>
      addout_9_21, aa(20)=>addout_9_20, aa(19)=>addout_9_19, aa(18)=>
      addout_9_18, aa(17)=>addout_9_17, aa(16)=>addout_9_16, aa(15)=>
      addout_9_15, aa(14)=>addout_9_14, aa(13)=>addout_9_13, aa(12)=>
      addout_9_12, aa(11)=>addout_9_11, aa(10)=>addout_9_10, aa(9)=>
      addout_9_9, aa(8)=>addout_9_8, aa(7)=>addout_9_7, aa(6)=>addout_9_6, 
      aa(5)=>addout_9_5, aa(4)=>addout_9_4, aa(3)=>addout_9_3, aa(2)=>
      addout_9_2, aa(1)=>addout_9_1, aa(0)=>addout_9_0, bb(31)=>nx5874, 
      bb(30)=>nx5874, bb(29)=>nx5874, bb(28)=>nx5872, bb(27)=>nx5872, bb(26)
      =>nx5872, bb(25)=>op2_10_25, bb(24)=>op2_10_24, bb(23)=>op2_10_23, 
      bb(22)=>op2_10_22, bb(21)=>op2_10_21, bb(20)=>op2_10_20, bb(19)=>
      op2_10_19, bb(18)=>op2_10_18, bb(17)=>op2_10_17, bb(16)=>op2_10_16, 
      bb(15)=>op2_10_15, bb(14)=>op2_10_14, bb(13)=>op2_10_13, bb(12)=>
      op2_10_12, bb(11)=>op2_10_11, bb(10)=>addout_31_31, bb(9)=>
      addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_10_31, ff(30)=>
      addout_10_30, ff(29)=>addout_10_29, ff(28)=>addout_10_28, ff(27)=>
      addout_10_27, ff(26)=>addout_10_26, ff(25)=>addout_10_25, ff(24)=>
      addout_10_24, ff(23)=>addout_10_23, ff(22)=>addout_10_22, ff(21)=>
      addout_10_21, ff(20)=>addout_10_20, ff(19)=>addout_10_19, ff(18)=>
      addout_10_18, ff(17)=>addout_10_17, ff(16)=>addout_10_16, ff(15)=>
      addout_10_15, ff(14)=>addout_10_14, ff(13)=>addout_10_13, ff(12)=>
      addout_10_12, ff(11)=>addout_10_11, ff(10)=>addout_10_10, ff(9)=>
      addout_10_9, ff(8)=>addout_10_8, ff(7)=>addout_10_7, ff(6)=>
      addout_10_6, ff(5)=>addout_10_5, ff(4)=>addout_10_4, ff(3)=>
      addout_10_3, ff(2)=>addout_10_2, ff(1)=>addout_10_1, ff(0)=>
      addout_10_0);
   loop3_11_fx : FC_nadder_32 port map ( aa(31)=>addout_10_31, aa(30)=>
      addout_10_30, aa(29)=>addout_10_29, aa(28)=>addout_10_28, aa(27)=>
      addout_10_27, aa(26)=>addout_10_26, aa(25)=>addout_10_25, aa(24)=>
      addout_10_24, aa(23)=>addout_10_23, aa(22)=>addout_10_22, aa(21)=>
      addout_10_21, aa(20)=>addout_10_20, aa(19)=>addout_10_19, aa(18)=>
      addout_10_18, aa(17)=>addout_10_17, aa(16)=>addout_10_16, aa(15)=>
      addout_10_15, aa(14)=>addout_10_14, aa(13)=>addout_10_13, aa(12)=>
      addout_10_12, aa(11)=>addout_10_11, aa(10)=>addout_10_10, aa(9)=>
      addout_10_9, aa(8)=>addout_10_8, aa(7)=>addout_10_7, aa(6)=>
      addout_10_6, aa(5)=>addout_10_5, aa(4)=>addout_10_4, aa(3)=>
      addout_10_3, aa(2)=>addout_10_2, aa(1)=>addout_10_1, aa(0)=>
      addout_10_0, bb(31)=>nx5878, bb(30)=>nx5878, bb(29)=>nx5876, bb(28)=>
      nx5876, bb(27)=>nx5876, bb(26)=>op2_11_26, bb(25)=>op2_11_25, bb(24)=>
      op2_11_24, bb(23)=>op2_11_23, bb(22)=>op2_11_22, bb(21)=>op2_11_21, 
      bb(20)=>op2_11_20, bb(19)=>op2_11_19, bb(18)=>op2_11_18, bb(17)=>
      op2_11_17, bb(16)=>op2_11_16, bb(15)=>op2_11_15, bb(14)=>op2_11_14, 
      bb(13)=>op2_11_13, bb(12)=>op2_11_12, bb(11)=>addout_31_31, bb(10)=>
      addout_31_31, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>
      addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_11_31, ff(30)=>addout_11_30, ff(29)=>addout_11_29, ff(28)=>
      addout_11_28, ff(27)=>addout_11_27, ff(26)=>addout_11_26, ff(25)=>
      addout_11_25, ff(24)=>addout_11_24, ff(23)=>addout_11_23, ff(22)=>
      addout_11_22, ff(21)=>addout_11_21, ff(20)=>addout_11_20, ff(19)=>
      addout_11_19, ff(18)=>addout_11_18, ff(17)=>addout_11_17, ff(16)=>
      addout_11_16, ff(15)=>addout_11_15, ff(14)=>addout_11_14, ff(13)=>
      addout_11_13, ff(12)=>addout_11_12, ff(11)=>addout_11_11, ff(10)=>
      addout_11_10, ff(9)=>addout_11_9, ff(8)=>addout_11_8, ff(7)=>
      addout_11_7, ff(6)=>addout_11_6, ff(5)=>addout_11_5, ff(4)=>
      addout_11_4, ff(3)=>addout_11_3, ff(2)=>addout_11_2, ff(1)=>
      addout_11_1, ff(0)=>addout_11_0);
   loop3_12_fx : FC_nadder_32 port map ( aa(31)=>addout_11_31, aa(30)=>
      addout_11_30, aa(29)=>addout_11_29, aa(28)=>addout_11_28, aa(27)=>
      addout_11_27, aa(26)=>addout_11_26, aa(25)=>addout_11_25, aa(24)=>
      addout_11_24, aa(23)=>addout_11_23, aa(22)=>addout_11_22, aa(21)=>
      addout_11_21, aa(20)=>addout_11_20, aa(19)=>addout_11_19, aa(18)=>
      addout_11_18, aa(17)=>addout_11_17, aa(16)=>addout_11_16, aa(15)=>
      addout_11_15, aa(14)=>addout_11_14, aa(13)=>addout_11_13, aa(12)=>
      addout_11_12, aa(11)=>addout_11_11, aa(10)=>addout_11_10, aa(9)=>
      addout_11_9, aa(8)=>addout_11_8, aa(7)=>addout_11_7, aa(6)=>
      addout_11_6, aa(5)=>addout_11_5, aa(4)=>addout_11_4, aa(3)=>
      addout_11_3, aa(2)=>addout_11_2, aa(1)=>addout_11_1, aa(0)=>
      addout_11_0, bb(31)=>nx5882, bb(30)=>nx5880, bb(29)=>nx5880, bb(28)=>
      nx5880, bb(27)=>op2_12_27, bb(26)=>op2_12_26, bb(25)=>op2_12_25, 
      bb(24)=>op2_12_24, bb(23)=>op2_12_23, bb(22)=>op2_12_22, bb(21)=>
      op2_12_21, bb(20)=>op2_12_20, bb(19)=>op2_12_19, bb(18)=>op2_12_18, 
      bb(17)=>op2_12_17, bb(16)=>op2_12_16, bb(15)=>op2_12_15, bb(14)=>
      op2_12_14, bb(13)=>op2_12_13, bb(12)=>addout_31_31, bb(11)=>
      addout_31_31, bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)=>
      addout_31_31, bb(7)=>addout_31_31, bb(6)=>addout_31_31, bb(5)=>
      addout_31_31, bb(4)=>addout_31_31, bb(3)=>addout_31_31, bb(2)=>
      addout_31_31, bb(1)=>addout_31_31, bb(0)=>addout_31_31, c_cin=>
      addout_31_31, ff(31)=>addout_12_31, ff(30)=>addout_12_30, ff(29)=>
      addout_12_29, ff(28)=>addout_12_28, ff(27)=>addout_12_27, ff(26)=>
      addout_12_26, ff(25)=>addout_12_25, ff(24)=>addout_12_24, ff(23)=>
      addout_12_23, ff(22)=>addout_12_22, ff(21)=>addout_12_21, ff(20)=>
      addout_12_20, ff(19)=>addout_12_19, ff(18)=>addout_12_18, ff(17)=>
      addout_12_17, ff(16)=>addout_12_16, ff(15)=>addout_12_15, ff(14)=>
      addout_12_14, ff(13)=>addout_12_13, ff(12)=>addout_12_12, ff(11)=>
      addout_12_11, ff(10)=>addout_12_10, ff(9)=>addout_12_9, ff(8)=>
      addout_12_8, ff(7)=>addout_12_7, ff(6)=>addout_12_6, ff(5)=>
      addout_12_5, ff(4)=>addout_12_4, ff(3)=>addout_12_3, ff(2)=>
      addout_12_2, ff(1)=>addout_12_1, ff(0)=>addout_12_0);
   loop3_13_fx : FC_nadder_32 port map ( aa(31)=>addout_12_31, aa(30)=>
      addout_12_30, aa(29)=>addout_12_29, aa(28)=>addout_12_28, aa(27)=>
      addout_12_27, aa(26)=>addout_12_26, aa(25)=>addout_12_25, aa(24)=>
      addout_12_24, aa(23)=>addout_12_23, aa(22)=>addout_12_22, aa(21)=>
      addout_12_21, aa(20)=>addout_12_20, aa(19)=>addout_12_19, aa(18)=>
      addout_12_18, aa(17)=>addout_12_17, aa(16)=>addout_12_16, aa(15)=>
      addout_12_15, aa(14)=>addout_12_14, aa(13)=>addout_12_13, aa(12)=>
      addout_12_12, aa(11)=>addout_12_11, aa(10)=>addout_12_10, aa(9)=>
      addout_12_9, aa(8)=>addout_12_8, aa(7)=>addout_12_7, aa(6)=>
      addout_12_6, aa(5)=>addout_12_5, aa(4)=>addout_12_4, aa(3)=>
      addout_12_3, aa(2)=>addout_12_2, aa(1)=>addout_12_1, aa(0)=>
      addout_12_0, bb(31)=>nx6480, bb(30)=>nx6480, bb(29)=>nx6480, bb(28)=>
      op2_13_28, bb(27)=>op2_13_27, bb(26)=>op2_13_26, bb(25)=>op2_13_25, 
      bb(24)=>op2_13_24, bb(23)=>op2_13_23, bb(22)=>op2_13_22, bb(21)=>
      op2_13_21, bb(20)=>op2_13_20, bb(19)=>op2_13_19, bb(18)=>op2_13_18, 
      bb(17)=>op2_13_17, bb(16)=>op2_13_16, bb(15)=>op2_13_15, bb(14)=>
      op2_13_14, bb(13)=>addout_31_31, bb(12)=>addout_31_31, bb(11)=>
      addout_31_31, bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)=>
      addout_31_31, bb(7)=>addout_31_31, bb(6)=>addout_31_31, bb(5)=>
      addout_31_31, bb(4)=>addout_31_31, bb(3)=>addout_31_31, bb(2)=>
      addout_31_31, bb(1)=>addout_31_31, bb(0)=>addout_31_31, c_cin=>
      addout_31_31, ff(31)=>addout_13_31, ff(30)=>addout_13_30, ff(29)=>
      addout_13_29, ff(28)=>addout_13_28, ff(27)=>addout_13_27, ff(26)=>
      addout_13_26, ff(25)=>addout_13_25, ff(24)=>addout_13_24, ff(23)=>
      addout_13_23, ff(22)=>addout_13_22, ff(21)=>addout_13_21, ff(20)=>
      addout_13_20, ff(19)=>addout_13_19, ff(18)=>addout_13_18, ff(17)=>
      addout_13_17, ff(16)=>addout_13_16, ff(15)=>addout_13_15, ff(14)=>
      addout_13_14, ff(13)=>addout_13_13, ff(12)=>addout_13_12, ff(11)=>
      addout_13_11, ff(10)=>addout_13_10, ff(9)=>addout_13_9, ff(8)=>
      addout_13_8, ff(7)=>addout_13_7, ff(6)=>addout_13_6, ff(5)=>
      addout_13_5, ff(4)=>addout_13_4, ff(3)=>addout_13_3, ff(2)=>
      addout_13_2, ff(1)=>addout_13_1, ff(0)=>addout_13_0);
   loop3_14_fx : FC_nadder_32 port map ( aa(31)=>addout_13_31, aa(30)=>
      addout_13_30, aa(29)=>addout_13_29, aa(28)=>addout_13_28, aa(27)=>
      addout_13_27, aa(26)=>addout_13_26, aa(25)=>addout_13_25, aa(24)=>
      addout_13_24, aa(23)=>addout_13_23, aa(22)=>addout_13_22, aa(21)=>
      addout_13_21, aa(20)=>addout_13_20, aa(19)=>addout_13_19, aa(18)=>
      addout_13_18, aa(17)=>addout_13_17, aa(16)=>addout_13_16, aa(15)=>
      addout_13_15, aa(14)=>addout_13_14, aa(13)=>addout_13_13, aa(12)=>
      addout_13_12, aa(11)=>addout_13_11, aa(10)=>addout_13_10, aa(9)=>
      addout_13_9, aa(8)=>addout_13_8, aa(7)=>addout_13_7, aa(6)=>
      addout_13_6, aa(5)=>addout_13_5, aa(4)=>addout_13_4, aa(3)=>
      addout_13_3, aa(2)=>addout_13_2, aa(1)=>addout_13_1, aa(0)=>
      addout_13_0, bb(31)=>nx6482, bb(30)=>nx6482, bb(29)=>nx6484, bb(28)=>
      nx5884, bb(27)=>nx5888, bb(26)=>nx5892, bb(25)=>nx5898, bb(24)=>nx5906, 
      bb(23)=>nx5914, bb(22)=>nx5922, bb(21)=>nx5932, bb(20)=>nx5942, bb(19)
      =>nx5952, bb(18)=>nx5964, bb(17)=>nx5976, bb(16)=>nx5988, bb(15)=>
      nx6002, bb(14)=>addout_31_31, bb(13)=>addout_31_31, bb(12)=>
      addout_31_31, bb(11)=>addout_31_31, bb(10)=>addout_31_31, bb(9)=>
      addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_14_31, ff(30)=>
      addout_14_30, ff(29)=>addout_14_29, ff(28)=>addout_14_28, ff(27)=>
      addout_14_27, ff(26)=>addout_14_26, ff(25)=>addout_14_25, ff(24)=>
      addout_14_24, ff(23)=>addout_14_23, ff(22)=>addout_14_22, ff(21)=>
      addout_14_21, ff(20)=>addout_14_20, ff(19)=>addout_14_19, ff(18)=>
      addout_14_18, ff(17)=>addout_14_17, ff(16)=>addout_14_16, ff(15)=>
      addout_14_15, ff(14)=>addout_14_14, ff(13)=>addout_14_13, ff(12)=>
      addout_14_12, ff(11)=>addout_14_11, ff(10)=>addout_14_10, ff(9)=>
      addout_14_9, ff(8)=>addout_14_8, ff(7)=>addout_14_7, ff(6)=>
      addout_14_6, ff(5)=>addout_14_5, ff(4)=>addout_14_4, ff(3)=>
      addout_14_3, ff(2)=>addout_14_2, ff(1)=>addout_14_1, ff(0)=>
      addout_14_0);
   loop3_15_fx : FC_nadder_32 port map ( aa(31)=>addout_14_31, aa(30)=>
      addout_14_30, aa(29)=>addout_14_29, aa(28)=>addout_14_28, aa(27)=>
      addout_14_27, aa(26)=>addout_14_26, aa(25)=>addout_14_25, aa(24)=>
      addout_14_24, aa(23)=>addout_14_23, aa(22)=>addout_14_22, aa(21)=>
      addout_14_21, aa(20)=>addout_14_20, aa(19)=>addout_14_19, aa(18)=>
      addout_14_18, aa(17)=>addout_14_17, aa(16)=>addout_14_16, aa(15)=>
      addout_14_15, aa(14)=>addout_14_14, aa(13)=>addout_14_13, aa(12)=>
      addout_14_12, aa(11)=>addout_14_11, aa(10)=>addout_14_10, aa(9)=>
      addout_14_9, aa(8)=>addout_14_8, aa(7)=>addout_14_7, aa(6)=>
      addout_14_6, aa(5)=>addout_14_5, aa(4)=>addout_14_4, aa(3)=>
      addout_14_3, aa(2)=>addout_14_2, aa(1)=>addout_14_1, aa(0)=>
      addout_14_0, bb(31)=>nx6482, bb(30)=>nx6484, bb(29)=>nx5884, bb(28)=>
      nx5888, bb(27)=>nx5892, bb(26)=>nx5898, bb(25)=>nx5906, bb(24)=>nx5914, 
      bb(23)=>nx5922, bb(22)=>nx5932, bb(21)=>nx5942, bb(20)=>nx5952, bb(19)
      =>nx5964, bb(18)=>nx5976, bb(17)=>nx5988, bb(16)=>nx6002, bb(15)=>
      addout_31_31, bb(14)=>addout_31_31, bb(13)=>addout_31_31, bb(12)=>
      addout_31_31, bb(11)=>addout_31_31, bb(10)=>addout_31_31, bb(9)=>
      addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_15_31, ff(30)=>
      addout_15_30, ff(29)=>addout_15_29, ff(28)=>addout_15_28, ff(27)=>
      addout_15_27, ff(26)=>addout_15_26, ff(25)=>addout_15_25, ff(24)=>
      addout_15_24, ff(23)=>addout_15_23, ff(22)=>addout_15_22, ff(21)=>
      addout_15_21, ff(20)=>addout_15_20, ff(19)=>addout_15_19, ff(18)=>
      addout_15_18, ff(17)=>addout_15_17, ff(16)=>addout_15_16, ff(15)=>
      addout_15_15, ff(14)=>addout_15_14, ff(13)=>addout_15_13, ff(12)=>
      addout_15_12, ff(11)=>addout_15_11, ff(10)=>addout_15_10, ff(9)=>
      addout_15_9, ff(8)=>addout_15_8, ff(7)=>addout_15_7, ff(6)=>
      addout_15_6, ff(5)=>addout_15_5, ff(4)=>addout_15_4, ff(3)=>
      addout_15_3, ff(2)=>addout_15_2, ff(1)=>addout_15_1, ff(0)=>
      addout_15_0);
   loop3_16_fx : FC_nadder_32 port map ( aa(31)=>addout_15_31, aa(30)=>
      addout_15_30, aa(29)=>addout_15_29, aa(28)=>addout_15_28, aa(27)=>
      addout_15_27, aa(26)=>addout_15_26, aa(25)=>addout_15_25, aa(24)=>
      addout_15_24, aa(23)=>addout_15_23, aa(22)=>addout_15_22, aa(21)=>
      addout_15_21, aa(20)=>addout_15_20, aa(19)=>addout_15_19, aa(18)=>
      addout_15_18, aa(17)=>addout_15_17, aa(16)=>addout_15_16, aa(15)=>
      addout_15_15, aa(14)=>addout_15_14, aa(13)=>addout_15_13, aa(12)=>
      addout_15_12, aa(11)=>addout_15_11, aa(10)=>addout_15_10, aa(9)=>
      addout_15_9, aa(8)=>addout_15_8, aa(7)=>addout_15_7, aa(6)=>
      addout_15_6, aa(5)=>addout_15_5, aa(4)=>addout_15_4, aa(3)=>
      addout_15_3, aa(2)=>addout_15_2, aa(1)=>addout_15_1, aa(0)=>
      addout_15_0, bb(31)=>nx6484, bb(30)=>nx5884, bb(29)=>nx5888, bb(28)=>
      nx5892, bb(27)=>nx5898, bb(26)=>nx5906, bb(25)=>nx5914, bb(24)=>nx5922, 
      bb(23)=>nx5932, bb(22)=>nx5942, bb(21)=>nx5952, bb(20)=>nx5964, bb(19)
      =>nx5976, bb(18)=>nx5988, bb(17)=>nx6002, bb(16)=>addout_31_31, bb(15)
      =>addout_31_31, bb(14)=>addout_31_31, bb(13)=>addout_31_31, bb(12)=>
      addout_31_31, bb(11)=>addout_31_31, bb(10)=>addout_31_31, bb(9)=>
      addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_16_31, ff(30)=>
      addout_16_30, ff(29)=>addout_16_29, ff(28)=>addout_16_28, ff(27)=>
      addout_16_27, ff(26)=>addout_16_26, ff(25)=>addout_16_25, ff(24)=>
      addout_16_24, ff(23)=>addout_16_23, ff(22)=>addout_16_22, ff(21)=>
      addout_16_21, ff(20)=>addout_16_20, ff(19)=>addout_16_19, ff(18)=>
      addout_16_18, ff(17)=>addout_16_17, ff(16)=>addout_16_16, ff(15)=>
      addout_16_15, ff(14)=>addout_16_14, ff(13)=>addout_16_13, ff(12)=>
      addout_16_12, ff(11)=>addout_16_11, ff(10)=>addout_16_10, ff(9)=>
      addout_16_9, ff(8)=>addout_16_8, ff(7)=>addout_16_7, ff(6)=>
      addout_16_6, ff(5)=>addout_16_5, ff(4)=>addout_16_4, ff(3)=>
      addout_16_3, ff(2)=>addout_16_2, ff(1)=>addout_16_1, ff(0)=>
      addout_16_0);
   loop3_17_fx : FC_nadder_32 port map ( aa(31)=>addout_16_31, aa(30)=>
      addout_16_30, aa(29)=>addout_16_29, aa(28)=>addout_16_28, aa(27)=>
      addout_16_27, aa(26)=>addout_16_26, aa(25)=>addout_16_25, aa(24)=>
      addout_16_24, aa(23)=>addout_16_23, aa(22)=>addout_16_22, aa(21)=>
      addout_16_21, aa(20)=>addout_16_20, aa(19)=>addout_16_19, aa(18)=>
      addout_16_18, aa(17)=>addout_16_17, aa(16)=>addout_16_16, aa(15)=>
      addout_16_15, aa(14)=>addout_16_14, aa(13)=>addout_16_13, aa(12)=>
      addout_16_12, aa(11)=>addout_16_11, aa(10)=>addout_16_10, aa(9)=>
      addout_16_9, aa(8)=>addout_16_8, aa(7)=>addout_16_7, aa(6)=>
      addout_16_6, aa(5)=>addout_16_5, aa(4)=>addout_16_4, aa(3)=>
      addout_16_3, aa(2)=>addout_16_2, aa(1)=>addout_16_1, aa(0)=>
      addout_16_0, bb(31)=>nx5886, bb(30)=>nx5890, bb(29)=>nx5894, bb(28)=>
      nx5900, bb(27)=>nx5908, bb(26)=>nx5916, bb(25)=>nx5924, bb(24)=>nx5934, 
      bb(23)=>nx5944, bb(22)=>nx5954, bb(21)=>nx5966, bb(20)=>nx5978, bb(19)
      =>nx5990, bb(18)=>nx6004, bb(17)=>addout_31_31, bb(16)=>addout_31_31, 
      bb(15)=>addout_31_31, bb(14)=>addout_31_31, bb(13)=>addout_31_31, 
      bb(12)=>addout_31_31, bb(11)=>addout_31_31, bb(10)=>addout_31_31, 
      bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_17_31, ff(30)=>
      addout_17_30, ff(29)=>addout_17_29, ff(28)=>addout_17_28, ff(27)=>
      addout_17_27, ff(26)=>addout_17_26, ff(25)=>addout_17_25, ff(24)=>
      addout_17_24, ff(23)=>addout_17_23, ff(22)=>addout_17_22, ff(21)=>
      addout_17_21, ff(20)=>addout_17_20, ff(19)=>addout_17_19, ff(18)=>
      addout_17_18, ff(17)=>addout_17_17, ff(16)=>addout_17_16, ff(15)=>
      addout_17_15, ff(14)=>addout_17_14, ff(13)=>addout_17_13, ff(12)=>
      addout_17_12, ff(11)=>addout_17_11, ff(10)=>addout_17_10, ff(9)=>
      addout_17_9, ff(8)=>addout_17_8, ff(7)=>addout_17_7, ff(6)=>
      addout_17_6, ff(5)=>addout_17_5, ff(4)=>addout_17_4, ff(3)=>
      addout_17_3, ff(2)=>addout_17_2, ff(1)=>addout_17_1, ff(0)=>
      addout_17_0);
   loop3_18_fx : FC_nadder_32 port map ( aa(31)=>addout_17_31, aa(30)=>
      addout_17_30, aa(29)=>addout_17_29, aa(28)=>addout_17_28, aa(27)=>
      addout_17_27, aa(26)=>addout_17_26, aa(25)=>addout_17_25, aa(24)=>
      addout_17_24, aa(23)=>addout_17_23, aa(22)=>addout_17_22, aa(21)=>
      addout_17_21, aa(20)=>addout_17_20, aa(19)=>addout_17_19, aa(18)=>
      addout_17_18, aa(17)=>addout_17_17, aa(16)=>addout_17_16, aa(15)=>
      addout_17_15, aa(14)=>addout_17_14, aa(13)=>addout_17_13, aa(12)=>
      addout_17_12, aa(11)=>addout_17_11, aa(10)=>addout_17_10, aa(9)=>
      addout_17_9, aa(8)=>addout_17_8, aa(7)=>addout_17_7, aa(6)=>
      addout_17_6, aa(5)=>addout_17_5, aa(4)=>addout_17_4, aa(3)=>
      addout_17_3, aa(2)=>addout_17_2, aa(1)=>addout_17_1, aa(0)=>
      addout_17_0, bb(31)=>nx5890, bb(30)=>nx5894, bb(29)=>nx5900, bb(28)=>
      nx5908, bb(27)=>nx5916, bb(26)=>nx5924, bb(25)=>nx5934, bb(24)=>nx5944, 
      bb(23)=>nx5954, bb(22)=>nx5966, bb(21)=>nx5978, bb(20)=>nx5990, bb(19)
      =>nx6004, bb(18)=>addout_31_31, bb(17)=>addout_31_31, bb(16)=>
      addout_31_31, bb(15)=>addout_31_31, bb(14)=>addout_31_31, bb(13)=>
      addout_31_31, bb(12)=>addout_31_31, bb(11)=>addout_31_31, bb(10)=>
      addout_31_31, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>
      addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_18_31, ff(30)=>addout_18_30, ff(29)=>addout_18_29, ff(28)=>
      addout_18_28, ff(27)=>addout_18_27, ff(26)=>addout_18_26, ff(25)=>
      addout_18_25, ff(24)=>addout_18_24, ff(23)=>addout_18_23, ff(22)=>
      addout_18_22, ff(21)=>addout_18_21, ff(20)=>addout_18_20, ff(19)=>
      addout_18_19, ff(18)=>addout_18_18, ff(17)=>addout_18_17, ff(16)=>
      addout_18_16, ff(15)=>addout_18_15, ff(14)=>addout_18_14, ff(13)=>
      addout_18_13, ff(12)=>addout_18_12, ff(11)=>addout_18_11, ff(10)=>
      addout_18_10, ff(9)=>addout_18_9, ff(8)=>addout_18_8, ff(7)=>
      addout_18_7, ff(6)=>addout_18_6, ff(5)=>addout_18_5, ff(4)=>
      addout_18_4, ff(3)=>addout_18_3, ff(2)=>addout_18_2, ff(1)=>
      addout_18_1, ff(0)=>addout_18_0);
   loop3_19_fx : FC_nadder_32 port map ( aa(31)=>addout_18_31, aa(30)=>
      addout_18_30, aa(29)=>addout_18_29, aa(28)=>addout_18_28, aa(27)=>
      addout_18_27, aa(26)=>addout_18_26, aa(25)=>addout_18_25, aa(24)=>
      addout_18_24, aa(23)=>addout_18_23, aa(22)=>addout_18_22, aa(21)=>
      addout_18_21, aa(20)=>addout_18_20, aa(19)=>addout_18_19, aa(18)=>
      addout_18_18, aa(17)=>addout_18_17, aa(16)=>addout_18_16, aa(15)=>
      addout_18_15, aa(14)=>addout_18_14, aa(13)=>addout_18_13, aa(12)=>
      addout_18_12, aa(11)=>addout_18_11, aa(10)=>addout_18_10, aa(9)=>
      addout_18_9, aa(8)=>addout_18_8, aa(7)=>addout_18_7, aa(6)=>
      addout_18_6, aa(5)=>addout_18_5, aa(4)=>addout_18_4, aa(3)=>
      addout_18_3, aa(2)=>addout_18_2, aa(1)=>addout_18_1, aa(0)=>
      addout_18_0, bb(31)=>nx5894, bb(30)=>nx5900, bb(29)=>nx5908, bb(28)=>
      nx5916, bb(27)=>nx5924, bb(26)=>nx5934, bb(25)=>nx5944, bb(24)=>nx5954, 
      bb(23)=>nx5966, bb(22)=>nx5978, bb(21)=>nx5990, bb(20)=>nx6004, bb(19)
      =>addout_31_31, bb(18)=>addout_31_31, bb(17)=>addout_31_31, bb(16)=>
      addout_31_31, bb(15)=>addout_31_31, bb(14)=>addout_31_31, bb(13)=>
      addout_31_31, bb(12)=>addout_31_31, bb(11)=>addout_31_31, bb(10)=>
      addout_31_31, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>
      addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_19_31, ff(30)=>addout_19_30, ff(29)=>addout_19_29, ff(28)=>
      addout_19_28, ff(27)=>addout_19_27, ff(26)=>addout_19_26, ff(25)=>
      addout_19_25, ff(24)=>addout_19_24, ff(23)=>addout_19_23, ff(22)=>
      addout_19_22, ff(21)=>addout_19_21, ff(20)=>addout_19_20, ff(19)=>
      addout_19_19, ff(18)=>addout_19_18, ff(17)=>addout_19_17, ff(16)=>
      addout_19_16, ff(15)=>addout_19_15, ff(14)=>addout_19_14, ff(13)=>
      addout_19_13, ff(12)=>addout_19_12, ff(11)=>addout_19_11, ff(10)=>
      addout_19_10, ff(9)=>addout_19_9, ff(8)=>addout_19_8, ff(7)=>
      addout_19_7, ff(6)=>addout_19_6, ff(5)=>addout_19_5, ff(4)=>
      addout_19_4, ff(3)=>addout_19_3, ff(2)=>addout_19_2, ff(1)=>
      addout_19_1, ff(0)=>addout_19_0);
   loop3_20_fx : FC_nadder_32 port map ( aa(31)=>addout_19_31, aa(30)=>
      addout_19_30, aa(29)=>addout_19_29, aa(28)=>addout_19_28, aa(27)=>
      addout_19_27, aa(26)=>addout_19_26, aa(25)=>addout_19_25, aa(24)=>
      addout_19_24, aa(23)=>addout_19_23, aa(22)=>addout_19_22, aa(21)=>
      addout_19_21, aa(20)=>addout_19_20, aa(19)=>addout_19_19, aa(18)=>
      addout_19_18, aa(17)=>addout_19_17, aa(16)=>addout_19_16, aa(15)=>
      addout_19_15, aa(14)=>addout_19_14, aa(13)=>addout_19_13, aa(12)=>
      addout_19_12, aa(11)=>addout_19_11, aa(10)=>addout_19_10, aa(9)=>
      addout_19_9, aa(8)=>addout_19_8, aa(7)=>addout_19_7, aa(6)=>
      addout_19_6, aa(5)=>addout_19_5, aa(4)=>addout_19_4, aa(3)=>
      addout_19_3, aa(2)=>addout_19_2, aa(1)=>addout_19_1, aa(0)=>
      addout_19_0, bb(31)=>nx5902, bb(30)=>nx5910, bb(29)=>nx5918, bb(28)=>
      nx5926, bb(27)=>nx5936, bb(26)=>nx5946, bb(25)=>nx5956, bb(24)=>nx5968, 
      bb(23)=>nx5980, bb(22)=>nx5992, bb(21)=>nx6006, bb(20)=>addout_31_31, 
      bb(19)=>addout_31_31, bb(18)=>addout_31_31, bb(17)=>addout_31_31, 
      bb(16)=>addout_31_31, bb(15)=>addout_31_31, bb(14)=>addout_31_31, 
      bb(13)=>addout_31_31, bb(12)=>addout_31_31, bb(11)=>addout_31_31, 
      bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)
      =>addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_20_31, ff(30)=>addout_20_30, ff(29)=>addout_20_29, ff(28)=>
      addout_20_28, ff(27)=>addout_20_27, ff(26)=>addout_20_26, ff(25)=>
      addout_20_25, ff(24)=>addout_20_24, ff(23)=>addout_20_23, ff(22)=>
      addout_20_22, ff(21)=>addout_20_21, ff(20)=>addout_20_20, ff(19)=>
      addout_20_19, ff(18)=>addout_20_18, ff(17)=>addout_20_17, ff(16)=>
      addout_20_16, ff(15)=>addout_20_15, ff(14)=>addout_20_14, ff(13)=>
      addout_20_13, ff(12)=>addout_20_12, ff(11)=>addout_20_11, ff(10)=>
      addout_20_10, ff(9)=>addout_20_9, ff(8)=>addout_20_8, ff(7)=>
      addout_20_7, ff(6)=>addout_20_6, ff(5)=>addout_20_5, ff(4)=>
      addout_20_4, ff(3)=>addout_20_3, ff(2)=>addout_20_2, ff(1)=>
      addout_20_1, ff(0)=>addout_20_0);
   loop3_21_fx : FC_nadder_32 port map ( aa(31)=>addout_20_31, aa(30)=>
      addout_20_30, aa(29)=>addout_20_29, aa(28)=>addout_20_28, aa(27)=>
      addout_20_27, aa(26)=>addout_20_26, aa(25)=>addout_20_25, aa(24)=>
      addout_20_24, aa(23)=>addout_20_23, aa(22)=>addout_20_22, aa(21)=>
      addout_20_21, aa(20)=>addout_20_20, aa(19)=>addout_20_19, aa(18)=>
      addout_20_18, aa(17)=>addout_20_17, aa(16)=>addout_20_16, aa(15)=>
      addout_20_15, aa(14)=>addout_20_14, aa(13)=>addout_20_13, aa(12)=>
      addout_20_12, aa(11)=>addout_20_11, aa(10)=>addout_20_10, aa(9)=>
      addout_20_9, aa(8)=>addout_20_8, aa(7)=>addout_20_7, aa(6)=>
      addout_20_6, aa(5)=>addout_20_5, aa(4)=>addout_20_4, aa(3)=>
      addout_20_3, aa(2)=>addout_20_2, aa(1)=>addout_20_1, aa(0)=>
      addout_20_0, bb(31)=>nx5910, bb(30)=>nx5918, bb(29)=>nx5926, bb(28)=>
      nx5936, bb(27)=>nx5946, bb(26)=>nx5956, bb(25)=>nx5968, bb(24)=>nx5980, 
      bb(23)=>nx5992, bb(22)=>nx6006, bb(21)=>addout_31_31, bb(20)=>
      addout_31_31, bb(19)=>addout_31_31, bb(18)=>addout_31_31, bb(17)=>
      addout_31_31, bb(16)=>addout_31_31, bb(15)=>addout_31_31, bb(14)=>
      addout_31_31, bb(13)=>addout_31_31, bb(12)=>addout_31_31, bb(11)=>
      addout_31_31, bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)=>
      addout_31_31, bb(7)=>addout_31_31, bb(6)=>addout_31_31, bb(5)=>
      addout_31_31, bb(4)=>addout_31_31, bb(3)=>addout_31_31, bb(2)=>
      addout_31_31, bb(1)=>addout_31_31, bb(0)=>addout_31_31, c_cin=>
      addout_31_31, ff(31)=>addout_21_31, ff(30)=>addout_21_30, ff(29)=>
      addout_21_29, ff(28)=>addout_21_28, ff(27)=>addout_21_27, ff(26)=>
      addout_21_26, ff(25)=>addout_21_25, ff(24)=>addout_21_24, ff(23)=>
      addout_21_23, ff(22)=>addout_21_22, ff(21)=>addout_21_21, ff(20)=>
      addout_21_20, ff(19)=>addout_21_19, ff(18)=>addout_21_18, ff(17)=>
      addout_21_17, ff(16)=>addout_21_16, ff(15)=>addout_21_15, ff(14)=>
      addout_21_14, ff(13)=>addout_21_13, ff(12)=>addout_21_12, ff(11)=>
      addout_21_11, ff(10)=>addout_21_10, ff(9)=>addout_21_9, ff(8)=>
      addout_21_8, ff(7)=>addout_21_7, ff(6)=>addout_21_6, ff(5)=>
      addout_21_5, ff(4)=>addout_21_4, ff(3)=>addout_21_3, ff(2)=>
      addout_21_2, ff(1)=>addout_21_1, ff(0)=>addout_21_0);
   loop3_22_fx : FC_nadder_32 port map ( aa(31)=>addout_21_31, aa(30)=>
      addout_21_30, aa(29)=>addout_21_29, aa(28)=>addout_21_28, aa(27)=>
      addout_21_27, aa(26)=>addout_21_26, aa(25)=>addout_21_25, aa(24)=>
      addout_21_24, aa(23)=>addout_21_23, aa(22)=>addout_21_22, aa(21)=>
      addout_21_21, aa(20)=>addout_21_20, aa(19)=>addout_21_19, aa(18)=>
      addout_21_18, aa(17)=>addout_21_17, aa(16)=>addout_21_16, aa(15)=>
      addout_21_15, aa(14)=>addout_21_14, aa(13)=>addout_21_13, aa(12)=>
      addout_21_12, aa(11)=>addout_21_11, aa(10)=>addout_21_10, aa(9)=>
      addout_21_9, aa(8)=>addout_21_8, aa(7)=>addout_21_7, aa(6)=>
      addout_21_6, aa(5)=>addout_21_5, aa(4)=>addout_21_4, aa(3)=>
      addout_21_3, aa(2)=>addout_21_2, aa(1)=>addout_21_1, aa(0)=>
      addout_21_0, bb(31)=>nx5918, bb(30)=>nx5926, bb(29)=>nx5936, bb(28)=>
      nx5946, bb(27)=>nx5956, bb(26)=>nx5968, bb(25)=>nx5980, bb(24)=>nx5992, 
      bb(23)=>nx6006, bb(22)=>addout_31_31, bb(21)=>addout_31_31, bb(20)=>
      addout_31_31, bb(19)=>addout_31_31, bb(18)=>addout_31_31, bb(17)=>
      addout_31_31, bb(16)=>addout_31_31, bb(15)=>addout_31_31, bb(14)=>
      addout_31_31, bb(13)=>addout_31_31, bb(12)=>addout_31_31, bb(11)=>
      addout_31_31, bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)=>
      addout_31_31, bb(7)=>addout_31_31, bb(6)=>addout_31_31, bb(5)=>
      addout_31_31, bb(4)=>addout_31_31, bb(3)=>addout_31_31, bb(2)=>
      addout_31_31, bb(1)=>addout_31_31, bb(0)=>addout_31_31, c_cin=>
      addout_31_31, ff(31)=>addout_22_31, ff(30)=>addout_22_30, ff(29)=>
      addout_22_29, ff(28)=>addout_22_28, ff(27)=>addout_22_27, ff(26)=>
      addout_22_26, ff(25)=>addout_22_25, ff(24)=>addout_22_24, ff(23)=>
      addout_22_23, ff(22)=>addout_22_22, ff(21)=>addout_22_21, ff(20)=>
      addout_22_20, ff(19)=>addout_22_19, ff(18)=>addout_22_18, ff(17)=>
      addout_22_17, ff(16)=>addout_22_16, ff(15)=>addout_22_15, ff(14)=>
      addout_22_14, ff(13)=>addout_22_13, ff(12)=>addout_22_12, ff(11)=>
      addout_22_11, ff(10)=>addout_22_10, ff(9)=>addout_22_9, ff(8)=>
      addout_22_8, ff(7)=>addout_22_7, ff(6)=>addout_22_6, ff(5)=>
      addout_22_5, ff(4)=>addout_22_4, ff(3)=>addout_22_3, ff(2)=>
      addout_22_2, ff(1)=>addout_22_1, ff(0)=>addout_22_0);
   loop3_23_fx : FC_nadder_32 port map ( aa(31)=>addout_22_31, aa(30)=>
      addout_22_30, aa(29)=>addout_22_29, aa(28)=>addout_22_28, aa(27)=>
      addout_22_27, aa(26)=>addout_22_26, aa(25)=>addout_22_25, aa(24)=>
      addout_22_24, aa(23)=>addout_22_23, aa(22)=>addout_22_22, aa(21)=>
      addout_22_21, aa(20)=>addout_22_20, aa(19)=>addout_22_19, aa(18)=>
      addout_22_18, aa(17)=>addout_22_17, aa(16)=>addout_22_16, aa(15)=>
      addout_22_15, aa(14)=>addout_22_14, aa(13)=>addout_22_13, aa(12)=>
      addout_22_12, aa(11)=>addout_22_11, aa(10)=>addout_22_10, aa(9)=>
      addout_22_9, aa(8)=>addout_22_8, aa(7)=>addout_22_7, aa(6)=>
      addout_22_6, aa(5)=>addout_22_5, aa(4)=>addout_22_4, aa(3)=>
      addout_22_3, aa(2)=>addout_22_2, aa(1)=>addout_22_1, aa(0)=>
      addout_22_0, bb(31)=>nx5928, bb(30)=>nx5938, bb(29)=>nx5948, bb(28)=>
      nx5958, bb(27)=>nx5970, bb(26)=>nx5982, bb(25)=>nx5994, bb(24)=>nx6008, 
      bb(23)=>addout_31_31, bb(22)=>addout_31_31, bb(21)=>addout_31_31, 
      bb(20)=>addout_31_31, bb(19)=>addout_31_31, bb(18)=>addout_31_31, 
      bb(17)=>addout_31_31, bb(16)=>addout_31_31, bb(15)=>addout_31_31, 
      bb(14)=>addout_31_31, bb(13)=>addout_31_31, bb(12)=>addout_31_31, 
      bb(11)=>addout_31_31, bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)
      =>addout_31_31, bb(7)=>addout_31_31, bb(6)=>addout_31_31, bb(5)=>
      addout_31_31, bb(4)=>addout_31_31, bb(3)=>addout_31_31, bb(2)=>
      addout_31_31, bb(1)=>addout_31_31, bb(0)=>addout_31_31, c_cin=>
      addout_31_31, ff(31)=>addout_23_31, ff(30)=>addout_23_30, ff(29)=>
      addout_23_29, ff(28)=>addout_23_28, ff(27)=>addout_23_27, ff(26)=>
      addout_23_26, ff(25)=>addout_23_25, ff(24)=>addout_23_24, ff(23)=>
      addout_23_23, ff(22)=>addout_23_22, ff(21)=>addout_23_21, ff(20)=>
      addout_23_20, ff(19)=>addout_23_19, ff(18)=>addout_23_18, ff(17)=>
      addout_23_17, ff(16)=>addout_23_16, ff(15)=>addout_23_15, ff(14)=>
      addout_23_14, ff(13)=>addout_23_13, ff(12)=>addout_23_12, ff(11)=>
      addout_23_11, ff(10)=>addout_23_10, ff(9)=>addout_23_9, ff(8)=>
      addout_23_8, ff(7)=>addout_23_7, ff(6)=>addout_23_6, ff(5)=>
      addout_23_5, ff(4)=>addout_23_4, ff(3)=>addout_23_3, ff(2)=>
      addout_23_2, ff(1)=>addout_23_1, ff(0)=>addout_23_0);
   loop3_24_fx : FC_nadder_32 port map ( aa(31)=>addout_23_31, aa(30)=>
      addout_23_30, aa(29)=>addout_23_29, aa(28)=>addout_23_28, aa(27)=>
      addout_23_27, aa(26)=>addout_23_26, aa(25)=>addout_23_25, aa(24)=>
      addout_23_24, aa(23)=>addout_23_23, aa(22)=>addout_23_22, aa(21)=>
      addout_23_21, aa(20)=>addout_23_20, aa(19)=>addout_23_19, aa(18)=>
      addout_23_18, aa(17)=>addout_23_17, aa(16)=>addout_23_16, aa(15)=>
      addout_23_15, aa(14)=>addout_23_14, aa(13)=>addout_23_13, aa(12)=>
      addout_23_12, aa(11)=>addout_23_11, aa(10)=>addout_23_10, aa(9)=>
      addout_23_9, aa(8)=>addout_23_8, aa(7)=>addout_23_7, aa(6)=>
      addout_23_6, aa(5)=>addout_23_5, aa(4)=>addout_23_4, aa(3)=>
      addout_23_3, aa(2)=>addout_23_2, aa(1)=>addout_23_1, aa(0)=>
      addout_23_0, bb(31)=>nx5938, bb(30)=>nx5948, bb(29)=>nx5958, bb(28)=>
      nx5970, bb(27)=>nx5982, bb(26)=>nx5994, bb(25)=>nx6008, bb(24)=>
      addout_31_31, bb(23)=>addout_31_31, bb(22)=>addout_31_31, bb(21)=>
      addout_31_31, bb(20)=>addout_31_31, bb(19)=>addout_31_31, bb(18)=>
      addout_31_31, bb(17)=>addout_31_31, bb(16)=>addout_31_31, bb(15)=>
      addout_31_31, bb(14)=>addout_31_31, bb(13)=>addout_31_31, bb(12)=>
      addout_31_31, bb(11)=>addout_31_31, bb(10)=>addout_31_31, bb(9)=>
      addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_24_31, ff(30)=>
      addout_24_30, ff(29)=>addout_24_29, ff(28)=>addout_24_28, ff(27)=>
      addout_24_27, ff(26)=>addout_24_26, ff(25)=>addout_24_25, ff(24)=>
      addout_24_24, ff(23)=>addout_24_23, ff(22)=>addout_24_22, ff(21)=>
      addout_24_21, ff(20)=>addout_24_20, ff(19)=>addout_24_19, ff(18)=>
      addout_24_18, ff(17)=>addout_24_17, ff(16)=>addout_24_16, ff(15)=>
      addout_24_15, ff(14)=>addout_24_14, ff(13)=>addout_24_13, ff(12)=>
      addout_24_12, ff(11)=>addout_24_11, ff(10)=>addout_24_10, ff(9)=>
      addout_24_9, ff(8)=>addout_24_8, ff(7)=>addout_24_7, ff(6)=>
      addout_24_6, ff(5)=>addout_24_5, ff(4)=>addout_24_4, ff(3)=>
      addout_24_3, ff(2)=>addout_24_2, ff(1)=>addout_24_1, ff(0)=>
      addout_24_0);
   loop3_25_fx : FC_nadder_32 port map ( aa(31)=>addout_24_31, aa(30)=>
      addout_24_30, aa(29)=>addout_24_29, aa(28)=>addout_24_28, aa(27)=>
      addout_24_27, aa(26)=>addout_24_26, aa(25)=>addout_24_25, aa(24)=>
      addout_24_24, aa(23)=>addout_24_23, aa(22)=>addout_24_22, aa(21)=>
      addout_24_21, aa(20)=>addout_24_20, aa(19)=>addout_24_19, aa(18)=>
      addout_24_18, aa(17)=>addout_24_17, aa(16)=>addout_24_16, aa(15)=>
      addout_24_15, aa(14)=>addout_24_14, aa(13)=>addout_24_13, aa(12)=>
      addout_24_12, aa(11)=>addout_24_11, aa(10)=>addout_24_10, aa(9)=>
      addout_24_9, aa(8)=>addout_24_8, aa(7)=>addout_24_7, aa(6)=>
      addout_24_6, aa(5)=>addout_24_5, aa(4)=>addout_24_4, aa(3)=>
      addout_24_3, aa(2)=>addout_24_2, aa(1)=>addout_24_1, aa(0)=>
      addout_24_0, bb(31)=>nx5948, bb(30)=>nx5958, bb(29)=>nx5970, bb(28)=>
      nx5982, bb(27)=>nx5994, bb(26)=>nx6008, bb(25)=>addout_31_31, bb(24)=>
      addout_31_31, bb(23)=>addout_31_31, bb(22)=>addout_31_31, bb(21)=>
      addout_31_31, bb(20)=>addout_31_31, bb(19)=>addout_31_31, bb(18)=>
      addout_31_31, bb(17)=>addout_31_31, bb(16)=>addout_31_31, bb(15)=>
      addout_31_31, bb(14)=>addout_31_31, bb(13)=>addout_31_31, bb(12)=>
      addout_31_31, bb(11)=>addout_31_31, bb(10)=>addout_31_31, bb(9)=>
      addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_25_31, ff(30)=>
      addout_25_30, ff(29)=>addout_25_29, ff(28)=>addout_25_28, ff(27)=>
      addout_25_27, ff(26)=>addout_25_26, ff(25)=>addout_25_25, ff(24)=>
      addout_25_24, ff(23)=>addout_25_23, ff(22)=>addout_25_22, ff(21)=>
      addout_25_21, ff(20)=>addout_25_20, ff(19)=>addout_25_19, ff(18)=>
      addout_25_18, ff(17)=>addout_25_17, ff(16)=>addout_25_16, ff(15)=>
      addout_25_15, ff(14)=>addout_25_14, ff(13)=>addout_25_13, ff(12)=>
      addout_25_12, ff(11)=>addout_25_11, ff(10)=>addout_25_10, ff(9)=>
      addout_25_9, ff(8)=>addout_25_8, ff(7)=>addout_25_7, ff(6)=>
      addout_25_6, ff(5)=>addout_25_5, ff(4)=>addout_25_4, ff(3)=>
      addout_25_3, ff(2)=>addout_25_2, ff(1)=>addout_25_1, ff(0)=>
      addout_25_0);
   loop3_26_fx : FC_nadder_32 port map ( aa(31)=>addout_25_31, aa(30)=>
      addout_25_30, aa(29)=>addout_25_29, aa(28)=>addout_25_28, aa(27)=>
      addout_25_27, aa(26)=>addout_25_26, aa(25)=>addout_25_25, aa(24)=>
      addout_25_24, aa(23)=>addout_25_23, aa(22)=>addout_25_22, aa(21)=>
      addout_25_21, aa(20)=>addout_25_20, aa(19)=>addout_25_19, aa(18)=>
      addout_25_18, aa(17)=>addout_25_17, aa(16)=>addout_25_16, aa(15)=>
      addout_25_15, aa(14)=>addout_25_14, aa(13)=>addout_25_13, aa(12)=>
      addout_25_12, aa(11)=>addout_25_11, aa(10)=>addout_25_10, aa(9)=>
      addout_25_9, aa(8)=>addout_25_8, aa(7)=>addout_25_7, aa(6)=>
      addout_25_6, aa(5)=>addout_25_5, aa(4)=>addout_25_4, aa(3)=>
      addout_25_3, aa(2)=>addout_25_2, aa(1)=>addout_25_1, aa(0)=>
      addout_25_0, bb(31)=>nx5960, bb(30)=>nx5972, bb(29)=>nx5984, bb(28)=>
      nx5996, bb(27)=>nx6010, bb(26)=>addout_31_31, bb(25)=>addout_31_31, 
      bb(24)=>addout_31_31, bb(23)=>addout_31_31, bb(22)=>addout_31_31, 
      bb(21)=>addout_31_31, bb(20)=>addout_31_31, bb(19)=>addout_31_31, 
      bb(18)=>addout_31_31, bb(17)=>addout_31_31, bb(16)=>addout_31_31, 
      bb(15)=>addout_31_31, bb(14)=>addout_31_31, bb(13)=>addout_31_31, 
      bb(12)=>addout_31_31, bb(11)=>addout_31_31, bb(10)=>addout_31_31, 
      bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>addout_31_31, bb(6)=>
      addout_31_31, bb(5)=>addout_31_31, bb(4)=>addout_31_31, bb(3)=>
      addout_31_31, bb(2)=>addout_31_31, bb(1)=>addout_31_31, bb(0)=>
      addout_31_31, c_cin=>addout_31_31, ff(31)=>addout_26_31, ff(30)=>
      addout_26_30, ff(29)=>addout_26_29, ff(28)=>addout_26_28, ff(27)=>
      addout_26_27, ff(26)=>addout_26_26, ff(25)=>addout_26_25, ff(24)=>
      addout_26_24, ff(23)=>addout_26_23, ff(22)=>addout_26_22, ff(21)=>
      addout_26_21, ff(20)=>addout_26_20, ff(19)=>addout_26_19, ff(18)=>
      addout_26_18, ff(17)=>addout_26_17, ff(16)=>addout_26_16, ff(15)=>
      addout_26_15, ff(14)=>addout_26_14, ff(13)=>addout_26_13, ff(12)=>
      addout_26_12, ff(11)=>addout_26_11, ff(10)=>addout_26_10, ff(9)=>
      addout_26_9, ff(8)=>addout_26_8, ff(7)=>addout_26_7, ff(6)=>
      addout_26_6, ff(5)=>addout_26_5, ff(4)=>addout_26_4, ff(3)=>
      addout_26_3, ff(2)=>addout_26_2, ff(1)=>addout_26_1, ff(0)=>
      addout_26_0);
   loop3_27_fx : FC_nadder_32 port map ( aa(31)=>addout_26_31, aa(30)=>
      addout_26_30, aa(29)=>addout_26_29, aa(28)=>addout_26_28, aa(27)=>
      addout_26_27, aa(26)=>addout_26_26, aa(25)=>addout_26_25, aa(24)=>
      addout_26_24, aa(23)=>addout_26_23, aa(22)=>addout_26_22, aa(21)=>
      addout_26_21, aa(20)=>addout_26_20, aa(19)=>addout_26_19, aa(18)=>
      addout_26_18, aa(17)=>addout_26_17, aa(16)=>addout_26_16, aa(15)=>
      addout_26_15, aa(14)=>addout_26_14, aa(13)=>addout_26_13, aa(12)=>
      addout_26_12, aa(11)=>addout_26_11, aa(10)=>addout_26_10, aa(9)=>
      addout_26_9, aa(8)=>addout_26_8, aa(7)=>addout_26_7, aa(6)=>
      addout_26_6, aa(5)=>addout_26_5, aa(4)=>addout_26_4, aa(3)=>
      addout_26_3, aa(2)=>addout_26_2, aa(1)=>addout_26_1, aa(0)=>
      addout_26_0, bb(31)=>nx5972, bb(30)=>nx5984, bb(29)=>nx5996, bb(28)=>
      nx6010, bb(27)=>addout_31_31, bb(26)=>addout_31_31, bb(25)=>
      addout_31_31, bb(24)=>addout_31_31, bb(23)=>addout_31_31, bb(22)=>
      addout_31_31, bb(21)=>addout_31_31, bb(20)=>addout_31_31, bb(19)=>
      addout_31_31, bb(18)=>addout_31_31, bb(17)=>addout_31_31, bb(16)=>
      addout_31_31, bb(15)=>addout_31_31, bb(14)=>addout_31_31, bb(13)=>
      addout_31_31, bb(12)=>addout_31_31, bb(11)=>addout_31_31, bb(10)=>
      addout_31_31, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>
      addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_27_31, ff(30)=>addout_27_30, ff(29)=>addout_27_29, ff(28)=>
      addout_27_28, ff(27)=>addout_27_27, ff(26)=>addout_27_26, ff(25)=>
      addout_27_25, ff(24)=>addout_27_24, ff(23)=>addout_27_23, ff(22)=>
      addout_27_22, ff(21)=>addout_27_21, ff(20)=>addout_27_20, ff(19)=>
      addout_27_19, ff(18)=>addout_27_18, ff(17)=>addout_27_17, ff(16)=>
      addout_27_16, ff(15)=>addout_27_15, ff(14)=>addout_27_14, ff(13)=>
      addout_27_13, ff(12)=>addout_27_12, ff(11)=>addout_27_11, ff(10)=>
      addout_27_10, ff(9)=>addout_27_9, ff(8)=>addout_27_8, ff(7)=>
      addout_27_7, ff(6)=>addout_27_6, ff(5)=>addout_27_5, ff(4)=>
      addout_27_4, ff(3)=>addout_27_3, ff(2)=>addout_27_2, ff(1)=>
      addout_27_1, ff(0)=>addout_27_0);
   loop3_28_fx : FC_nadder_32 port map ( aa(31)=>addout_27_31, aa(30)=>
      addout_27_30, aa(29)=>addout_27_29, aa(28)=>addout_27_28, aa(27)=>
      addout_27_27, aa(26)=>addout_27_26, aa(25)=>addout_27_25, aa(24)=>
      addout_27_24, aa(23)=>addout_27_23, aa(22)=>addout_27_22, aa(21)=>
      addout_27_21, aa(20)=>addout_27_20, aa(19)=>addout_27_19, aa(18)=>
      addout_27_18, aa(17)=>addout_27_17, aa(16)=>addout_27_16, aa(15)=>
      addout_27_15, aa(14)=>addout_27_14, aa(13)=>addout_27_13, aa(12)=>
      addout_27_12, aa(11)=>addout_27_11, aa(10)=>addout_27_10, aa(9)=>
      addout_27_9, aa(8)=>addout_27_8, aa(7)=>addout_27_7, aa(6)=>
      addout_27_6, aa(5)=>addout_27_5, aa(4)=>addout_27_4, aa(3)=>
      addout_27_3, aa(2)=>addout_27_2, aa(1)=>addout_27_1, aa(0)=>
      addout_27_0, bb(31)=>nx5984, bb(30)=>nx5996, bb(29)=>nx6010, bb(28)=>
      addout_31_31, bb(27)=>addout_31_31, bb(26)=>addout_31_31, bb(25)=>
      addout_31_31, bb(24)=>addout_31_31, bb(23)=>addout_31_31, bb(22)=>
      addout_31_31, bb(21)=>addout_31_31, bb(20)=>addout_31_31, bb(19)=>
      addout_31_31, bb(18)=>addout_31_31, bb(17)=>addout_31_31, bb(16)=>
      addout_31_31, bb(15)=>addout_31_31, bb(14)=>addout_31_31, bb(13)=>
      addout_31_31, bb(12)=>addout_31_31, bb(11)=>addout_31_31, bb(10)=>
      addout_31_31, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)=>
      addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_28_31, ff(30)=>addout_28_30, ff(29)=>addout_28_29, ff(28)=>
      addout_28_28, ff(27)=>addout_28_27, ff(26)=>addout_28_26, ff(25)=>
      addout_28_25, ff(24)=>addout_28_24, ff(23)=>addout_28_23, ff(22)=>
      addout_28_22, ff(21)=>addout_28_21, ff(20)=>addout_28_20, ff(19)=>
      addout_28_19, ff(18)=>addout_28_18, ff(17)=>addout_28_17, ff(16)=>
      addout_28_16, ff(15)=>addout_28_15, ff(14)=>addout_28_14, ff(13)=>
      addout_28_13, ff(12)=>addout_28_12, ff(11)=>addout_28_11, ff(10)=>
      addout_28_10, ff(9)=>addout_28_9, ff(8)=>addout_28_8, ff(7)=>
      addout_28_7, ff(6)=>addout_28_6, ff(5)=>addout_28_5, ff(4)=>
      addout_28_4, ff(3)=>addout_28_3, ff(2)=>addout_28_2, ff(1)=>
      addout_28_1, ff(0)=>addout_28_0);
   loop3_29_fx : FC_nadder_32 port map ( aa(31)=>addout_28_31, aa(30)=>
      addout_28_30, aa(29)=>addout_28_29, aa(28)=>addout_28_28, aa(27)=>
      addout_28_27, aa(26)=>addout_28_26, aa(25)=>addout_28_25, aa(24)=>
      addout_28_24, aa(23)=>addout_28_23, aa(22)=>addout_28_22, aa(21)=>
      addout_28_21, aa(20)=>addout_28_20, aa(19)=>addout_28_19, aa(18)=>
      addout_28_18, aa(17)=>addout_28_17, aa(16)=>addout_28_16, aa(15)=>
      addout_28_15, aa(14)=>addout_28_14, aa(13)=>addout_28_13, aa(12)=>
      addout_28_12, aa(11)=>addout_28_11, aa(10)=>addout_28_10, aa(9)=>
      addout_28_9, aa(8)=>addout_28_8, aa(7)=>addout_28_7, aa(6)=>
      addout_28_6, aa(5)=>addout_28_5, aa(4)=>addout_28_4, aa(3)=>
      addout_28_3, aa(2)=>addout_28_2, aa(1)=>addout_28_1, aa(0)=>
      addout_28_0, bb(31)=>nx5998, bb(30)=>nx6012, bb(29)=>addout_31_31, 
      bb(28)=>addout_31_31, bb(27)=>addout_31_31, bb(26)=>addout_31_31, 
      bb(25)=>addout_31_31, bb(24)=>addout_31_31, bb(23)=>addout_31_31, 
      bb(22)=>addout_31_31, bb(21)=>addout_31_31, bb(20)=>addout_31_31, 
      bb(19)=>addout_31_31, bb(18)=>addout_31_31, bb(17)=>addout_31_31, 
      bb(16)=>addout_31_31, bb(15)=>addout_31_31, bb(14)=>addout_31_31, 
      bb(13)=>addout_31_31, bb(12)=>addout_31_31, bb(11)=>addout_31_31, 
      bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)=>addout_31_31, bb(7)
      =>addout_31_31, bb(6)=>addout_31_31, bb(5)=>addout_31_31, bb(4)=>
      addout_31_31, bb(3)=>addout_31_31, bb(2)=>addout_31_31, bb(1)=>
      addout_31_31, bb(0)=>addout_31_31, c_cin=>addout_31_31, ff(31)=>
      addout_29_31, ff(30)=>addout_29_30, ff(29)=>addout_29_29, ff(28)=>
      addout_29_28, ff(27)=>addout_29_27, ff(26)=>addout_29_26, ff(25)=>
      addout_29_25, ff(24)=>addout_29_24, ff(23)=>addout_29_23, ff(22)=>
      addout_29_22, ff(21)=>addout_29_21, ff(20)=>addout_29_20, ff(19)=>
      addout_29_19, ff(18)=>addout_29_18, ff(17)=>addout_29_17, ff(16)=>
      addout_29_16, ff(15)=>addout_29_15, ff(14)=>addout_29_14, ff(13)=>
      addout_29_13, ff(12)=>addout_29_12, ff(11)=>addout_29_11, ff(10)=>
      addout_29_10, ff(9)=>addout_29_9, ff(8)=>addout_29_8, ff(7)=>
      addout_29_7, ff(6)=>addout_29_6, ff(5)=>addout_29_5, ff(4)=>
      addout_29_4, ff(3)=>addout_29_3, ff(2)=>addout_29_2, ff(1)=>
      addout_29_1, ff(0)=>addout_29_0);
   loop3_30_fx : FC_nadder_32 port map ( aa(31)=>addout_29_31, aa(30)=>
      addout_29_30, aa(29)=>addout_29_29, aa(28)=>addout_29_28, aa(27)=>
      addout_29_27, aa(26)=>addout_29_26, aa(25)=>addout_29_25, aa(24)=>
      addout_29_24, aa(23)=>addout_29_23, aa(22)=>addout_29_22, aa(21)=>
      addout_29_21, aa(20)=>addout_29_20, aa(19)=>addout_29_19, aa(18)=>
      addout_29_18, aa(17)=>addout_29_17, aa(16)=>addout_29_16, aa(15)=>
      addout_29_15, aa(14)=>addout_29_14, aa(13)=>addout_29_13, aa(12)=>
      addout_29_12, aa(11)=>addout_29_11, aa(10)=>addout_29_10, aa(9)=>
      addout_29_9, aa(8)=>addout_29_8, aa(7)=>addout_29_7, aa(6)=>
      addout_29_6, aa(5)=>addout_29_5, aa(4)=>addout_29_4, aa(3)=>
      addout_29_3, aa(2)=>addout_29_2, aa(1)=>addout_29_1, aa(0)=>
      addout_29_0, bb(31)=>nx6012, bb(30)=>addout_31_31, bb(29)=>
      addout_31_31, bb(28)=>addout_31_31, bb(27)=>addout_31_31, bb(26)=>
      addout_31_31, bb(25)=>addout_31_31, bb(24)=>addout_31_31, bb(23)=>
      addout_31_31, bb(22)=>addout_31_31, bb(21)=>addout_31_31, bb(20)=>
      addout_31_31, bb(19)=>addout_31_31, bb(18)=>addout_31_31, bb(17)=>
      addout_31_31, bb(16)=>addout_31_31, bb(15)=>addout_31_31, bb(14)=>
      addout_31_31, bb(13)=>addout_31_31, bb(12)=>addout_31_31, bb(11)=>
      addout_31_31, bb(10)=>addout_31_31, bb(9)=>addout_31_31, bb(8)=>
      addout_31_31, bb(7)=>addout_31_31, bb(6)=>addout_31_31, bb(5)=>
      addout_31_31, bb(4)=>addout_31_31, bb(3)=>addout_31_31, bb(2)=>
      addout_31_31, bb(1)=>addout_31_31, bb(0)=>addout_31_31, c_cin=>
      addout_31_31, ff(31)=>F(31), ff(30)=>F(30), ff(29)=>F(29), ff(28)=>
      F(28), ff(27)=>F(27), ff(26)=>F(26), ff(25)=>F(25), ff(24)=>F(24), 
      ff(23)=>F(23), ff(22)=>F(22), ff(21)=>F(21), ff(20)=>F(20), ff(19)=>
      F(19), ff(18)=>F(18), ff(17)=>F(17), ff(16)=>F(16), ff(15)=>F(15), 
      ff(14)=>F(14), ff(13)=>F(13), ff(12)=>F(12), ff(11)=>F(11), ff(10)=>
      F(10), ff(9)=>F(9), ff(8)=>F(8), ff(7)=>F(7), ff(6)=>F(6), ff(5)=>F(5), 
      ff(4)=>F(4), ff(3)=>F(3), ff(2)=>F(2), ff(1)=>F(1), ff(0)=>F(0));
   ix5404 : fake_gnd port map ( Y=>addout_31_31);
   ix5769 : inv02 port map ( Y=>nx5770, A=>nx5768);
   ix5771 : inv02 port map ( Y=>nx5772, A=>nx5768);
   ix5773 : inv02 port map ( Y=>nx5774, A=>nx5768);
   ix5775 : inv02 port map ( Y=>nx5776, A=>nx5768);
   ix5777 : inv02 port map ( Y=>nx5778, A=>nx5768);
   ix5779 : inv02 port map ( Y=>nx5780, A=>nx5768);
   ix5783 : inv02 port map ( Y=>nx5784, A=>nx5782);
   ix5785 : inv02 port map ( Y=>nx5786, A=>nx5782);
   ix5787 : inv02 port map ( Y=>nx5788, A=>nx5782);
   ix5789 : inv02 port map ( Y=>nx5790, A=>nx5782);
   ix5791 : inv02 port map ( Y=>nx5792, A=>nx5782);
   ix5795 : inv02 port map ( Y=>nx5796, A=>nx5794);
   ix5797 : inv02 port map ( Y=>nx5798, A=>nx5794);
   ix5799 : inv02 port map ( Y=>nx5800, A=>nx5794);
   ix5801 : inv02 port map ( Y=>nx5802, A=>nx5794);
   ix5803 : inv02 port map ( Y=>nx5804, A=>nx5794);
   ix5807 : inv02 port map ( Y=>nx5808, A=>nx5806);
   ix5809 : inv02 port map ( Y=>nx5810, A=>nx5806);
   ix5811 : inv02 port map ( Y=>nx5812, A=>nx5806);
   ix5813 : inv02 port map ( Y=>nx5814, A=>nx5806);
   ix5815 : inv02 port map ( Y=>nx5816, A=>nx5806);
   ix5819 : inv02 port map ( Y=>nx5820, A=>nx5818);
   ix5821 : inv02 port map ( Y=>nx5822, A=>nx5818);
   ix5823 : inv02 port map ( Y=>nx5824, A=>nx5818);
   ix5825 : inv02 port map ( Y=>nx5826, A=>nx5818);
   ix5829 : inv02 port map ( Y=>nx5830, A=>nx5828);
   ix5831 : inv02 port map ( Y=>nx5832, A=>nx5828);
   ix5833 : inv02 port map ( Y=>nx5834, A=>nx5828);
   ix5835 : inv02 port map ( Y=>nx5836, A=>nx5828);
   ix5839 : inv02 port map ( Y=>nx5840, A=>nx5838);
   ix5841 : inv02 port map ( Y=>nx5842, A=>nx5838);
   ix5843 : inv02 port map ( Y=>nx5844, A=>nx5838);
   ix5845 : inv02 port map ( Y=>nx5846, A=>nx5838);
   ix5849 : inv02 port map ( Y=>nx5850, A=>nx5848);
   ix5851 : inv02 port map ( Y=>nx5852, A=>nx5848);
   ix5853 : inv02 port map ( Y=>nx5854, A=>nx5848);
   ix5857 : inv02 port map ( Y=>nx5858, A=>nx5856);
   ix5859 : inv02 port map ( Y=>nx5860, A=>nx5856);
   ix5861 : inv02 port map ( Y=>nx5862, A=>nx5856);
   ix5865 : inv02 port map ( Y=>nx5866, A=>nx5864);
   ix5867 : inv02 port map ( Y=>nx5868, A=>nx5864);
   ix5869 : inv02 port map ( Y=>nx5870, A=>nx5864);
   ix5871 : buf02 port map ( Y=>nx5872, A=>op2_10_26);
   ix5873 : buf02 port map ( Y=>nx5874, A=>op2_10_26);
   ix5875 : buf02 port map ( Y=>nx5876, A=>op2_11_27);
   ix5877 : buf02 port map ( Y=>nx5878, A=>op2_11_27);
   ix5879 : buf02 port map ( Y=>nx5880, A=>op2_12_28);
   ix5881 : buf02 port map ( Y=>nx5882, A=>op2_12_28);
   ix5883 : buf02 port map ( Y=>nx5884, A=>op2_14_28);
   ix5885 : buf02 port map ( Y=>nx5886, A=>op2_14_28);
   ix5887 : buf02 port map ( Y=>nx5888, A=>op2_14_27);
   ix5889 : buf02 port map ( Y=>nx5890, A=>op2_14_27);
   ix5891 : buf02 port map ( Y=>nx5892, A=>op2_14_26);
   ix5893 : buf02 port map ( Y=>nx5894, A=>op2_14_26);
   ix5897 : inv02 port map ( Y=>nx5898, A=>nx5896);
   ix5899 : inv02 port map ( Y=>nx5900, A=>nx5896);
   ix5901 : inv02 port map ( Y=>nx5902, A=>nx5896);
   ix5905 : inv02 port map ( Y=>nx5906, A=>nx5904);
   ix5907 : inv02 port map ( Y=>nx5908, A=>nx5904);
   ix5909 : inv02 port map ( Y=>nx5910, A=>nx5904);
   ix5913 : inv02 port map ( Y=>nx5914, A=>nx5912);
   ix5915 : inv02 port map ( Y=>nx5916, A=>nx5912);
   ix5917 : inv02 port map ( Y=>nx5918, A=>nx5912);
   ix5921 : inv02 port map ( Y=>nx5922, A=>nx5920);
   ix5923 : inv02 port map ( Y=>nx5924, A=>nx5920);
   ix5925 : inv02 port map ( Y=>nx5926, A=>nx5920);
   ix5927 : inv02 port map ( Y=>nx5928, A=>nx5920);
   ix5931 : inv02 port map ( Y=>nx5932, A=>nx5930);
   ix5933 : inv02 port map ( Y=>nx5934, A=>nx5930);
   ix5935 : inv02 port map ( Y=>nx5936, A=>nx5930);
   ix5937 : inv02 port map ( Y=>nx5938, A=>nx5930);
   ix5941 : inv02 port map ( Y=>nx5942, A=>nx5940);
   ix5943 : inv02 port map ( Y=>nx5944, A=>nx5940);
   ix5945 : inv02 port map ( Y=>nx5946, A=>nx5940);
   ix5947 : inv02 port map ( Y=>nx5948, A=>nx5940);
   ix5951 : inv02 port map ( Y=>nx5952, A=>nx5950);
   ix5953 : inv02 port map ( Y=>nx5954, A=>nx5950);
   ix5955 : inv02 port map ( Y=>nx5956, A=>nx5950);
   ix5957 : inv02 port map ( Y=>nx5958, A=>nx5950);
   ix5959 : inv02 port map ( Y=>nx5960, A=>nx5950);
   ix5963 : inv02 port map ( Y=>nx5964, A=>nx5962);
   ix5965 : inv02 port map ( Y=>nx5966, A=>nx5962);
   ix5967 : inv02 port map ( Y=>nx5968, A=>nx5962);
   ix5969 : inv02 port map ( Y=>nx5970, A=>nx5962);
   ix5971 : inv02 port map ( Y=>nx5972, A=>nx5962);
   ix5975 : inv02 port map ( Y=>nx5976, A=>nx5974);
   ix5977 : inv02 port map ( Y=>nx5978, A=>nx5974);
   ix5979 : inv02 port map ( Y=>nx5980, A=>nx5974);
   ix5981 : inv02 port map ( Y=>nx5982, A=>nx5974);
   ix5983 : inv02 port map ( Y=>nx5984, A=>nx5974);
   ix5987 : inv02 port map ( Y=>nx5988, A=>nx5986);
   ix5989 : inv02 port map ( Y=>nx5990, A=>nx5986);
   ix5991 : inv02 port map ( Y=>nx5992, A=>nx5986);
   ix5993 : inv02 port map ( Y=>nx5994, A=>nx5986);
   ix5995 : inv02 port map ( Y=>nx5996, A=>nx5986);
   ix5997 : inv02 port map ( Y=>nx5998, A=>nx5986);
   ix6001 : inv02 port map ( Y=>nx6002, A=>nx6000);
   ix6003 : inv02 port map ( Y=>nx6004, A=>nx6000);
   ix6005 : inv02 port map ( Y=>nx6006, A=>nx6000);
   ix6007 : inv02 port map ( Y=>nx6008, A=>nx6000);
   ix6009 : inv02 port map ( Y=>nx6010, A=>nx6000);
   ix6011 : inv02 port map ( Y=>nx6012, A=>nx6000);
   ix6015 : inv02 port map ( Y=>nx6016, A=>nx6014);
   ix6017 : inv02 port map ( Y=>nx6018, A=>nx6014);
   ix6019 : inv02 port map ( Y=>nx6020, A=>nx6014);
   ix6021 : inv02 port map ( Y=>nx6022, A=>nx6014);
   ix6023 : inv02 port map ( Y=>nx6024, A=>nx6014);
   ix6025 : inv02 port map ( Y=>nx6026, A=>nx6014);
   ix481 : and02 port map ( Y=>op1_0, A0=>nx6346, A1=>nx6474);
   ix483 : and02 port map ( Y=>op1_1, A0=>nx6338, A1=>nx6474);
   ix485 : and02 port map ( Y=>op1_2, A0=>nx6330, A1=>nx6474);
   ix487 : and02 port map ( Y=>op1_3, A0=>nx6322, A1=>nx6474);
   ix489 : and02 port map ( Y=>op1_4, A0=>nx6314, A1=>nx6474);
   ix491 : and02 port map ( Y=>op1_5, A0=>nx6306, A1=>nx6474);
   ix493 : and02 port map ( Y=>op1_6, A0=>nx6298, A1=>nx6474);
   ix495 : and02 port map ( Y=>op1_7, A0=>nx6290, A1=>nx6476);
   ix497 : and02 port map ( Y=>op1_8, A0=>nx6282, A1=>nx6476);
   ix499 : and02 port map ( Y=>op1_9, A0=>nx6274, A1=>nx6476);
   ix501 : and02 port map ( Y=>op1_10, A0=>nx6266, A1=>nx6476);
   ix503 : and02 port map ( Y=>op1_11, A0=>nx6258, A1=>nx6476);
   ix505 : and02 port map ( Y=>op1_12, A0=>nx6250, A1=>nx6476);
   ix507 : and02 port map ( Y=>op1_13, A0=>nx6242, A1=>nx6476);
   ix509 : and02 port map ( Y=>op1_14, A0=>nx6234, A1=>nx6478);
   ix511 : nand02 port map ( Y=>nx6014, A0=>nx6478, A1=>nx6226);
   ix1 : nand02 port map ( Y=>nx6000, A0=>nx6354, A1=>nx6346);
   ix3 : nand02 port map ( Y=>nx5986, A0=>nx6354, A1=>nx6338);
   ix5 : nand02 port map ( Y=>nx5974, A0=>nx6354, A1=>nx6330);
   ix7 : nand02 port map ( Y=>nx5962, A0=>nx6354, A1=>nx6322);
   ix9 : nand02 port map ( Y=>nx5950, A0=>nx6354, A1=>nx6314);
   ix11 : nand02 port map ( Y=>nx5940, A0=>nx6354, A1=>nx6306);
   ix13 : nand02 port map ( Y=>nx5930, A0=>nx6354, A1=>nx6298);
   ix15 : nand02 port map ( Y=>nx5920, A0=>nx6356, A1=>nx6290);
   ix17 : nand02 port map ( Y=>nx5912, A0=>nx6356, A1=>nx6282);
   ix19 : nand02 port map ( Y=>nx5904, A0=>nx6356, A1=>nx6274);
   ix21 : nand02 port map ( Y=>nx5896, A0=>nx6356, A1=>nx6266);
   ix23 : and02 port map ( Y=>op2_14_26, A0=>nx6356, A1=>nx6258);
   ix25 : and02 port map ( Y=>op2_14_27, A0=>nx6356, A1=>nx6250);
   ix27 : and02 port map ( Y=>op2_14_28, A0=>nx6356, A1=>nx6242);
   ix29 : and02 port map ( Y=>op2_14_29, A0=>nx6358, A1=>nx6234);
   ix31 : and02 port map ( Y=>op2_14_30, A0=>nx6358, A1=>nx6226);
   ix33 : and02 port map ( Y=>op2_13_14, A0=>nx6362, A1=>nx6346);
   ix35 : and02 port map ( Y=>op2_13_15, A0=>nx6362, A1=>nx6338);
   ix37 : and02 port map ( Y=>op2_13_16, A0=>nx6362, A1=>nx6330);
   ix39 : and02 port map ( Y=>op2_13_17, A0=>nx6362, A1=>nx6322);
   ix41 : and02 port map ( Y=>op2_13_18, A0=>nx6362, A1=>nx6314);
   ix43 : and02 port map ( Y=>op2_13_19, A0=>nx6362, A1=>nx6306);
   ix45 : and02 port map ( Y=>op2_13_20, A0=>nx6362, A1=>nx6298);
   ix47 : and02 port map ( Y=>op2_13_21, A0=>nx6364, A1=>nx6290);
   ix49 : and02 port map ( Y=>op2_13_22, A0=>nx6364, A1=>nx6282);
   ix51 : and02 port map ( Y=>op2_13_23, A0=>nx6364, A1=>nx6274);
   ix53 : and02 port map ( Y=>op2_13_24, A0=>nx6364, A1=>nx6266);
   ix55 : and02 port map ( Y=>op2_13_25, A0=>nx6364, A1=>nx6258);
   ix57 : and02 port map ( Y=>op2_13_26, A0=>nx6364, A1=>nx6250);
   ix59 : and02 port map ( Y=>op2_13_27, A0=>nx6364, A1=>nx6242);
   ix61 : and02 port map ( Y=>op2_13_28, A0=>nx6366, A1=>nx6234);
   ix63 : and02 port map ( Y=>op2_13_29, A0=>nx6366, A1=>nx6226);
   ix65 : and02 port map ( Y=>op2_12_13, A0=>nx6370, A1=>nx6346);
   ix67 : and02 port map ( Y=>op2_12_14, A0=>nx6370, A1=>nx6338);
   ix69 : and02 port map ( Y=>op2_12_15, A0=>nx6370, A1=>nx6330);
   ix71 : and02 port map ( Y=>op2_12_16, A0=>nx6370, A1=>nx6322);
   ix73 : and02 port map ( Y=>op2_12_17, A0=>nx6370, A1=>nx6314);
   ix75 : and02 port map ( Y=>op2_12_18, A0=>nx6370, A1=>nx6306);
   ix77 : and02 port map ( Y=>op2_12_19, A0=>nx6370, A1=>nx6298);
   ix79 : and02 port map ( Y=>op2_12_20, A0=>nx6372, A1=>nx6290);
   ix81 : and02 port map ( Y=>op2_12_21, A0=>nx6372, A1=>nx6282);
   ix83 : and02 port map ( Y=>op2_12_22, A0=>nx6372, A1=>nx6274);
   ix85 : and02 port map ( Y=>op2_12_23, A0=>nx6372, A1=>nx6266);
   ix87 : and02 port map ( Y=>op2_12_24, A0=>nx6372, A1=>nx6258);
   ix89 : and02 port map ( Y=>op2_12_25, A0=>nx6372, A1=>nx6250);
   ix91 : and02 port map ( Y=>op2_12_26, A0=>nx6372, A1=>nx6242);
   ix93 : and02 port map ( Y=>op2_12_27, A0=>nx6374, A1=>nx6234);
   ix95 : and02 port map ( Y=>op2_12_28, A0=>nx6374, A1=>nx6226);
   ix97 : and02 port map ( Y=>op2_11_12, A0=>nx6378, A1=>nx6346);
   ix99 : and02 port map ( Y=>op2_11_13, A0=>nx6378, A1=>nx6338);
   ix101 : and02 port map ( Y=>op2_11_14, A0=>nx6378, A1=>nx6330);
   ix103 : and02 port map ( Y=>op2_11_15, A0=>nx6378, A1=>nx6322);
   ix105 : and02 port map ( Y=>op2_11_16, A0=>nx6378, A1=>nx6314);
   ix107 : and02 port map ( Y=>op2_11_17, A0=>nx6378, A1=>nx6306);
   ix109 : and02 port map ( Y=>op2_11_18, A0=>nx6378, A1=>nx6298);
   ix111 : and02 port map ( Y=>op2_11_19, A0=>nx6380, A1=>nx6290);
   ix113 : and02 port map ( Y=>op2_11_20, A0=>nx6380, A1=>nx6282);
   ix115 : and02 port map ( Y=>op2_11_21, A0=>nx6380, A1=>nx6274);
   ix117 : and02 port map ( Y=>op2_11_22, A0=>nx6380, A1=>nx6266);
   ix119 : and02 port map ( Y=>op2_11_23, A0=>nx6380, A1=>nx6258);
   ix121 : and02 port map ( Y=>op2_11_24, A0=>nx6380, A1=>nx6250);
   ix123 : and02 port map ( Y=>op2_11_25, A0=>nx6380, A1=>nx6242);
   ix125 : and02 port map ( Y=>op2_11_26, A0=>nx6382, A1=>nx6234);
   ix127 : and02 port map ( Y=>op2_11_27, A0=>nx6382, A1=>nx6226);
   ix129 : and02 port map ( Y=>op2_10_11, A0=>nx6386, A1=>nx6346);
   ix131 : and02 port map ( Y=>op2_10_12, A0=>nx6386, A1=>nx6338);
   ix133 : and02 port map ( Y=>op2_10_13, A0=>nx6386, A1=>nx6330);
   ix135 : and02 port map ( Y=>op2_10_14, A0=>nx6386, A1=>nx6322);
   ix137 : and02 port map ( Y=>op2_10_15, A0=>nx6386, A1=>nx6314);
   ix139 : and02 port map ( Y=>op2_10_16, A0=>nx6386, A1=>nx6306);
   ix141 : and02 port map ( Y=>op2_10_17, A0=>nx6386, A1=>nx6298);
   ix143 : and02 port map ( Y=>op2_10_18, A0=>nx6388, A1=>nx6290);
   ix145 : and02 port map ( Y=>op2_10_19, A0=>nx6388, A1=>nx6282);
   ix147 : and02 port map ( Y=>op2_10_20, A0=>nx6388, A1=>nx6274);
   ix149 : and02 port map ( Y=>op2_10_21, A0=>nx6388, A1=>nx6266);
   ix151 : and02 port map ( Y=>op2_10_22, A0=>nx6388, A1=>nx6258);
   ix153 : and02 port map ( Y=>op2_10_23, A0=>nx6388, A1=>nx6250);
   ix155 : and02 port map ( Y=>op2_10_24, A0=>nx6388, A1=>nx6242);
   ix157 : and02 port map ( Y=>op2_10_25, A0=>nx6390, A1=>nx6234);
   ix159 : and02 port map ( Y=>op2_10_26, A0=>nx6390, A1=>nx6226);
   ix161 : and02 port map ( Y=>op2_9_10, A0=>nx6394, A1=>nx6346);
   ix163 : and02 port map ( Y=>op2_9_11, A0=>nx6394, A1=>nx6338);
   ix165 : and02 port map ( Y=>op2_9_12, A0=>nx6394, A1=>nx6330);
   ix167 : and02 port map ( Y=>op2_9_13, A0=>nx6394, A1=>nx6322);
   ix169 : and02 port map ( Y=>op2_9_14, A0=>nx6394, A1=>nx6314);
   ix171 : and02 port map ( Y=>op2_9_15, A0=>nx6394, A1=>nx6306);
   ix173 : and02 port map ( Y=>op2_9_16, A0=>nx6394, A1=>nx6298);
   ix175 : and02 port map ( Y=>op2_9_17, A0=>nx6396, A1=>nx6290);
   ix177 : and02 port map ( Y=>op2_9_18, A0=>nx6396, A1=>nx6282);
   ix179 : and02 port map ( Y=>op2_9_19, A0=>nx6396, A1=>nx6274);
   ix181 : and02 port map ( Y=>op2_9_20, A0=>nx6396, A1=>nx6266);
   ix183 : and02 port map ( Y=>op2_9_21, A0=>nx6396, A1=>nx6258);
   ix185 : and02 port map ( Y=>op2_9_22, A0=>nx6396, A1=>nx6250);
   ix187 : and02 port map ( Y=>op2_9_23, A0=>nx6396, A1=>nx6242);
   ix189 : and02 port map ( Y=>op2_9_24, A0=>nx6398, A1=>nx6234);
   ix191 : nand02 port map ( Y=>nx5864, A0=>nx6398, A1=>nx6226);
   ix193 : and02 port map ( Y=>op2_8_9, A0=>nx6402, A1=>nx6348);
   ix195 : and02 port map ( Y=>op2_8_10, A0=>nx6402, A1=>nx6340);
   ix197 : and02 port map ( Y=>op2_8_11, A0=>nx6402, A1=>nx6332);
   ix199 : and02 port map ( Y=>op2_8_12, A0=>nx6402, A1=>nx6324);
   ix201 : and02 port map ( Y=>op2_8_13, A0=>nx6402, A1=>nx6316);
   ix203 : and02 port map ( Y=>op2_8_14, A0=>nx6402, A1=>nx6308);
   ix205 : and02 port map ( Y=>op2_8_15, A0=>nx6402, A1=>nx6300);
   ix207 : and02 port map ( Y=>op2_8_16, A0=>nx6404, A1=>nx6292);
   ix209 : and02 port map ( Y=>op2_8_17, A0=>nx6404, A1=>nx6284);
   ix211 : and02 port map ( Y=>op2_8_18, A0=>nx6404, A1=>nx6276);
   ix213 : and02 port map ( Y=>op2_8_19, A0=>nx6404, A1=>nx6268);
   ix215 : and02 port map ( Y=>op2_8_20, A0=>nx6404, A1=>nx6260);
   ix217 : and02 port map ( Y=>op2_8_21, A0=>nx6404, A1=>nx6252);
   ix219 : and02 port map ( Y=>op2_8_22, A0=>nx6404, A1=>nx6244);
   ix221 : and02 port map ( Y=>op2_8_23, A0=>nx6406, A1=>nx6236);
   ix223 : nand02 port map ( Y=>nx5856, A0=>nx6406, A1=>nx6228);
   ix225 : and02 port map ( Y=>op2_7_8, A0=>nx6410, A1=>nx6348);
   ix227 : and02 port map ( Y=>op2_7_9, A0=>nx6410, A1=>nx6340);
   ix229 : and02 port map ( Y=>op2_7_10, A0=>nx6410, A1=>nx6332);
   ix231 : and02 port map ( Y=>op2_7_11, A0=>nx6410, A1=>nx6324);
   ix233 : and02 port map ( Y=>op2_7_12, A0=>nx6410, A1=>nx6316);
   ix235 : and02 port map ( Y=>op2_7_13, A0=>nx6410, A1=>nx6308);
   ix237 : and02 port map ( Y=>op2_7_14, A0=>nx6410, A1=>nx6300);
   ix239 : and02 port map ( Y=>op2_7_15, A0=>nx6412, A1=>nx6292);
   ix241 : and02 port map ( Y=>op2_7_16, A0=>nx6412, A1=>nx6284);
   ix243 : and02 port map ( Y=>op2_7_17, A0=>nx6412, A1=>nx6276);
   ix245 : and02 port map ( Y=>op2_7_18, A0=>nx6412, A1=>nx6268);
   ix247 : and02 port map ( Y=>op2_7_19, A0=>nx6412, A1=>nx6260);
   ix249 : and02 port map ( Y=>op2_7_20, A0=>nx6412, A1=>nx6252);
   ix251 : and02 port map ( Y=>op2_7_21, A0=>nx6412, A1=>nx6244);
   ix253 : and02 port map ( Y=>op2_7_22, A0=>nx6414, A1=>nx6236);
   ix255 : nand02 port map ( Y=>nx5848, A0=>nx6414, A1=>nx6228);
   ix257 : and02 port map ( Y=>op2_6_7, A0=>nx6418, A1=>nx6348);
   ix259 : and02 port map ( Y=>op2_6_8, A0=>nx6418, A1=>nx6340);
   ix261 : and02 port map ( Y=>op2_6_9, A0=>nx6418, A1=>nx6332);
   ix263 : and02 port map ( Y=>op2_6_10, A0=>nx6418, A1=>nx6324);
   ix265 : and02 port map ( Y=>op2_6_11, A0=>nx6418, A1=>nx6316);
   ix267 : and02 port map ( Y=>op2_6_12, A0=>nx6418, A1=>nx6308);
   ix269 : and02 port map ( Y=>op2_6_13, A0=>nx6418, A1=>nx6300);
   ix271 : and02 port map ( Y=>op2_6_14, A0=>nx6420, A1=>nx6292);
   ix273 : and02 port map ( Y=>op2_6_15, A0=>nx6420, A1=>nx6284);
   ix275 : and02 port map ( Y=>op2_6_16, A0=>nx6420, A1=>nx6276);
   ix277 : and02 port map ( Y=>op2_6_17, A0=>nx6420, A1=>nx6268);
   ix279 : and02 port map ( Y=>op2_6_18, A0=>nx6420, A1=>nx6260);
   ix281 : and02 port map ( Y=>op2_6_19, A0=>nx6420, A1=>nx6252);
   ix283 : and02 port map ( Y=>op2_6_20, A0=>nx6420, A1=>nx6244);
   ix285 : and02 port map ( Y=>op2_6_21, A0=>nx6422, A1=>nx6236);
   ix287 : nand02 port map ( Y=>nx5838, A0=>nx6422, A1=>nx6228);
   ix289 : and02 port map ( Y=>op2_5_6, A0=>nx6426, A1=>nx6348);
   ix291 : and02 port map ( Y=>op2_5_7, A0=>nx6426, A1=>nx6340);
   ix293 : and02 port map ( Y=>op2_5_8, A0=>nx6426, A1=>nx6332);
   ix295 : and02 port map ( Y=>op2_5_9, A0=>nx6426, A1=>nx6324);
   ix297 : and02 port map ( Y=>op2_5_10, A0=>nx6426, A1=>nx6316);
   ix299 : and02 port map ( Y=>op2_5_11, A0=>nx6426, A1=>nx6308);
   ix301 : and02 port map ( Y=>op2_5_12, A0=>nx6426, A1=>nx6300);
   ix303 : and02 port map ( Y=>op2_5_13, A0=>nx6428, A1=>nx6292);
   ix305 : and02 port map ( Y=>op2_5_14, A0=>nx6428, A1=>nx6284);
   ix307 : and02 port map ( Y=>op2_5_15, A0=>nx6428, A1=>nx6276);
   ix309 : and02 port map ( Y=>op2_5_16, A0=>nx6428, A1=>nx6268);
   ix311 : and02 port map ( Y=>op2_5_17, A0=>nx6428, A1=>nx6260);
   ix313 : and02 port map ( Y=>op2_5_18, A0=>nx6428, A1=>nx6252);
   ix315 : and02 port map ( Y=>op2_5_19, A0=>nx6428, A1=>nx6244);
   ix317 : and02 port map ( Y=>op2_5_20, A0=>nx6430, A1=>nx6236);
   ix319 : nand02 port map ( Y=>nx5828, A0=>nx6430, A1=>nx6228);
   ix321 : and02 port map ( Y=>op2_4_5, A0=>nx6434, A1=>nx6348);
   ix323 : and02 port map ( Y=>op2_4_6, A0=>nx6434, A1=>nx6340);
   ix325 : and02 port map ( Y=>op2_4_7, A0=>nx6434, A1=>nx6332);
   ix327 : and02 port map ( Y=>op2_4_8, A0=>nx6434, A1=>nx6324);
   ix329 : and02 port map ( Y=>op2_4_9, A0=>nx6434, A1=>nx6316);
   ix331 : and02 port map ( Y=>op2_4_10, A0=>nx6434, A1=>nx6308);
   ix333 : and02 port map ( Y=>op2_4_11, A0=>nx6434, A1=>nx6300);
   ix335 : and02 port map ( Y=>op2_4_12, A0=>nx6436, A1=>nx6292);
   ix337 : and02 port map ( Y=>op2_4_13, A0=>nx6436, A1=>nx6284);
   ix339 : and02 port map ( Y=>op2_4_14, A0=>nx6436, A1=>nx6276);
   ix341 : and02 port map ( Y=>op2_4_15, A0=>nx6436, A1=>nx6268);
   ix343 : and02 port map ( Y=>op2_4_16, A0=>nx6436, A1=>nx6260);
   ix345 : and02 port map ( Y=>op2_4_17, A0=>nx6436, A1=>nx6252);
   ix347 : and02 port map ( Y=>op2_4_18, A0=>nx6436, A1=>nx6244);
   ix349 : and02 port map ( Y=>op2_4_19, A0=>nx6438, A1=>nx6236);
   ix351 : nand02 port map ( Y=>nx5818, A0=>nx6438, A1=>nx6228);
   ix353 : and02 port map ( Y=>op2_3_4, A0=>nx6442, A1=>nx6348);
   ix355 : and02 port map ( Y=>op2_3_5, A0=>nx6442, A1=>nx6340);
   ix357 : and02 port map ( Y=>op2_3_6, A0=>nx6442, A1=>nx6332);
   ix359 : and02 port map ( Y=>op2_3_7, A0=>nx6442, A1=>nx6324);
   ix361 : and02 port map ( Y=>op2_3_8, A0=>nx6442, A1=>nx6316);
   ix363 : and02 port map ( Y=>op2_3_9, A0=>nx6442, A1=>nx6308);
   ix365 : and02 port map ( Y=>op2_3_10, A0=>nx6442, A1=>nx6300);
   ix367 : and02 port map ( Y=>op2_3_11, A0=>nx6444, A1=>nx6292);
   ix369 : and02 port map ( Y=>op2_3_12, A0=>nx6444, A1=>nx6284);
   ix371 : and02 port map ( Y=>op2_3_13, A0=>nx6444, A1=>nx6276);
   ix373 : and02 port map ( Y=>op2_3_14, A0=>nx6444, A1=>nx6268);
   ix375 : and02 port map ( Y=>op2_3_15, A0=>nx6444, A1=>nx6260);
   ix377 : and02 port map ( Y=>op2_3_16, A0=>nx6444, A1=>nx6252);
   ix379 : and02 port map ( Y=>op2_3_17, A0=>nx6444, A1=>nx6244);
   ix381 : and02 port map ( Y=>op2_3_18, A0=>nx6446, A1=>nx6236);
   ix383 : nand02 port map ( Y=>nx5806, A0=>nx6446, A1=>nx6228);
   ix385 : and02 port map ( Y=>op2_2_3, A0=>nx6450, A1=>nx6348);
   ix387 : and02 port map ( Y=>op2_2_4, A0=>nx6450, A1=>nx6340);
   ix389 : and02 port map ( Y=>op2_2_5, A0=>nx6450, A1=>nx6332);
   ix391 : and02 port map ( Y=>op2_2_6, A0=>nx6450, A1=>nx6324);
   ix393 : and02 port map ( Y=>op2_2_7, A0=>nx6450, A1=>nx6316);
   ix395 : and02 port map ( Y=>op2_2_8, A0=>nx6450, A1=>nx6308);
   ix397 : and02 port map ( Y=>op2_2_9, A0=>nx6450, A1=>nx6300);
   ix399 : and02 port map ( Y=>op2_2_10, A0=>nx6452, A1=>nx6292);
   ix401 : and02 port map ( Y=>op2_2_11, A0=>nx6452, A1=>nx6284);
   ix403 : and02 port map ( Y=>op2_2_12, A0=>nx6452, A1=>nx6276);
   ix405 : and02 port map ( Y=>op2_2_13, A0=>nx6452, A1=>nx6268);
   ix407 : and02 port map ( Y=>op2_2_14, A0=>nx6452, A1=>nx6260);
   ix409 : and02 port map ( Y=>op2_2_15, A0=>nx6452, A1=>nx6252);
   ix411 : and02 port map ( Y=>op2_2_16, A0=>nx6452, A1=>nx6244);
   ix413 : and02 port map ( Y=>op2_2_17, A0=>nx6454, A1=>nx6236);
   ix415 : nand02 port map ( Y=>nx5794, A0=>nx6454, A1=>nx6228);
   ix417 : and02 port map ( Y=>op2_1_2, A0=>nx6458, A1=>nx6350);
   ix419 : and02 port map ( Y=>op2_1_3, A0=>nx6458, A1=>nx6342);
   ix421 : and02 port map ( Y=>op2_1_4, A0=>nx6458, A1=>nx6334);
   ix423 : and02 port map ( Y=>op2_1_5, A0=>nx6458, A1=>nx6326);
   ix425 : and02 port map ( Y=>op2_1_6, A0=>nx6458, A1=>nx6318);
   ix427 : and02 port map ( Y=>op2_1_7, A0=>nx6458, A1=>nx6310);
   ix429 : and02 port map ( Y=>op2_1_8, A0=>nx6458, A1=>nx6302);
   ix431 : and02 port map ( Y=>op2_1_9, A0=>nx6460, A1=>nx6294);
   ix433 : and02 port map ( Y=>op2_1_10, A0=>nx6460, A1=>nx6286);
   ix435 : and02 port map ( Y=>op2_1_11, A0=>nx6460, A1=>nx6278);
   ix437 : and02 port map ( Y=>op2_1_12, A0=>nx6460, A1=>nx6270);
   ix439 : and02 port map ( Y=>op2_1_13, A0=>nx6460, A1=>nx6262);
   ix441 : and02 port map ( Y=>op2_1_14, A0=>nx6460, A1=>nx6254);
   ix443 : and02 port map ( Y=>op2_1_15, A0=>nx6460, A1=>nx6246);
   ix445 : and02 port map ( Y=>op2_1_16, A0=>nx6462, A1=>nx6238);
   ix447 : nand02 port map ( Y=>nx5782, A0=>nx6462, A1=>nx6230);
   ix449 : and02 port map ( Y=>op2_0_1, A0=>nx6466, A1=>nx6350);
   ix451 : and02 port map ( Y=>op2_0_2, A0=>nx6466, A1=>nx6342);
   ix453 : and02 port map ( Y=>op2_0_3, A0=>nx6466, A1=>nx6334);
   ix455 : and02 port map ( Y=>op2_0_4, A0=>nx6466, A1=>nx6326);
   ix457 : and02 port map ( Y=>op2_0_5, A0=>nx6466, A1=>nx6318);
   ix459 : and02 port map ( Y=>op2_0_6, A0=>nx6466, A1=>nx6310);
   ix461 : and02 port map ( Y=>op2_0_7, A0=>nx6466, A1=>nx6302);
   ix463 : and02 port map ( Y=>op2_0_8, A0=>nx6468, A1=>nx6294);
   ix465 : and02 port map ( Y=>op2_0_9, A0=>nx6468, A1=>nx6286);
   ix467 : and02 port map ( Y=>op2_0_10, A0=>nx6468, A1=>nx6278);
   ix469 : and02 port map ( Y=>op2_0_11, A0=>nx6468, A1=>nx6270);
   ix471 : and02 port map ( Y=>op2_0_12, A0=>nx6468, A1=>nx6262);
   ix473 : and02 port map ( Y=>op2_0_13, A0=>nx6468, A1=>nx6254);
   ix475 : and02 port map ( Y=>op2_0_14, A0=>nx6468, A1=>nx6246);
   ix477 : and02 port map ( Y=>op2_0_15, A0=>nx6470, A1=>nx6238);
   ix479 : nand02 port map ( Y=>nx5768, A0=>nx6470, A1=>nx6230);
   ix6223 : inv01 port map ( Y=>nx6224, A=>A(15));
   ix6225 : inv02 port map ( Y=>nx6226, A=>nx6224);
   ix6227 : inv02 port map ( Y=>nx6228, A=>nx6224);
   ix6229 : inv02 port map ( Y=>nx6230, A=>nx6224);
   ix6231 : inv01 port map ( Y=>nx6232, A=>A(14));
   ix6233 : inv02 port map ( Y=>nx6234, A=>nx6232);
   ix6235 : inv02 port map ( Y=>nx6236, A=>nx6232);
   ix6237 : inv02 port map ( Y=>nx6238, A=>nx6232);
   ix6239 : inv01 port map ( Y=>nx6240, A=>A(13));
   ix6241 : inv02 port map ( Y=>nx6242, A=>nx6240);
   ix6243 : inv02 port map ( Y=>nx6244, A=>nx6240);
   ix6245 : inv02 port map ( Y=>nx6246, A=>nx6240);
   ix6247 : inv01 port map ( Y=>nx6248, A=>A(12));
   ix6249 : inv02 port map ( Y=>nx6250, A=>nx6248);
   ix6251 : inv02 port map ( Y=>nx6252, A=>nx6248);
   ix6253 : inv02 port map ( Y=>nx6254, A=>nx6248);
   ix6255 : inv01 port map ( Y=>nx6256, A=>A(11));
   ix6257 : inv02 port map ( Y=>nx6258, A=>nx6256);
   ix6259 : inv02 port map ( Y=>nx6260, A=>nx6256);
   ix6261 : inv02 port map ( Y=>nx6262, A=>nx6256);
   ix6263 : inv01 port map ( Y=>nx6264, A=>A(10));
   ix6265 : inv02 port map ( Y=>nx6266, A=>nx6264);
   ix6267 : inv02 port map ( Y=>nx6268, A=>nx6264);
   ix6269 : inv02 port map ( Y=>nx6270, A=>nx6264);
   ix6271 : inv01 port map ( Y=>nx6272, A=>A(9));
   ix6273 : inv02 port map ( Y=>nx6274, A=>nx6272);
   ix6275 : inv02 port map ( Y=>nx6276, A=>nx6272);
   ix6277 : inv02 port map ( Y=>nx6278, A=>nx6272);
   ix6279 : inv01 port map ( Y=>nx6280, A=>A(8));
   ix6281 : inv02 port map ( Y=>nx6282, A=>nx6280);
   ix6283 : inv02 port map ( Y=>nx6284, A=>nx6280);
   ix6285 : inv02 port map ( Y=>nx6286, A=>nx6280);
   ix6287 : inv01 port map ( Y=>nx6288, A=>A(7));
   ix6289 : inv02 port map ( Y=>nx6290, A=>nx6288);
   ix6291 : inv02 port map ( Y=>nx6292, A=>nx6288);
   ix6293 : inv02 port map ( Y=>nx6294, A=>nx6288);
   ix6295 : inv01 port map ( Y=>nx6296, A=>A(6));
   ix6297 : inv02 port map ( Y=>nx6298, A=>nx6296);
   ix6299 : inv02 port map ( Y=>nx6300, A=>nx6296);
   ix6301 : inv02 port map ( Y=>nx6302, A=>nx6296);
   ix6303 : inv01 port map ( Y=>nx6304, A=>A(5));
   ix6305 : inv02 port map ( Y=>nx6306, A=>nx6304);
   ix6307 : inv02 port map ( Y=>nx6308, A=>nx6304);
   ix6309 : inv02 port map ( Y=>nx6310, A=>nx6304);
   ix6311 : inv01 port map ( Y=>nx6312, A=>A(4));
   ix6313 : inv02 port map ( Y=>nx6314, A=>nx6312);
   ix6315 : inv02 port map ( Y=>nx6316, A=>nx6312);
   ix6317 : inv02 port map ( Y=>nx6318, A=>nx6312);
   ix6319 : inv01 port map ( Y=>nx6320, A=>A(3));
   ix6321 : inv02 port map ( Y=>nx6322, A=>nx6320);
   ix6323 : inv02 port map ( Y=>nx6324, A=>nx6320);
   ix6325 : inv02 port map ( Y=>nx6326, A=>nx6320);
   ix6327 : inv01 port map ( Y=>nx6328, A=>A(2));
   ix6329 : inv02 port map ( Y=>nx6330, A=>nx6328);
   ix6331 : inv02 port map ( Y=>nx6332, A=>nx6328);
   ix6333 : inv02 port map ( Y=>nx6334, A=>nx6328);
   ix6335 : inv01 port map ( Y=>nx6336, A=>A(1));
   ix6337 : inv02 port map ( Y=>nx6338, A=>nx6336);
   ix6339 : inv02 port map ( Y=>nx6340, A=>nx6336);
   ix6341 : inv02 port map ( Y=>nx6342, A=>nx6336);
   ix6343 : inv01 port map ( Y=>nx6344, A=>A(0));
   ix6345 : inv02 port map ( Y=>nx6346, A=>nx6344);
   ix6347 : inv02 port map ( Y=>nx6348, A=>nx6344);
   ix6349 : inv02 port map ( Y=>nx6350, A=>nx6344);
   ix6351 : inv01 port map ( Y=>nx6352, A=>B(15));
   ix6353 : inv01 port map ( Y=>nx6354, A=>nx6352);
   ix6355 : inv01 port map ( Y=>nx6356, A=>nx6352);
   ix6357 : inv01 port map ( Y=>nx6358, A=>nx6352);
   ix6359 : inv01 port map ( Y=>nx6360, A=>B(14));
   ix6361 : inv01 port map ( Y=>nx6362, A=>nx6360);
   ix6363 : inv01 port map ( Y=>nx6364, A=>nx6360);
   ix6365 : inv01 port map ( Y=>nx6366, A=>nx6360);
   ix6367 : inv01 port map ( Y=>nx6368, A=>B(13));
   ix6369 : inv01 port map ( Y=>nx6370, A=>nx6368);
   ix6371 : inv01 port map ( Y=>nx6372, A=>nx6368);
   ix6373 : inv01 port map ( Y=>nx6374, A=>nx6368);
   ix6375 : inv01 port map ( Y=>nx6376, A=>B(12));
   ix6377 : inv01 port map ( Y=>nx6378, A=>nx6376);
   ix6379 : inv01 port map ( Y=>nx6380, A=>nx6376);
   ix6381 : inv01 port map ( Y=>nx6382, A=>nx6376);
   ix6383 : inv01 port map ( Y=>nx6384, A=>B(11));
   ix6385 : inv01 port map ( Y=>nx6386, A=>nx6384);
   ix6387 : inv01 port map ( Y=>nx6388, A=>nx6384);
   ix6389 : inv01 port map ( Y=>nx6390, A=>nx6384);
   ix6391 : inv01 port map ( Y=>nx6392, A=>B(10));
   ix6393 : inv01 port map ( Y=>nx6394, A=>nx6392);
   ix6395 : inv01 port map ( Y=>nx6396, A=>nx6392);
   ix6397 : inv01 port map ( Y=>nx6398, A=>nx6392);
   ix6399 : inv01 port map ( Y=>nx6400, A=>B(9));
   ix6401 : inv01 port map ( Y=>nx6402, A=>nx6400);
   ix6403 : inv01 port map ( Y=>nx6404, A=>nx6400);
   ix6405 : inv01 port map ( Y=>nx6406, A=>nx6400);
   ix6407 : inv01 port map ( Y=>nx6408, A=>B(8));
   ix6409 : inv01 port map ( Y=>nx6410, A=>nx6408);
   ix6411 : inv01 port map ( Y=>nx6412, A=>nx6408);
   ix6413 : inv01 port map ( Y=>nx6414, A=>nx6408);
   ix6415 : inv01 port map ( Y=>nx6416, A=>B(7));
   ix6417 : inv01 port map ( Y=>nx6418, A=>nx6416);
   ix6419 : inv01 port map ( Y=>nx6420, A=>nx6416);
   ix6421 : inv01 port map ( Y=>nx6422, A=>nx6416);
   ix6423 : inv01 port map ( Y=>nx6424, A=>B(6));
   ix6425 : inv01 port map ( Y=>nx6426, A=>nx6424);
   ix6427 : inv01 port map ( Y=>nx6428, A=>nx6424);
   ix6429 : inv01 port map ( Y=>nx6430, A=>nx6424);
   ix6431 : inv01 port map ( Y=>nx6432, A=>B(5));
   ix6433 : inv01 port map ( Y=>nx6434, A=>nx6432);
   ix6435 : inv01 port map ( Y=>nx6436, A=>nx6432);
   ix6437 : inv01 port map ( Y=>nx6438, A=>nx6432);
   ix6439 : inv01 port map ( Y=>nx6440, A=>B(4));
   ix6441 : inv01 port map ( Y=>nx6442, A=>nx6440);
   ix6443 : inv01 port map ( Y=>nx6444, A=>nx6440);
   ix6445 : inv01 port map ( Y=>nx6446, A=>nx6440);
   ix6447 : inv01 port map ( Y=>nx6448, A=>B(3));
   ix6449 : inv01 port map ( Y=>nx6450, A=>nx6448);
   ix6451 : inv01 port map ( Y=>nx6452, A=>nx6448);
   ix6453 : inv01 port map ( Y=>nx6454, A=>nx6448);
   ix6455 : inv01 port map ( Y=>nx6456, A=>B(2));
   ix6457 : inv01 port map ( Y=>nx6458, A=>nx6456);
   ix6459 : inv01 port map ( Y=>nx6460, A=>nx6456);
   ix6461 : inv01 port map ( Y=>nx6462, A=>nx6456);
   ix6463 : inv01 port map ( Y=>nx6464, A=>B(1));
   ix6465 : inv01 port map ( Y=>nx6466, A=>nx6464);
   ix6467 : inv01 port map ( Y=>nx6468, A=>nx6464);
   ix6469 : inv01 port map ( Y=>nx6470, A=>nx6464);
   ix6471 : inv01 port map ( Y=>nx6472, A=>B(0));
   ix6473 : inv02 port map ( Y=>nx6474, A=>nx6472);
   ix6475 : inv02 port map ( Y=>nx6476, A=>nx6472);
   ix6477 : inv02 port map ( Y=>nx6478, A=>nx6472);
   ix6479 : buf02 port map ( Y=>nx6480, A=>op2_13_29);
   ix6481 : buf02 port map ( Y=>nx6482, A=>op2_14_30);
   ix6483 : buf02 port map ( Y=>nx6484, A=>op2_14_29);
end Flow ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Convolution is
   port (
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      QImgStat : IN std_logic ;
      ACK : OUT std_logic ;
      LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
      ImgAddress : IN std_logic_vector (12 DOWNTO 0) ;
      OutputImg0 : IN std_logic_vector (79 DOWNTO 0) ;
      OutputImg1 : IN std_logic_vector (79 DOWNTO 0) ;
      OutputImg2 : IN std_logic_vector (79 DOWNTO 0) ;
      OutputImg3 : IN std_logic_vector (79 DOWNTO 0) ;
      OutputImg4 : IN std_logic_vector (79 DOWNTO 0) ;
      outFilter0 : IN std_logic_vector (399 DOWNTO 0) ;
      outFilter1 : IN std_logic_vector (399 DOWNTO 0) ;
      ConvOuput : OUT std_logic_vector (15 DOWNTO 0)) ;
end Convolution ;

architecture ConvArch of Convolution is
   component Multiplier_16
      port (
         A : IN std_logic_vector (15 DOWNTO 0) ;
         B : IN std_logic_vector (15 DOWNTO 0) ;
         F : OUT std_logic_vector (31 DOWNTO 0)) ;
   end component ;
   component my_nadder_16
      port (
         a : IN std_logic_vector (15 DOWNTO 0) ;
         b : IN std_logic_vector (15 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (15 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component Counter_3
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (2 DOWNTO 0) ;
         input : IN std_logic_vector (2 DOWNTO 0)) ;
   end component ;
   signal ACK_EXMPLR, ConvOuput_15_EXMPLR, FilterToAlu_399, FilterToAlu_398, 
      FilterToAlu_397, FilterToAlu_396, FilterToAlu_395, FilterToAlu_394, 
      FilterToAlu_393, FilterToAlu_392, FilterToAlu_391, FilterToAlu_390, 
      FilterToAlu_389, FilterToAlu_388, FilterToAlu_387, FilterToAlu_386, 
      FilterToAlu_385, FilterToAlu_384, FilterToAlu_383, FilterToAlu_382, 
      FilterToAlu_381, FilterToAlu_380, FilterToAlu_379, FilterToAlu_378, 
      FilterToAlu_377, FilterToAlu_376, FilterToAlu_375, FilterToAlu_374, 
      FilterToAlu_373, FilterToAlu_372, FilterToAlu_371, FilterToAlu_370, 
      FilterToAlu_369, FilterToAlu_368, FilterToAlu_367, FilterToAlu_366, 
      FilterToAlu_365, FilterToAlu_364, FilterToAlu_363, FilterToAlu_362, 
      FilterToAlu_361, FilterToAlu_360, FilterToAlu_359, FilterToAlu_358, 
      FilterToAlu_357, FilterToAlu_356, FilterToAlu_355, FilterToAlu_354, 
      FilterToAlu_353, FilterToAlu_352, FilterToAlu_351, FilterToAlu_350, 
      FilterToAlu_349, FilterToAlu_348, FilterToAlu_347, FilterToAlu_346, 
      FilterToAlu_345, FilterToAlu_344, FilterToAlu_343, FilterToAlu_342, 
      FilterToAlu_341, FilterToAlu_340, FilterToAlu_339, FilterToAlu_338, 
      FilterToAlu_337, FilterToAlu_336, FilterToAlu_335, FilterToAlu_334, 
      FilterToAlu_333, FilterToAlu_332, FilterToAlu_331, FilterToAlu_330, 
      FilterToAlu_329, FilterToAlu_328, FilterToAlu_327, FilterToAlu_326, 
      FilterToAlu_325, FilterToAlu_324, FilterToAlu_323, FilterToAlu_322, 
      FilterToAlu_321, FilterToAlu_320, FilterToAlu_319, FilterToAlu_318, 
      FilterToAlu_317, FilterToAlu_316, FilterToAlu_315, FilterToAlu_314, 
      FilterToAlu_313, FilterToAlu_312, FilterToAlu_311, FilterToAlu_310, 
      FilterToAlu_309, FilterToAlu_308, FilterToAlu_307, FilterToAlu_306, 
      FilterToAlu_305, FilterToAlu_304, FilterToAlu_303, FilterToAlu_302, 
      FilterToAlu_301, FilterToAlu_300, FilterToAlu_299, FilterToAlu_298, 
      FilterToAlu_297, FilterToAlu_296, FilterToAlu_295, FilterToAlu_294, 
      FilterToAlu_293, FilterToAlu_292, FilterToAlu_291, FilterToAlu_290, 
      FilterToAlu_289, FilterToAlu_288, FilterToAlu_287, FilterToAlu_286, 
      FilterToAlu_285, FilterToAlu_284, FilterToAlu_283, FilterToAlu_282, 
      FilterToAlu_281, FilterToAlu_280, FilterToAlu_279, FilterToAlu_278, 
      FilterToAlu_277, FilterToAlu_276, FilterToAlu_275, FilterToAlu_274, 
      FilterToAlu_273, FilterToAlu_272, FilterToAlu_271, FilterToAlu_270, 
      FilterToAlu_269, FilterToAlu_268, FilterToAlu_267, FilterToAlu_266, 
      FilterToAlu_265, FilterToAlu_264, FilterToAlu_263, FilterToAlu_262, 
      FilterToAlu_261, FilterToAlu_260, FilterToAlu_259, FilterToAlu_258, 
      FilterToAlu_257, FilterToAlu_256, FilterToAlu_255, FilterToAlu_254, 
      FilterToAlu_253, FilterToAlu_252, FilterToAlu_251, FilterToAlu_250, 
      FilterToAlu_249, FilterToAlu_248, FilterToAlu_247, FilterToAlu_246, 
      FilterToAlu_245, FilterToAlu_244, FilterToAlu_243, FilterToAlu_242, 
      FilterToAlu_241, FilterToAlu_240, FilterToAlu_239, FilterToAlu_238, 
      FilterToAlu_237, FilterToAlu_236, FilterToAlu_235, FilterToAlu_234, 
      FilterToAlu_233, FilterToAlu_232, FilterToAlu_231, FilterToAlu_230, 
      FilterToAlu_229, FilterToAlu_228, FilterToAlu_227, FilterToAlu_226, 
      FilterToAlu_225, FilterToAlu_224, FilterToAlu_223, FilterToAlu_222, 
      FilterToAlu_221, FilterToAlu_220, FilterToAlu_219, FilterToAlu_218, 
      FilterToAlu_217, FilterToAlu_216, FilterToAlu_215, FilterToAlu_214, 
      FilterToAlu_213, FilterToAlu_212, FilterToAlu_211, FilterToAlu_210, 
      FilterToAlu_209, FilterToAlu_208, FilterToAlu_207, FilterToAlu_206, 
      FilterToAlu_205, FilterToAlu_204, FilterToAlu_203, FilterToAlu_202, 
      FilterToAlu_201, FilterToAlu_200, FilterToAlu_199, FilterToAlu_198, 
      FilterToAlu_197, FilterToAlu_196, FilterToAlu_195, FilterToAlu_194, 
      FilterToAlu_193, FilterToAlu_192, FilterToAlu_191, FilterToAlu_190, 
      FilterToAlu_189, FilterToAlu_188, FilterToAlu_187, FilterToAlu_186, 
      FilterToAlu_185, FilterToAlu_184, FilterToAlu_183, FilterToAlu_182, 
      FilterToAlu_181, FilterToAlu_180, FilterToAlu_179, FilterToAlu_178, 
      FilterToAlu_177, FilterToAlu_176, FilterToAlu_175, FilterToAlu_174, 
      FilterToAlu_173, FilterToAlu_172, FilterToAlu_171, FilterToAlu_170, 
      FilterToAlu_169, FilterToAlu_168, FilterToAlu_167, FilterToAlu_166, 
      FilterToAlu_165, FilterToAlu_164, FilterToAlu_163, FilterToAlu_162, 
      FilterToAlu_161, FilterToAlu_160, FilterToAlu_159, FilterToAlu_158, 
      FilterToAlu_157, FilterToAlu_156, FilterToAlu_155, FilterToAlu_154, 
      FilterToAlu_153, FilterToAlu_152, FilterToAlu_151, FilterToAlu_150, 
      FilterToAlu_149, FilterToAlu_148, FilterToAlu_147, FilterToAlu_146, 
      FilterToAlu_145, FilterToAlu_144, FilterToAlu_143, FilterToAlu_142, 
      FilterToAlu_141, FilterToAlu_140, FilterToAlu_139, FilterToAlu_138, 
      FilterToAlu_137, FilterToAlu_136, FilterToAlu_135, FilterToAlu_134, 
      FilterToAlu_133, FilterToAlu_132, FilterToAlu_131, FilterToAlu_130, 
      FilterToAlu_129, FilterToAlu_128, FilterToAlu_127, FilterToAlu_126, 
      FilterToAlu_125, FilterToAlu_124, FilterToAlu_123, FilterToAlu_122, 
      FilterToAlu_121, FilterToAlu_120, FilterToAlu_119, FilterToAlu_118, 
      FilterToAlu_117, FilterToAlu_116, FilterToAlu_115, FilterToAlu_114, 
      FilterToAlu_113, FilterToAlu_112, FilterToAlu_111, FilterToAlu_110, 
      FilterToAlu_109, FilterToAlu_108, FilterToAlu_107, FilterToAlu_106, 
      FilterToAlu_105, FilterToAlu_104, FilterToAlu_103, FilterToAlu_102, 
      FilterToAlu_101, FilterToAlu_100, FilterToAlu_99, FilterToAlu_98, 
      FilterToAlu_97, FilterToAlu_96, FilterToAlu_95, FilterToAlu_94, 
      FilterToAlu_93, FilterToAlu_92, FilterToAlu_91, FilterToAlu_90, 
      FilterToAlu_89, FilterToAlu_88, FilterToAlu_87, FilterToAlu_86, 
      FilterToAlu_85, FilterToAlu_84, FilterToAlu_83, FilterToAlu_82, 
      FilterToAlu_81, FilterToAlu_80, FilterToAlu_79, FilterToAlu_78, 
      FilterToAlu_77, FilterToAlu_76, FilterToAlu_75, FilterToAlu_74, 
      FilterToAlu_73, FilterToAlu_72, FilterToAlu_71, FilterToAlu_70, 
      FilterToAlu_69, FilterToAlu_68, FilterToAlu_67, FilterToAlu_66, 
      FilterToAlu_65, FilterToAlu_64, FilterToAlu_63, FilterToAlu_62, 
      FilterToAlu_61, FilterToAlu_60, FilterToAlu_59, FilterToAlu_58, 
      FilterToAlu_57, FilterToAlu_56, FilterToAlu_55, FilterToAlu_54, 
      FilterToAlu_53, FilterToAlu_52, FilterToAlu_51, FilterToAlu_50, 
      FilterToAlu_49, FilterToAlu_48, FilterToAlu_47, FilterToAlu_46, 
      FilterToAlu_45, FilterToAlu_44, FilterToAlu_43, FilterToAlu_42, 
      FilterToAlu_41, FilterToAlu_40, FilterToAlu_39, FilterToAlu_38, 
      FilterToAlu_37, FilterToAlu_36, FilterToAlu_35, FilterToAlu_34, 
      FilterToAlu_33, FilterToAlu_32, FilterToAlu_31, FilterToAlu_30, 
      FilterToAlu_29, FilterToAlu_28, FilterToAlu_27, FilterToAlu_26, 
      FilterToAlu_25, FilterToAlu_24, FilterToAlu_23, FilterToAlu_22, 
      FilterToAlu_21, FilterToAlu_20, FilterToAlu_19, FilterToAlu_18, 
      FilterToAlu_17, FilterToAlu_16, FilterToAlu_15, FilterToAlu_14, 
      FilterToAlu_13, FilterToAlu_12, FilterToAlu_11, FilterToAlu_10, 
      FilterToAlu_9, FilterToAlu_8, FilterToAlu_7, FilterToAlu_6, 
      FilterToAlu_5, FilterToAlu_4, FilterToAlu_3, FilterToAlu_2, 
      FilterToAlu_1, FilterToAlu_0, MultiplierOut_792, MultiplierOut_791, 
      MultiplierOut_790, MultiplierOut_789, MultiplierOut_788, 
      MultiplierOut_787, MultiplierOut_786, MultiplierOut_785, 
      MultiplierOut_784, MultiplierOut_783, MultiplierOut_782, 
      MultiplierOut_781, MultiplierOut_780, MultiplierOut_779, 
      MultiplierOut_778, MultiplierOut_777, MultiplierOut_760, 
      MultiplierOut_759, MultiplierOut_758, MultiplierOut_757, 
      MultiplierOut_756, MultiplierOut_755, MultiplierOut_754, 
      MultiplierOut_753, MultiplierOut_752, MultiplierOut_751, 
      MultiplierOut_750, MultiplierOut_749, MultiplierOut_748, 
      MultiplierOut_747, MultiplierOut_746, MultiplierOut_745, 
      MultiplierOut_728, MultiplierOut_727, MultiplierOut_726, 
      MultiplierOut_725, MultiplierOut_724, MultiplierOut_723, 
      MultiplierOut_722, MultiplierOut_721, MultiplierOut_720, 
      MultiplierOut_719, MultiplierOut_718, MultiplierOut_717, 
      MultiplierOut_716, MultiplierOut_715, MultiplierOut_714, 
      MultiplierOut_713, MultiplierOut_696, MultiplierOut_695, 
      MultiplierOut_694, MultiplierOut_693, MultiplierOut_692, 
      MultiplierOut_691, MultiplierOut_690, MultiplierOut_689, 
      MultiplierOut_688, MultiplierOut_687, MultiplierOut_686, 
      MultiplierOut_685, MultiplierOut_684, MultiplierOut_683, 
      MultiplierOut_682, MultiplierOut_681, MultiplierOut_664, 
      MultiplierOut_663, MultiplierOut_662, MultiplierOut_661, 
      MultiplierOut_660, MultiplierOut_659, MultiplierOut_658, 
      MultiplierOut_657, MultiplierOut_656, MultiplierOut_655, 
      MultiplierOut_654, MultiplierOut_653, MultiplierOut_652, 
      MultiplierOut_651, MultiplierOut_650, MultiplierOut_649, 
      MultiplierOut_632, MultiplierOut_631, MultiplierOut_630, 
      MultiplierOut_629, MultiplierOut_628, MultiplierOut_627, 
      MultiplierOut_626, MultiplierOut_625, MultiplierOut_624, 
      MultiplierOut_623, MultiplierOut_622, MultiplierOut_621, 
      MultiplierOut_620, MultiplierOut_619, MultiplierOut_618, 
      MultiplierOut_617, MultiplierOut_600, MultiplierOut_599, 
      MultiplierOut_598, MultiplierOut_597, MultiplierOut_596, 
      MultiplierOut_595, MultiplierOut_594, MultiplierOut_593, 
      MultiplierOut_592, MultiplierOut_591, MultiplierOut_590, 
      MultiplierOut_589, MultiplierOut_588, MultiplierOut_587, 
      MultiplierOut_586, MultiplierOut_585, MultiplierOut_568, 
      MultiplierOut_567, MultiplierOut_566, MultiplierOut_565, 
      MultiplierOut_564, MultiplierOut_563, MultiplierOut_562, 
      MultiplierOut_561, MultiplierOut_560, MultiplierOut_559, 
      MultiplierOut_558, MultiplierOut_557, MultiplierOut_556, 
      MultiplierOut_555, MultiplierOut_554, MultiplierOut_553, 
      MultiplierOut_536, MultiplierOut_535, MultiplierOut_534, 
      MultiplierOut_533, MultiplierOut_532, MultiplierOut_531, 
      MultiplierOut_530, MultiplierOut_529, MultiplierOut_528, 
      MultiplierOut_527, MultiplierOut_526, MultiplierOut_525, 
      MultiplierOut_524, MultiplierOut_523, MultiplierOut_522, 
      MultiplierOut_521, MultiplierOut_504, MultiplierOut_503, 
      MultiplierOut_502, MultiplierOut_501, MultiplierOut_500, 
      MultiplierOut_499, MultiplierOut_498, MultiplierOut_497, 
      MultiplierOut_496, MultiplierOut_495, MultiplierOut_494, 
      MultiplierOut_493, MultiplierOut_492, MultiplierOut_491, 
      MultiplierOut_490, MultiplierOut_489, MultiplierOut_472, 
      MultiplierOut_471, MultiplierOut_470, MultiplierOut_469, 
      MultiplierOut_468, MultiplierOut_467, MultiplierOut_466, 
      MultiplierOut_465, MultiplierOut_464, MultiplierOut_463, 
      MultiplierOut_462, MultiplierOut_461, MultiplierOut_460, 
      MultiplierOut_459, MultiplierOut_458, MultiplierOut_457, 
      MultiplierOut_440, MultiplierOut_439, MultiplierOut_438, 
      MultiplierOut_437, MultiplierOut_436, MultiplierOut_435, 
      MultiplierOut_434, MultiplierOut_433, MultiplierOut_432, 
      MultiplierOut_431, MultiplierOut_430, MultiplierOut_429, 
      MultiplierOut_428, MultiplierOut_427, MultiplierOut_426, 
      MultiplierOut_425, MultiplierOut_408, MultiplierOut_407, 
      MultiplierOut_406, MultiplierOut_405, MultiplierOut_404, 
      MultiplierOut_403, MultiplierOut_402, MultiplierOut_401, 
      MultiplierOut_400, MultiplierOut_399, MultiplierOut_398, 
      MultiplierOut_397, MultiplierOut_396, MultiplierOut_395, 
      MultiplierOut_394, MultiplierOut_393, MultiplierOut_376, 
      MultiplierOut_375, MultiplierOut_374, MultiplierOut_373, 
      MultiplierOut_372, MultiplierOut_371, MultiplierOut_370, 
      MultiplierOut_369, MultiplierOut_368, MultiplierOut_367, 
      MultiplierOut_366, MultiplierOut_365, MultiplierOut_364, 
      MultiplierOut_363, MultiplierOut_362, MultiplierOut_361, 
      MultiplierOut_344, MultiplierOut_343, MultiplierOut_342, 
      MultiplierOut_341, MultiplierOut_340, MultiplierOut_339, 
      MultiplierOut_338, MultiplierOut_337, MultiplierOut_336, 
      MultiplierOut_335, MultiplierOut_334, MultiplierOut_333, 
      MultiplierOut_332, MultiplierOut_331, MultiplierOut_330, 
      MultiplierOut_329, MultiplierOut_312, MultiplierOut_311, 
      MultiplierOut_310, MultiplierOut_309, MultiplierOut_308, 
      MultiplierOut_307, MultiplierOut_306, MultiplierOut_305, 
      MultiplierOut_304, MultiplierOut_303, MultiplierOut_302, 
      MultiplierOut_301, MultiplierOut_300, MultiplierOut_299, 
      MultiplierOut_298, MultiplierOut_297, MultiplierOut_280, 
      MultiplierOut_279, MultiplierOut_278, MultiplierOut_277, 
      MultiplierOut_276, MultiplierOut_275, MultiplierOut_274, 
      MultiplierOut_273, MultiplierOut_272, MultiplierOut_271, 
      MultiplierOut_270, MultiplierOut_269, MultiplierOut_268, 
      MultiplierOut_267, MultiplierOut_266, MultiplierOut_265, 
      MultiplierOut_248, MultiplierOut_247, MultiplierOut_246, 
      MultiplierOut_245, MultiplierOut_244, MultiplierOut_243, 
      MultiplierOut_242, MultiplierOut_241, MultiplierOut_240, 
      MultiplierOut_239, MultiplierOut_238, MultiplierOut_237, 
      MultiplierOut_236, MultiplierOut_235, MultiplierOut_234, 
      MultiplierOut_233, MultiplierOut_216, MultiplierOut_215, 
      MultiplierOut_214, MultiplierOut_213, MultiplierOut_212, 
      MultiplierOut_211, MultiplierOut_210, MultiplierOut_209, 
      MultiplierOut_208, MultiplierOut_207, MultiplierOut_206, 
      MultiplierOut_205, MultiplierOut_204, MultiplierOut_203, 
      MultiplierOut_202, MultiplierOut_201, MultiplierOut_184, 
      MultiplierOut_183, MultiplierOut_182, MultiplierOut_181, 
      MultiplierOut_180, MultiplierOut_179, MultiplierOut_178, 
      MultiplierOut_177, MultiplierOut_176, MultiplierOut_175, 
      MultiplierOut_174, MultiplierOut_173, MultiplierOut_172, 
      MultiplierOut_171, MultiplierOut_170, MultiplierOut_169, 
      MultiplierOut_152, MultiplierOut_151, MultiplierOut_150, 
      MultiplierOut_149, MultiplierOut_148, MultiplierOut_147, 
      MultiplierOut_146, MultiplierOut_145, MultiplierOut_144, 
      MultiplierOut_143, MultiplierOut_142, MultiplierOut_141, 
      MultiplierOut_140, MultiplierOut_139, MultiplierOut_138, 
      MultiplierOut_137, MultiplierOut_120, MultiplierOut_119, 
      MultiplierOut_118, MultiplierOut_117, MultiplierOut_116, 
      MultiplierOut_115, MultiplierOut_114, MultiplierOut_113, 
      MultiplierOut_112, MultiplierOut_111, MultiplierOut_110, 
      MultiplierOut_109, MultiplierOut_108, MultiplierOut_107, 
      MultiplierOut_106, MultiplierOut_105, MultiplierOut_88, 
      MultiplierOut_87, MultiplierOut_86, MultiplierOut_85, MultiplierOut_84, 
      MultiplierOut_83, MultiplierOut_82, MultiplierOut_81, MultiplierOut_80, 
      MultiplierOut_79, MultiplierOut_78, MultiplierOut_77, MultiplierOut_76, 
      MultiplierOut_75, MultiplierOut_74, MultiplierOut_73, MultiplierOut_56, 
      MultiplierOut_55, MultiplierOut_54, MultiplierOut_53, MultiplierOut_52, 
      MultiplierOut_51, MultiplierOut_50, MultiplierOut_49, MultiplierOut_48, 
      MultiplierOut_47, MultiplierOut_46, MultiplierOut_45, MultiplierOut_44, 
      MultiplierOut_43, MultiplierOut_42, MultiplierOut_41, MultiplierOut_24, 
      MultiplierOut_23, MultiplierOut_22, MultiplierOut_21, MultiplierOut_20, 
      MultiplierOut_19, MultiplierOut_18, MultiplierOut_17, MultiplierOut_16, 
      MultiplierOut_15, MultiplierOut_14, MultiplierOut_13, MultiplierOut_12, 
      MultiplierOut_11, MultiplierOut_10, MultiplierOut_9, AddOutputLvL1_191, 
      AddOutputLvL1_190, AddOutputLvL1_189, AddOutputLvL1_188, 
      AddOutputLvL1_187, AddOutputLvL1_186, AddOutputLvL1_185, 
      AddOutputLvL1_184, AddOutputLvL1_183, AddOutputLvL1_182, 
      AddOutputLvL1_181, AddOutputLvL1_180, AddOutputLvL1_179, 
      AddOutputLvL1_178, AddOutputLvL1_177, AddOutputLvL1_176, 
      AddOutputLvL1_175, AddOutputLvL1_174, AddOutputLvL1_173, 
      AddOutputLvL1_172, AddOutputLvL1_171, AddOutputLvL1_170, 
      AddOutputLvL1_169, AddOutputLvL1_168, AddOutputLvL1_167, 
      AddOutputLvL1_166, AddOutputLvL1_165, AddOutputLvL1_164, 
      AddOutputLvL1_163, AddOutputLvL1_162, AddOutputLvL1_161, 
      AddOutputLvL1_160, AddOutputLvL1_159, AddOutputLvL1_158, 
      AddOutputLvL1_157, AddOutputLvL1_156, AddOutputLvL1_155, 
      AddOutputLvL1_154, AddOutputLvL1_153, AddOutputLvL1_152, 
      AddOutputLvL1_151, AddOutputLvL1_150, AddOutputLvL1_149, 
      AddOutputLvL1_148, AddOutputLvL1_147, AddOutputLvL1_146, 
      AddOutputLvL1_145, AddOutputLvL1_144, AddOutputLvL1_143, 
      AddOutputLvL1_142, AddOutputLvL1_141, AddOutputLvL1_140, 
      AddOutputLvL1_139, AddOutputLvL1_138, AddOutputLvL1_137, 
      AddOutputLvL1_136, AddOutputLvL1_135, AddOutputLvL1_134, 
      AddOutputLvL1_133, AddOutputLvL1_132, AddOutputLvL1_131, 
      AddOutputLvL1_130, AddOutputLvL1_129, AddOutputLvL1_128, 
      AddOutputLvL1_127, AddOutputLvL1_126, AddOutputLvL1_125, 
      AddOutputLvL1_124, AddOutputLvL1_123, AddOutputLvL1_122, 
      AddOutputLvL1_121, AddOutputLvL1_120, AddOutputLvL1_119, 
      AddOutputLvL1_118, AddOutputLvL1_117, AddOutputLvL1_116, 
      AddOutputLvL1_115, AddOutputLvL1_114, AddOutputLvL1_113, 
      AddOutputLvL1_112, AddOutputLvL1_111, AddOutputLvL1_110, 
      AddOutputLvL1_109, AddOutputLvL1_108, AddOutputLvL1_107, 
      AddOutputLvL1_106, AddOutputLvL1_105, AddOutputLvL1_104, 
      AddOutputLvL1_103, AddOutputLvL1_102, AddOutputLvL1_101, 
      AddOutputLvL1_100, AddOutputLvL1_99, AddOutputLvL1_98, 
      AddOutputLvL1_97, AddOutputLvL1_96, AddOutputLvL1_95, AddOutputLvL1_94, 
      AddOutputLvL1_93, AddOutputLvL1_92, AddOutputLvL1_91, AddOutputLvL1_90, 
      AddOutputLvL1_89, AddOutputLvL1_88, AddOutputLvL1_87, AddOutputLvL1_86, 
      AddOutputLvL1_85, AddOutputLvL1_84, AddOutputLvL1_83, AddOutputLvL1_82, 
      AddOutputLvL1_81, AddOutputLvL1_80, AddOutputLvL1_79, AddOutputLvL1_78, 
      AddOutputLvL1_77, AddOutputLvL1_76, AddOutputLvL1_75, AddOutputLvL1_74, 
      AddOutputLvL1_73, AddOutputLvL1_72, AddOutputLvL1_71, AddOutputLvL1_70, 
      AddOutputLvL1_69, AddOutputLvL1_68, AddOutputLvL1_67, AddOutputLvL1_66, 
      AddOutputLvL1_65, AddOutputLvL1_64, AddOutputLvL1_63, AddOutputLvL1_62, 
      AddOutputLvL1_61, AddOutputLvL1_60, AddOutputLvL1_59, AddOutputLvL1_58, 
      AddOutputLvL1_57, AddOutputLvL1_56, AddOutputLvL1_55, AddOutputLvL1_54, 
      AddOutputLvL1_53, AddOutputLvL1_52, AddOutputLvL1_51, AddOutputLvL1_50, 
      AddOutputLvL1_49, AddOutputLvL1_48, AddOutputLvL1_47, AddOutputLvL1_46, 
      AddOutputLvL1_45, AddOutputLvL1_44, AddOutputLvL1_43, AddOutputLvL1_42, 
      AddOutputLvL1_41, AddOutputLvL1_40, AddOutputLvL1_39, AddOutputLvL1_38, 
      AddOutputLvL1_37, AddOutputLvL1_36, AddOutputLvL1_35, AddOutputLvL1_34, 
      AddOutputLvL1_33, AddOutputLvL1_32, AddOutputLvL1_31, AddOutputLvL1_30, 
      AddOutputLvL1_29, AddOutputLvL1_28, AddOutputLvL1_27, AddOutputLvL1_26, 
      AddOutputLvL1_25, AddOutputLvL1_24, AddOutputLvL1_23, AddOutputLvL1_22, 
      AddOutputLvL1_21, AddOutputLvL1_20, AddOutputLvL1_19, AddOutputLvL1_18, 
      AddOutputLvL1_17, AddOutputLvL1_16, AddOutputLvL1_15, AddOutputLvL1_14, 
      AddOutputLvL1_13, AddOutputLvL1_12, AddOutputLvL1_11, AddOutputLvL1_10, 
      AddOutputLvL1_9, AddOutputLvL1_8, AddOutputLvL1_7, AddOutputLvL1_6, 
      AddOutputLvL1_5, AddOutputLvL1_4, AddOutputLvL1_3, AddOutputLvL1_2, 
      AddOutputLvL1_1, AddOutputLvL1_0, AddOutputLvL2_95, AddOutputLvL2_94, 
      AddOutputLvL2_93, AddOutputLvL2_92, AddOutputLvL2_91, AddOutputLvL2_90, 
      AddOutputLvL2_89, AddOutputLvL2_88, AddOutputLvL2_87, AddOutputLvL2_86, 
      AddOutputLvL2_85, AddOutputLvL2_84, AddOutputLvL2_83, AddOutputLvL2_82, 
      AddOutputLvL2_81, AddOutputLvL2_80, AddOutputLvL2_79, AddOutputLvL2_78, 
      AddOutputLvL2_77, AddOutputLvL2_76, AddOutputLvL2_75, AddOutputLvL2_74, 
      AddOutputLvL2_73, AddOutputLvL2_72, AddOutputLvL2_71, AddOutputLvL2_70, 
      AddOutputLvL2_69, AddOutputLvL2_68, AddOutputLvL2_67, AddOutputLvL2_66, 
      AddOutputLvL2_65, AddOutputLvL2_64, AddOutputLvL2_63, AddOutputLvL2_62, 
      AddOutputLvL2_61, AddOutputLvL2_60, AddOutputLvL2_59, AddOutputLvL2_58, 
      AddOutputLvL2_57, AddOutputLvL2_56, AddOutputLvL2_55, AddOutputLvL2_54, 
      AddOutputLvL2_53, AddOutputLvL2_52, AddOutputLvL2_51, AddOutputLvL2_50, 
      AddOutputLvL2_49, AddOutputLvL2_48, AddOutputLvL2_47, AddOutputLvL2_46, 
      AddOutputLvL2_45, AddOutputLvL2_44, AddOutputLvL2_43, AddOutputLvL2_42, 
      AddOutputLvL2_41, AddOutputLvL2_40, AddOutputLvL2_39, AddOutputLvL2_38, 
      AddOutputLvL2_37, AddOutputLvL2_36, AddOutputLvL2_35, AddOutputLvL2_34, 
      AddOutputLvL2_33, AddOutputLvL2_32, AddOutputLvL2_31, AddOutputLvL2_30, 
      AddOutputLvL2_29, AddOutputLvL2_28, AddOutputLvL2_27, AddOutputLvL2_26, 
      AddOutputLvL2_25, AddOutputLvL2_24, AddOutputLvL2_23, AddOutputLvL2_22, 
      AddOutputLvL2_21, AddOutputLvL2_20, AddOutputLvL2_19, AddOutputLvL2_18, 
      AddOutputLvL2_17, AddOutputLvL2_16, AddOutputLvL2_15, AddOutputLvL2_14, 
      AddOutputLvL2_13, AddOutputLvL2_12, AddOutputLvL2_11, AddOutputLvL2_10, 
      AddOutputLvL2_9, AddOutputLvL2_8, AddOutputLvL2_7, AddOutputLvL2_6, 
      AddOutputLvL2_5, AddOutputLvL2_4, AddOutputLvL2_3, AddOutputLvL2_2, 
      AddOutputLvL2_1, AddOutputLvL2_0, AddOutputLvL3_47, AddOutputLvL3_46, 
      AddOutputLvL3_45, AddOutputLvL3_44, AddOutputLvL3_43, AddOutputLvL3_42, 
      AddOutputLvL3_41, AddOutputLvL3_40, AddOutputLvL3_39, AddOutputLvL3_38, 
      AddOutputLvL3_37, AddOutputLvL3_36, AddOutputLvL3_35, AddOutputLvL3_34, 
      AddOutputLvL3_33, AddOutputLvL3_32, AddOutputLvL3_31, AddOutputLvL3_30, 
      AddOutputLvL3_29, AddOutputLvL3_28, AddOutputLvL3_27, AddOutputLvL3_26, 
      AddOutputLvL3_25, AddOutputLvL3_24, AddOutputLvL3_23, AddOutputLvL3_22, 
      AddOutputLvL3_21, AddOutputLvL3_20, AddOutputLvL3_19, AddOutputLvL3_18, 
      AddOutputLvL3_17, AddOutputLvL3_16, AddOutputLvL3_15, AddOutputLvL3_14, 
      AddOutputLvL3_13, AddOutputLvL3_12, AddOutputLvL3_11, AddOutputLvL3_10, 
      AddOutputLvL3_9, AddOutputLvL3_8, AddOutputLvL3_7, AddOutputLvL3_6, 
      AddOutputLvL3_5, AddOutputLvL3_4, AddOutputLvL3_3, AddOutputLvL3_2, 
      AddOutputLvL3_1, AddOutputLvL3_0, AddOut33_15, AddOut33_14, 
      AddOut33_13, AddOut33_12, AddOut33_11, AddOut33_10, AddOut33_9, 
      AddOut33_8, AddOut33_7, AddOut33_6, AddOut33_5, AddOut33_4, AddOut33_3, 
      AddOut33_2, AddOut33_1, AddOut33_0, AddOut55_15, AddOut55_14, 
      AddOut55_13, AddOut55_12, AddOut55_11, AddOut55_10, AddOut55_9, 
      AddOut55_8, AddOut55_7, AddOut55_6, AddOut55_5, AddOut55_4, AddOut55_3, 
      AddOut55_2, AddOut55_1, AddOut55_0, Final55_15, Final55_14, Final55_13, 
      Final55_12, Final55_11, Final55_10, Final55_9, Final55_8, Final55_7, 
      Final55_6, Final55_5, Final55_4, Final55_3, Final55_2, Final55_1, 
      Final55_0, CounterOut_2, CounterOut_1, CounterOut_0, 
      SecondInputToMult_143, SecondInputToMult_142, SecondInputToMult_141, 
      SecondInputToMult_140, SecondInputToMult_139, SecondInputToMult_138, 
      SecondInputToMult_137, SecondInputToMult_136, SecondInputToMult_135, 
      SecondInputToMult_134, SecondInputToMult_133, SecondInputToMult_132, 
      SecondInputToMult_131, SecondInputToMult_130, SecondInputToMult_129, 
      SecondInputToMult_128, SecondInputToMult_127, SecondInputToMult_126, 
      SecondInputToMult_125, SecondInputToMult_124, SecondInputToMult_123, 
      SecondInputToMult_122, SecondInputToMult_121, SecondInputToMult_120, 
      SecondInputToMult_119, SecondInputToMult_118, SecondInputToMult_117, 
      SecondInputToMult_116, SecondInputToMult_115, SecondInputToMult_114, 
      SecondInputToMult_113, SecondInputToMult_112, SecondInputToMult_111, 
      SecondInputToMult_110, SecondInputToMult_109, SecondInputToMult_108, 
      SecondInputToMult_107, SecondInputToMult_106, SecondInputToMult_105, 
      SecondInputToMult_104, SecondInputToMult_103, SecondInputToMult_102, 
      SecondInputToMult_101, SecondInputToMult_100, SecondInputToMult_99, 
      SecondInputToMult_98, SecondInputToMult_97, SecondInputToMult_96, 
      SecondInputToMult_95, SecondInputToMult_94, SecondInputToMult_93, 
      SecondInputToMult_92, SecondInputToMult_91, SecondInputToMult_90, 
      SecondInputToMult_89, SecondInputToMult_88, SecondInputToMult_87, 
      SecondInputToMult_86, SecondInputToMult_85, SecondInputToMult_84, 
      SecondInputToMult_83, SecondInputToMult_82, SecondInputToMult_81, 
      SecondInputToMult_80, SecondInputToMult_79, SecondInputToMult_78, 
      SecondInputToMult_77, SecondInputToMult_76, SecondInputToMult_75, 
      SecondInputToMult_74, SecondInputToMult_73, SecondInputToMult_72, 
      SecondInputToMult_71, SecondInputToMult_70, SecondInputToMult_69, 
      SecondInputToMult_68, SecondInputToMult_67, SecondInputToMult_66, 
      SecondInputToMult_65, SecondInputToMult_64, SecondInputToMult_63, 
      SecondInputToMult_62, SecondInputToMult_61, SecondInputToMult_60, 
      SecondInputToMult_59, SecondInputToMult_58, SecondInputToMult_57, 
      SecondInputToMult_56, SecondInputToMult_55, SecondInputToMult_54, 
      SecondInputToMult_53, SecondInputToMult_52, SecondInputToMult_51, 
      SecondInputToMult_50, SecondInputToMult_49, SecondInputToMult_48, 
      CountereEN, CountereRST, GND0, nx6, nx12, nx20, nx32, nx34, nx48, nx68, 
      nx98, nx116, nx134, nx152, nx170, nx188, nx206, nx224, nx510, nx516, 
      nx3552, nx3562, nx7936, nx8052, nx8072, nx8090, nx8108, nx8126, nx8144, 
      nx8162, nx8180, nx8198, nx8216, nx8234, nx8252, nx8270, nx8288, nx8306, 
      nx8324, nx8342, nx8360, nx8378, nx8396, nx8414, nx8432, nx8450, nx8468, 
      nx8486, nx8495, nx8501, nx8511, nx8514, nx8517, nx8520, nx8523, nx8525, 
      nx8528, nx8530, nx8534, nx8536, nx8540, nx8542, nx8546, nx8548, nx8552, 
      nx8554, nx8558, nx8560, nx8564, nx8566, nx8569, nx8571, nx8586, nx8588, 
      nx8590, nx8592, nx8594, nx8596, nx8598, nx8600, nx8602, nx8604, nx8606, 
      nx8608, nx8610, nx8612, nx8614, nx8616, nx8618, nx8620, nx8622, nx8624, 
      nx8626, nx8628, nx8630, nx8632, nx8634, nx8636, nx8638, nx8640, nx8642, 
      nx8644, nx8646, nx8648, nx8650, nx8652, nx8654, nx8656, nx8658, nx8660, 
      nx8662, nx8664, nx8666, nx8668, nx8670, nx8672, nx8674, nx8676, nx8678, 
      nx8680, nx8682, nx8684, nx8686, nx8688, nx8690, nx8692, nx8696, nx8698, 
      nx8700, nx8702, nx8704, nx8706, nx8708, nx8710, nx8712, nx8714, nx8716, 
      nx8718, nx8720, nx8722, nx8724, nx8726, nx8728, nx8730, nx8732, nx8734, 
      nx8736, nx8738, nx8740, nx8742, nx8744, nx8746, nx8748, nx8750, nx8752, 
      nx8754, nx8756, nx8758, nx8760, nx8762, nx8764, nx8766, nx8768, nx8770, 
      nx8772, nx8774, nx8776, nx8778, nx8780, nx8782, nx8784, nx8786, nx8788, 
      nx8790, nx8792, nx8794, nx8796, nx8798, nx8800, nx8802, nx8804, nx8806, 
      nx8808, nx8810, nx8812, nx8814, nx8816, nx8818, nx8820, nx8822, nx8824, 
      nx8826, nx8828, nx8830, nx8832, nx8834, nx8836, nx8838, nx8840, nx8842, 
      nx8844, nx8846, nx8852, nx8854, nx8856, nx8858, nx8860, nx8862, nx8864, 
      nx8866, nx8868, nx8870, nx8872, nx8874, nx8876, nx8878, nx8880, nx8882, 
      nx8884, nx8886, nx8888, nx8890, nx8892, nx8894, nx8896, nx8898, nx8900, 
      nx8902, nx8904, nx8906, nx8908, nx8910, nx8912, nx8914, nx8916, nx8918, 
      nx8920, nx8922, nx8924, nx8926: std_logic ;
   
   signal DANGLING : std_logic_vector (423 downto 0 );

begin
   ACK <= ACK_EXMPLR ;
   ConvOuput(15) <= ConvOuput_15_EXMPLR ;
   loop3_0_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_15, A(14)=>
      FilterToAlu_14, A(13)=>FilterToAlu_13, A(12)=>FilterToAlu_12, A(11)=>
      FilterToAlu_11, A(10)=>FilterToAlu_10, A(9)=>FilterToAlu_9, A(8)=>
      FilterToAlu_8, A(7)=>FilterToAlu_7, A(6)=>FilterToAlu_6, A(5)=>
      FilterToAlu_5, A(4)=>FilterToAlu_4, A(3)=>FilterToAlu_3, A(2)=>
      FilterToAlu_2, A(1)=>FilterToAlu_1, A(0)=>FilterToAlu_0, B(15)=>
      OutputImg0(15), B(14)=>OutputImg0(14), B(13)=>OutputImg0(13), B(12)=>
      OutputImg0(12), B(11)=>OutputImg0(11), B(10)=>OutputImg0(10), B(9)=>
      OutputImg0(9), B(8)=>OutputImg0(8), B(7)=>OutputImg0(7), B(6)=>
      OutputImg0(6), B(5)=>OutputImg0(5), B(4)=>OutputImg0(4), B(3)=>
      OutputImg0(3), B(2)=>OutputImg0(2), B(1)=>OutputImg0(1), B(0)=>
      OutputImg0(0), F(31)=>DANGLING(0), F(30)=>DANGLING(1), F(29)=>DANGLING
      (2), F(28)=>DANGLING(3), F(27)=>DANGLING(4), F(26)=>DANGLING(5), F(25)
      =>DANGLING(6), F(24)=>MultiplierOut_24, F(23)=>MultiplierOut_23, F(22)
      =>MultiplierOut_22, F(21)=>MultiplierOut_21, F(20)=>MultiplierOut_20, 
      F(19)=>MultiplierOut_19, F(18)=>MultiplierOut_18, F(17)=>
      MultiplierOut_17, F(16)=>MultiplierOut_16, F(15)=>MultiplierOut_15, 
      F(14)=>MultiplierOut_14, F(13)=>MultiplierOut_13, F(12)=>
      MultiplierOut_12, F(11)=>MultiplierOut_11, F(10)=>MultiplierOut_10, 
      F(9)=>MultiplierOut_9, F(8)=>DANGLING(7), F(7)=>DANGLING(8), F(6)=>
      DANGLING(9), F(5)=>DANGLING(10), F(4)=>DANGLING(11), F(3)=>DANGLING(12
      ), F(2)=>DANGLING(13), F(1)=>DANGLING(14), F(0)=>DANGLING(15));
   loop3_1_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_31, A(14)=>
      FilterToAlu_30, A(13)=>FilterToAlu_29, A(12)=>FilterToAlu_28, A(11)=>
      FilterToAlu_27, A(10)=>FilterToAlu_26, A(9)=>FilterToAlu_25, A(8)=>
      FilterToAlu_24, A(7)=>FilterToAlu_23, A(6)=>FilterToAlu_22, A(5)=>
      FilterToAlu_21, A(4)=>FilterToAlu_20, A(3)=>FilterToAlu_19, A(2)=>
      FilterToAlu_18, A(1)=>FilterToAlu_17, A(0)=>FilterToAlu_16, B(15)=>
      OutputImg0(31), B(14)=>OutputImg0(30), B(13)=>OutputImg0(29), B(12)=>
      OutputImg0(28), B(11)=>OutputImg0(27), B(10)=>OutputImg0(26), B(9)=>
      OutputImg0(25), B(8)=>OutputImg0(24), B(7)=>OutputImg0(23), B(6)=>
      OutputImg0(22), B(5)=>OutputImg0(21), B(4)=>OutputImg0(20), B(3)=>
      OutputImg0(19), B(2)=>OutputImg0(18), B(1)=>OutputImg0(17), B(0)=>
      OutputImg0(16), F(31)=>DANGLING(16), F(30)=>DANGLING(17), F(29)=>
      DANGLING(18), F(28)=>DANGLING(19), F(27)=>DANGLING(20), F(26)=>
      DANGLING(21), F(25)=>DANGLING(22), F(24)=>MultiplierOut_56, F(23)=>
      MultiplierOut_55, F(22)=>MultiplierOut_54, F(21)=>MultiplierOut_53, 
      F(20)=>MultiplierOut_52, F(19)=>MultiplierOut_51, F(18)=>
      MultiplierOut_50, F(17)=>MultiplierOut_49, F(16)=>MultiplierOut_48, 
      F(15)=>MultiplierOut_47, F(14)=>MultiplierOut_46, F(13)=>
      MultiplierOut_45, F(12)=>MultiplierOut_44, F(11)=>MultiplierOut_43, 
      F(10)=>MultiplierOut_42, F(9)=>MultiplierOut_41, F(8)=>DANGLING(23), 
      F(7)=>DANGLING(24), F(6)=>DANGLING(25), F(5)=>DANGLING(26), F(4)=>
      DANGLING(27), F(3)=>DANGLING(28), F(2)=>DANGLING(29), F(1)=>DANGLING(
      30), F(0)=>DANGLING(31));
   loop3_2_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_47, A(14)=>
      FilterToAlu_46, A(13)=>FilterToAlu_45, A(12)=>FilterToAlu_44, A(11)=>
      FilterToAlu_43, A(10)=>FilterToAlu_42, A(9)=>FilterToAlu_41, A(8)=>
      FilterToAlu_40, A(7)=>FilterToAlu_39, A(6)=>FilterToAlu_38, A(5)=>
      FilterToAlu_37, A(4)=>FilterToAlu_36, A(3)=>FilterToAlu_35, A(2)=>
      FilterToAlu_34, A(1)=>FilterToAlu_33, A(0)=>FilterToAlu_32, B(15)=>
      OutputImg0(47), B(14)=>OutputImg0(46), B(13)=>OutputImg0(45), B(12)=>
      OutputImg0(44), B(11)=>OutputImg0(43), B(10)=>OutputImg0(42), B(9)=>
      OutputImg0(41), B(8)=>OutputImg0(40), B(7)=>OutputImg0(39), B(6)=>
      OutputImg0(38), B(5)=>OutputImg0(37), B(4)=>OutputImg0(36), B(3)=>
      OutputImg0(35), B(2)=>OutputImg0(34), B(1)=>OutputImg0(33), B(0)=>
      OutputImg0(32), F(31)=>DANGLING(32), F(30)=>DANGLING(33), F(29)=>
      DANGLING(34), F(28)=>DANGLING(35), F(27)=>DANGLING(36), F(26)=>
      DANGLING(37), F(25)=>DANGLING(38), F(24)=>MultiplierOut_88, F(23)=>
      MultiplierOut_87, F(22)=>MultiplierOut_86, F(21)=>MultiplierOut_85, 
      F(20)=>MultiplierOut_84, F(19)=>MultiplierOut_83, F(18)=>
      MultiplierOut_82, F(17)=>MultiplierOut_81, F(16)=>MultiplierOut_80, 
      F(15)=>MultiplierOut_79, F(14)=>MultiplierOut_78, F(13)=>
      MultiplierOut_77, F(12)=>MultiplierOut_76, F(11)=>MultiplierOut_75, 
      F(10)=>MultiplierOut_74, F(9)=>MultiplierOut_73, F(8)=>DANGLING(39), 
      F(7)=>DANGLING(40), F(6)=>DANGLING(41), F(5)=>DANGLING(42), F(4)=>
      DANGLING(43), F(3)=>DANGLING(44), F(2)=>DANGLING(45), F(1)=>DANGLING(
      46), F(0)=>DANGLING(47));
   loop3_3_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_63, A(14)=>
      FilterToAlu_62, A(13)=>FilterToAlu_61, A(12)=>FilterToAlu_60, A(11)=>
      FilterToAlu_59, A(10)=>FilterToAlu_58, A(9)=>FilterToAlu_57, A(8)=>
      FilterToAlu_56, A(7)=>FilterToAlu_55, A(6)=>FilterToAlu_54, A(5)=>
      FilterToAlu_53, A(4)=>FilterToAlu_52, A(3)=>FilterToAlu_51, A(2)=>
      FilterToAlu_50, A(1)=>FilterToAlu_49, A(0)=>FilterToAlu_48, B(15)=>
      SecondInputToMult_63, B(14)=>SecondInputToMult_62, B(13)=>
      SecondInputToMult_61, B(12)=>SecondInputToMult_60, B(11)=>
      SecondInputToMult_59, B(10)=>SecondInputToMult_58, B(9)=>
      SecondInputToMult_57, B(8)=>SecondInputToMult_56, B(7)=>
      SecondInputToMult_55, B(6)=>SecondInputToMult_54, B(5)=>
      SecondInputToMult_53, B(4)=>SecondInputToMult_52, B(3)=>
      SecondInputToMult_51, B(2)=>SecondInputToMult_50, B(1)=>
      SecondInputToMult_49, B(0)=>SecondInputToMult_48, F(31)=>DANGLING(48), 
      F(30)=>DANGLING(49), F(29)=>DANGLING(50), F(28)=>DANGLING(51), F(27)=>
      DANGLING(52), F(26)=>DANGLING(53), F(25)=>DANGLING(54), F(24)=>
      MultiplierOut_120, F(23)=>MultiplierOut_119, F(22)=>MultiplierOut_118, 
      F(21)=>MultiplierOut_117, F(20)=>MultiplierOut_116, F(19)=>
      MultiplierOut_115, F(18)=>MultiplierOut_114, F(17)=>MultiplierOut_113, 
      F(16)=>MultiplierOut_112, F(15)=>MultiplierOut_111, F(14)=>
      MultiplierOut_110, F(13)=>MultiplierOut_109, F(12)=>MultiplierOut_108, 
      F(11)=>MultiplierOut_107, F(10)=>MultiplierOut_106, F(9)=>
      MultiplierOut_105, F(8)=>DANGLING(55), F(7)=>DANGLING(56), F(6)=>
      DANGLING(57), F(5)=>DANGLING(58), F(4)=>DANGLING(59), F(3)=>DANGLING(
      60), F(2)=>DANGLING(61), F(1)=>DANGLING(62), F(0)=>DANGLING(63));
   loop3_4_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_79, A(14)=>
      FilterToAlu_78, A(13)=>FilterToAlu_77, A(12)=>FilterToAlu_76, A(11)=>
      FilterToAlu_75, A(10)=>FilterToAlu_74, A(9)=>FilterToAlu_73, A(8)=>
      FilterToAlu_72, A(7)=>FilterToAlu_71, A(6)=>FilterToAlu_70, A(5)=>
      FilterToAlu_69, A(4)=>FilterToAlu_68, A(3)=>FilterToAlu_67, A(2)=>
      FilterToAlu_66, A(1)=>FilterToAlu_65, A(0)=>FilterToAlu_64, B(15)=>
      SecondInputToMult_79, B(14)=>SecondInputToMult_78, B(13)=>
      SecondInputToMult_77, B(12)=>SecondInputToMult_76, B(11)=>
      SecondInputToMult_75, B(10)=>SecondInputToMult_74, B(9)=>
      SecondInputToMult_73, B(8)=>SecondInputToMult_72, B(7)=>
      SecondInputToMult_71, B(6)=>SecondInputToMult_70, B(5)=>
      SecondInputToMult_69, B(4)=>SecondInputToMult_68, B(3)=>
      SecondInputToMult_67, B(2)=>SecondInputToMult_66, B(1)=>
      SecondInputToMult_65, B(0)=>SecondInputToMult_64, F(31)=>DANGLING(64), 
      F(30)=>DANGLING(65), F(29)=>DANGLING(66), F(28)=>DANGLING(67), F(27)=>
      DANGLING(68), F(26)=>DANGLING(69), F(25)=>DANGLING(70), F(24)=>
      MultiplierOut_152, F(23)=>MultiplierOut_151, F(22)=>MultiplierOut_150, 
      F(21)=>MultiplierOut_149, F(20)=>MultiplierOut_148, F(19)=>
      MultiplierOut_147, F(18)=>MultiplierOut_146, F(17)=>MultiplierOut_145, 
      F(16)=>MultiplierOut_144, F(15)=>MultiplierOut_143, F(14)=>
      MultiplierOut_142, F(13)=>MultiplierOut_141, F(12)=>MultiplierOut_140, 
      F(11)=>MultiplierOut_139, F(10)=>MultiplierOut_138, F(9)=>
      MultiplierOut_137, F(8)=>DANGLING(71), F(7)=>DANGLING(72), F(6)=>
      DANGLING(73), F(5)=>DANGLING(74), F(4)=>DANGLING(75), F(3)=>DANGLING(
      76), F(2)=>DANGLING(77), F(1)=>DANGLING(78), F(0)=>DANGLING(79));
   loop3_5_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_95, A(14)=>
      FilterToAlu_94, A(13)=>FilterToAlu_93, A(12)=>FilterToAlu_92, A(11)=>
      FilterToAlu_91, A(10)=>FilterToAlu_90, A(9)=>FilterToAlu_89, A(8)=>
      FilterToAlu_88, A(7)=>FilterToAlu_87, A(6)=>FilterToAlu_86, A(5)=>
      FilterToAlu_85, A(4)=>FilterToAlu_84, A(3)=>FilterToAlu_83, A(2)=>
      FilterToAlu_82, A(1)=>FilterToAlu_81, A(0)=>FilterToAlu_80, B(15)=>
      SecondInputToMult_95, B(14)=>SecondInputToMult_94, B(13)=>
      SecondInputToMult_93, B(12)=>SecondInputToMult_92, B(11)=>
      SecondInputToMult_91, B(10)=>SecondInputToMult_90, B(9)=>
      SecondInputToMult_89, B(8)=>SecondInputToMult_88, B(7)=>
      SecondInputToMult_87, B(6)=>SecondInputToMult_86, B(5)=>
      SecondInputToMult_85, B(4)=>SecondInputToMult_84, B(3)=>
      SecondInputToMult_83, B(2)=>SecondInputToMult_82, B(1)=>
      SecondInputToMult_81, B(0)=>SecondInputToMult_80, F(31)=>DANGLING(80), 
      F(30)=>DANGLING(81), F(29)=>DANGLING(82), F(28)=>DANGLING(83), F(27)=>
      DANGLING(84), F(26)=>DANGLING(85), F(25)=>DANGLING(86), F(24)=>
      MultiplierOut_184, F(23)=>MultiplierOut_183, F(22)=>MultiplierOut_182, 
      F(21)=>MultiplierOut_181, F(20)=>MultiplierOut_180, F(19)=>
      MultiplierOut_179, F(18)=>MultiplierOut_178, F(17)=>MultiplierOut_177, 
      F(16)=>MultiplierOut_176, F(15)=>MultiplierOut_175, F(14)=>
      MultiplierOut_174, F(13)=>MultiplierOut_173, F(12)=>MultiplierOut_172, 
      F(11)=>MultiplierOut_171, F(10)=>MultiplierOut_170, F(9)=>
      MultiplierOut_169, F(8)=>DANGLING(87), F(7)=>DANGLING(88), F(6)=>
      DANGLING(89), F(5)=>DANGLING(90), F(4)=>DANGLING(91), F(3)=>DANGLING(
      92), F(2)=>DANGLING(93), F(1)=>DANGLING(94), F(0)=>DANGLING(95));
   loop3_6_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_111, A(14)=>
      FilterToAlu_110, A(13)=>FilterToAlu_109, A(12)=>FilterToAlu_108, A(11)
      =>FilterToAlu_107, A(10)=>FilterToAlu_106, A(9)=>FilterToAlu_105, A(8)
      =>FilterToAlu_104, A(7)=>FilterToAlu_103, A(6)=>FilterToAlu_102, A(5)
      =>FilterToAlu_101, A(4)=>FilterToAlu_100, A(3)=>FilterToAlu_99, A(2)=>
      FilterToAlu_98, A(1)=>FilterToAlu_97, A(0)=>FilterToAlu_96, B(15)=>
      SecondInputToMult_111, B(14)=>SecondInputToMult_110, B(13)=>
      SecondInputToMult_109, B(12)=>SecondInputToMult_108, B(11)=>
      SecondInputToMult_107, B(10)=>SecondInputToMult_106, B(9)=>
      SecondInputToMult_105, B(8)=>SecondInputToMult_104, B(7)=>
      SecondInputToMult_103, B(6)=>SecondInputToMult_102, B(5)=>
      SecondInputToMult_101, B(4)=>SecondInputToMult_100, B(3)=>
      SecondInputToMult_99, B(2)=>SecondInputToMult_98, B(1)=>
      SecondInputToMult_97, B(0)=>SecondInputToMult_96, F(31)=>DANGLING(96), 
      F(30)=>DANGLING(97), F(29)=>DANGLING(98), F(28)=>DANGLING(99), F(27)=>
      DANGLING(100), F(26)=>DANGLING(101), F(25)=>DANGLING(102), F(24)=>
      MultiplierOut_216, F(23)=>MultiplierOut_215, F(22)=>MultiplierOut_214, 
      F(21)=>MultiplierOut_213, F(20)=>MultiplierOut_212, F(19)=>
      MultiplierOut_211, F(18)=>MultiplierOut_210, F(17)=>MultiplierOut_209, 
      F(16)=>MultiplierOut_208, F(15)=>MultiplierOut_207, F(14)=>
      MultiplierOut_206, F(13)=>MultiplierOut_205, F(12)=>MultiplierOut_204, 
      F(11)=>MultiplierOut_203, F(10)=>MultiplierOut_202, F(9)=>
      MultiplierOut_201, F(8)=>DANGLING(103), F(7)=>DANGLING(104), F(6)=>
      DANGLING(105), F(5)=>DANGLING(106), F(4)=>DANGLING(107), F(3)=>
      DANGLING(108), F(2)=>DANGLING(109), F(1)=>DANGLING(110), F(0)=>
      DANGLING(111));
   loop3_7_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_127, A(14)=>
      FilterToAlu_126, A(13)=>FilterToAlu_125, A(12)=>FilterToAlu_124, A(11)
      =>FilterToAlu_123, A(10)=>FilterToAlu_122, A(9)=>FilterToAlu_121, A(8)
      =>FilterToAlu_120, A(7)=>FilterToAlu_119, A(6)=>FilterToAlu_118, A(5)
      =>FilterToAlu_117, A(4)=>FilterToAlu_116, A(3)=>FilterToAlu_115, A(2)
      =>FilterToAlu_114, A(1)=>FilterToAlu_113, A(0)=>FilterToAlu_112, B(15)
      =>SecondInputToMult_127, B(14)=>SecondInputToMult_126, B(13)=>
      SecondInputToMult_125, B(12)=>SecondInputToMult_124, B(11)=>
      SecondInputToMult_123, B(10)=>SecondInputToMult_122, B(9)=>
      SecondInputToMult_121, B(8)=>SecondInputToMult_120, B(7)=>
      SecondInputToMult_119, B(6)=>SecondInputToMult_118, B(5)=>
      SecondInputToMult_117, B(4)=>SecondInputToMult_116, B(3)=>
      SecondInputToMult_115, B(2)=>SecondInputToMult_114, B(1)=>
      SecondInputToMult_113, B(0)=>SecondInputToMult_112, F(31)=>DANGLING(
      112), F(30)=>DANGLING(113), F(29)=>DANGLING(114), F(28)=>DANGLING(115), 
      F(27)=>DANGLING(116), F(26)=>DANGLING(117), F(25)=>DANGLING(118), 
      F(24)=>MultiplierOut_248, F(23)=>MultiplierOut_247, F(22)=>
      MultiplierOut_246, F(21)=>MultiplierOut_245, F(20)=>MultiplierOut_244, 
      F(19)=>MultiplierOut_243, F(18)=>MultiplierOut_242, F(17)=>
      MultiplierOut_241, F(16)=>MultiplierOut_240, F(15)=>MultiplierOut_239, 
      F(14)=>MultiplierOut_238, F(13)=>MultiplierOut_237, F(12)=>
      MultiplierOut_236, F(11)=>MultiplierOut_235, F(10)=>MultiplierOut_234, 
      F(9)=>MultiplierOut_233, F(8)=>DANGLING(119), F(7)=>DANGLING(120), 
      F(6)=>DANGLING(121), F(5)=>DANGLING(122), F(4)=>DANGLING(123), F(3)=>
      DANGLING(124), F(2)=>DANGLING(125), F(1)=>DANGLING(126), F(0)=>
      DANGLING(127));
   loop3_8_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_143, A(14)=>
      FilterToAlu_142, A(13)=>FilterToAlu_141, A(12)=>FilterToAlu_140, A(11)
      =>FilterToAlu_139, A(10)=>FilterToAlu_138, A(9)=>FilterToAlu_137, A(8)
      =>FilterToAlu_136, A(7)=>FilterToAlu_135, A(6)=>FilterToAlu_134, A(5)
      =>FilterToAlu_133, A(4)=>FilterToAlu_132, A(3)=>FilterToAlu_131, A(2)
      =>FilterToAlu_130, A(1)=>FilterToAlu_129, A(0)=>FilterToAlu_128, B(15)
      =>SecondInputToMult_143, B(14)=>SecondInputToMult_142, B(13)=>
      SecondInputToMult_141, B(12)=>SecondInputToMult_140, B(11)=>
      SecondInputToMult_139, B(10)=>SecondInputToMult_138, B(9)=>
      SecondInputToMult_137, B(8)=>SecondInputToMult_136, B(7)=>
      SecondInputToMult_135, B(6)=>SecondInputToMult_134, B(5)=>
      SecondInputToMult_133, B(4)=>SecondInputToMult_132, B(3)=>
      SecondInputToMult_131, B(2)=>SecondInputToMult_130, B(1)=>
      SecondInputToMult_129, B(0)=>SecondInputToMult_128, F(31)=>DANGLING(
      128), F(30)=>DANGLING(129), F(29)=>DANGLING(130), F(28)=>DANGLING(131), 
      F(27)=>DANGLING(132), F(26)=>DANGLING(133), F(25)=>DANGLING(134), 
      F(24)=>MultiplierOut_280, F(23)=>MultiplierOut_279, F(22)=>
      MultiplierOut_278, F(21)=>MultiplierOut_277, F(20)=>MultiplierOut_276, 
      F(19)=>MultiplierOut_275, F(18)=>MultiplierOut_274, F(17)=>
      MultiplierOut_273, F(16)=>MultiplierOut_272, F(15)=>MultiplierOut_271, 
      F(14)=>MultiplierOut_270, F(13)=>MultiplierOut_269, F(12)=>
      MultiplierOut_268, F(11)=>MultiplierOut_267, F(10)=>MultiplierOut_266, 
      F(9)=>MultiplierOut_265, F(8)=>DANGLING(135), F(7)=>DANGLING(136), 
      F(6)=>DANGLING(137), F(5)=>DANGLING(138), F(4)=>DANGLING(139), F(3)=>
      DANGLING(140), F(2)=>DANGLING(141), F(1)=>DANGLING(142), F(0)=>
      DANGLING(143));
   loop5_9_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_159, A(14)=>
      FilterToAlu_158, A(13)=>FilterToAlu_157, A(12)=>FilterToAlu_156, A(11)
      =>FilterToAlu_155, A(10)=>FilterToAlu_154, A(9)=>FilterToAlu_153, A(8)
      =>FilterToAlu_152, A(7)=>FilterToAlu_151, A(6)=>FilterToAlu_150, A(5)
      =>FilterToAlu_149, A(4)=>FilterToAlu_148, A(3)=>FilterToAlu_147, A(2)
      =>FilterToAlu_146, A(1)=>FilterToAlu_145, A(0)=>FilterToAlu_144, B(15)
      =>OutputImg1(79), B(14)=>OutputImg1(78), B(13)=>OutputImg1(77), B(12)
      =>OutputImg1(76), B(11)=>OutputImg1(75), B(10)=>OutputImg1(74), B(9)=>
      OutputImg1(73), B(8)=>OutputImg1(72), B(7)=>OutputImg1(71), B(6)=>
      OutputImg1(70), B(5)=>OutputImg1(69), B(4)=>OutputImg1(68), B(3)=>
      OutputImg1(67), B(2)=>OutputImg1(66), B(1)=>OutputImg1(65), B(0)=>
      OutputImg1(64), F(31)=>DANGLING(144), F(30)=>DANGLING(145), F(29)=>
      DANGLING(146), F(28)=>DANGLING(147), F(27)=>DANGLING(148), F(26)=>
      DANGLING(149), F(25)=>DANGLING(150), F(24)=>MultiplierOut_312, F(23)=>
      MultiplierOut_311, F(22)=>MultiplierOut_310, F(21)=>MultiplierOut_309, 
      F(20)=>MultiplierOut_308, F(19)=>MultiplierOut_307, F(18)=>
      MultiplierOut_306, F(17)=>MultiplierOut_305, F(16)=>MultiplierOut_304, 
      F(15)=>MultiplierOut_303, F(14)=>MultiplierOut_302, F(13)=>
      MultiplierOut_301, F(12)=>MultiplierOut_300, F(11)=>MultiplierOut_299, 
      F(10)=>MultiplierOut_298, F(9)=>MultiplierOut_297, F(8)=>DANGLING(151), 
      F(7)=>DANGLING(152), F(6)=>DANGLING(153), F(5)=>DANGLING(154), F(4)=>
      DANGLING(155), F(3)=>DANGLING(156), F(2)=>DANGLING(157), F(1)=>
      DANGLING(158), F(0)=>DANGLING(159));
   loop5_10_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_175, A(14)
      =>FilterToAlu_174, A(13)=>FilterToAlu_173, A(12)=>FilterToAlu_172, 
      A(11)=>FilterToAlu_171, A(10)=>FilterToAlu_170, A(9)=>FilterToAlu_169, 
      A(8)=>FilterToAlu_168, A(7)=>FilterToAlu_167, A(6)=>FilterToAlu_166, 
      A(5)=>FilterToAlu_165, A(4)=>FilterToAlu_164, A(3)=>FilterToAlu_163, 
      A(2)=>FilterToAlu_162, A(1)=>FilterToAlu_161, A(0)=>FilterToAlu_160, 
      B(15)=>OutputImg2(15), B(14)=>OutputImg2(14), B(13)=>OutputImg2(13), 
      B(12)=>OutputImg2(12), B(11)=>OutputImg2(11), B(10)=>OutputImg2(10), 
      B(9)=>OutputImg2(9), B(8)=>OutputImg2(8), B(7)=>OutputImg2(7), B(6)=>
      OutputImg2(6), B(5)=>OutputImg2(5), B(4)=>OutputImg2(4), B(3)=>
      OutputImg2(3), B(2)=>OutputImg2(2), B(1)=>OutputImg2(1), B(0)=>
      OutputImg2(0), F(31)=>DANGLING(160), F(30)=>DANGLING(161), F(29)=>
      DANGLING(162), F(28)=>DANGLING(163), F(27)=>DANGLING(164), F(26)=>
      DANGLING(165), F(25)=>DANGLING(166), F(24)=>MultiplierOut_344, F(23)=>
      MultiplierOut_343, F(22)=>MultiplierOut_342, F(21)=>MultiplierOut_341, 
      F(20)=>MultiplierOut_340, F(19)=>MultiplierOut_339, F(18)=>
      MultiplierOut_338, F(17)=>MultiplierOut_337, F(16)=>MultiplierOut_336, 
      F(15)=>MultiplierOut_335, F(14)=>MultiplierOut_334, F(13)=>
      MultiplierOut_333, F(12)=>MultiplierOut_332, F(11)=>MultiplierOut_331, 
      F(10)=>MultiplierOut_330, F(9)=>MultiplierOut_329, F(8)=>DANGLING(167), 
      F(7)=>DANGLING(168), F(6)=>DANGLING(169), F(5)=>DANGLING(170), F(4)=>
      DANGLING(171), F(3)=>DANGLING(172), F(2)=>DANGLING(173), F(1)=>
      DANGLING(174), F(0)=>DANGLING(175));
   loop5_11_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_191, A(14)
      =>FilterToAlu_190, A(13)=>FilterToAlu_189, A(12)=>FilterToAlu_188, 
      A(11)=>FilterToAlu_187, A(10)=>FilterToAlu_186, A(9)=>FilterToAlu_185, 
      A(8)=>FilterToAlu_184, A(7)=>FilterToAlu_183, A(6)=>FilterToAlu_182, 
      A(5)=>FilterToAlu_181, A(4)=>FilterToAlu_180, A(3)=>FilterToAlu_179, 
      A(2)=>FilterToAlu_178, A(1)=>FilterToAlu_177, A(0)=>FilterToAlu_176, 
      B(15)=>OutputImg2(31), B(14)=>OutputImg2(30), B(13)=>OutputImg2(29), 
      B(12)=>OutputImg2(28), B(11)=>OutputImg2(27), B(10)=>OutputImg2(26), 
      B(9)=>OutputImg2(25), B(8)=>OutputImg2(24), B(7)=>OutputImg2(23), B(6)
      =>OutputImg2(22), B(5)=>OutputImg2(21), B(4)=>OutputImg2(20), B(3)=>
      OutputImg2(19), B(2)=>OutputImg2(18), B(1)=>OutputImg2(17), B(0)=>
      OutputImg2(16), F(31)=>DANGLING(176), F(30)=>DANGLING(177), F(29)=>
      DANGLING(178), F(28)=>DANGLING(179), F(27)=>DANGLING(180), F(26)=>
      DANGLING(181), F(25)=>DANGLING(182), F(24)=>MultiplierOut_376, F(23)=>
      MultiplierOut_375, F(22)=>MultiplierOut_374, F(21)=>MultiplierOut_373, 
      F(20)=>MultiplierOut_372, F(19)=>MultiplierOut_371, F(18)=>
      MultiplierOut_370, F(17)=>MultiplierOut_369, F(16)=>MultiplierOut_368, 
      F(15)=>MultiplierOut_367, F(14)=>MultiplierOut_366, F(13)=>
      MultiplierOut_365, F(12)=>MultiplierOut_364, F(11)=>MultiplierOut_363, 
      F(10)=>MultiplierOut_362, F(9)=>MultiplierOut_361, F(8)=>DANGLING(183), 
      F(7)=>DANGLING(184), F(6)=>DANGLING(185), F(5)=>DANGLING(186), F(4)=>
      DANGLING(187), F(3)=>DANGLING(188), F(2)=>DANGLING(189), F(1)=>
      DANGLING(190), F(0)=>DANGLING(191));
   loop5_12_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_207, A(14)
      =>FilterToAlu_206, A(13)=>FilterToAlu_205, A(12)=>FilterToAlu_204, 
      A(11)=>FilterToAlu_203, A(10)=>FilterToAlu_202, A(9)=>FilterToAlu_201, 
      A(8)=>FilterToAlu_200, A(7)=>FilterToAlu_199, A(6)=>FilterToAlu_198, 
      A(5)=>FilterToAlu_197, A(4)=>FilterToAlu_196, A(3)=>FilterToAlu_195, 
      A(2)=>FilterToAlu_194, A(1)=>FilterToAlu_193, A(0)=>FilterToAlu_192, 
      B(15)=>OutputImg2(47), B(14)=>OutputImg2(46), B(13)=>OutputImg2(45), 
      B(12)=>OutputImg2(44), B(11)=>OutputImg2(43), B(10)=>OutputImg2(42), 
      B(9)=>OutputImg2(41), B(8)=>OutputImg2(40), B(7)=>OutputImg2(39), B(6)
      =>OutputImg2(38), B(5)=>OutputImg2(37), B(4)=>OutputImg2(36), B(3)=>
      OutputImg2(35), B(2)=>OutputImg2(34), B(1)=>OutputImg2(33), B(0)=>
      OutputImg2(32), F(31)=>DANGLING(192), F(30)=>DANGLING(193), F(29)=>
      DANGLING(194), F(28)=>DANGLING(195), F(27)=>DANGLING(196), F(26)=>
      DANGLING(197), F(25)=>DANGLING(198), F(24)=>MultiplierOut_408, F(23)=>
      MultiplierOut_407, F(22)=>MultiplierOut_406, F(21)=>MultiplierOut_405, 
      F(20)=>MultiplierOut_404, F(19)=>MultiplierOut_403, F(18)=>
      MultiplierOut_402, F(17)=>MultiplierOut_401, F(16)=>MultiplierOut_400, 
      F(15)=>MultiplierOut_399, F(14)=>MultiplierOut_398, F(13)=>
      MultiplierOut_397, F(12)=>MultiplierOut_396, F(11)=>MultiplierOut_395, 
      F(10)=>MultiplierOut_394, F(9)=>MultiplierOut_393, F(8)=>DANGLING(199), 
      F(7)=>DANGLING(200), F(6)=>DANGLING(201), F(5)=>DANGLING(202), F(4)=>
      DANGLING(203), F(3)=>DANGLING(204), F(2)=>DANGLING(205), F(1)=>
      DANGLING(206), F(0)=>DANGLING(207));
   loop5_13_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_223, A(14)
      =>FilterToAlu_222, A(13)=>FilterToAlu_221, A(12)=>FilterToAlu_220, 
      A(11)=>FilterToAlu_219, A(10)=>FilterToAlu_218, A(9)=>FilterToAlu_217, 
      A(8)=>FilterToAlu_216, A(7)=>FilterToAlu_215, A(6)=>FilterToAlu_214, 
      A(5)=>FilterToAlu_213, A(4)=>FilterToAlu_212, A(3)=>FilterToAlu_211, 
      A(2)=>FilterToAlu_210, A(1)=>FilterToAlu_209, A(0)=>FilterToAlu_208, 
      B(15)=>OutputImg2(63), B(14)=>OutputImg2(62), B(13)=>OutputImg2(61), 
      B(12)=>OutputImg2(60), B(11)=>OutputImg2(59), B(10)=>OutputImg2(58), 
      B(9)=>OutputImg2(57), B(8)=>OutputImg2(56), B(7)=>OutputImg2(55), B(6)
      =>OutputImg2(54), B(5)=>OutputImg2(53), B(4)=>OutputImg2(52), B(3)=>
      OutputImg2(51), B(2)=>OutputImg2(50), B(1)=>OutputImg2(49), B(0)=>
      OutputImg2(48), F(31)=>DANGLING(208), F(30)=>DANGLING(209), F(29)=>
      DANGLING(210), F(28)=>DANGLING(211), F(27)=>DANGLING(212), F(26)=>
      DANGLING(213), F(25)=>DANGLING(214), F(24)=>MultiplierOut_440, F(23)=>
      MultiplierOut_439, F(22)=>MultiplierOut_438, F(21)=>MultiplierOut_437, 
      F(20)=>MultiplierOut_436, F(19)=>MultiplierOut_435, F(18)=>
      MultiplierOut_434, F(17)=>MultiplierOut_433, F(16)=>MultiplierOut_432, 
      F(15)=>MultiplierOut_431, F(14)=>MultiplierOut_430, F(13)=>
      MultiplierOut_429, F(12)=>MultiplierOut_428, F(11)=>MultiplierOut_427, 
      F(10)=>MultiplierOut_426, F(9)=>MultiplierOut_425, F(8)=>DANGLING(215), 
      F(7)=>DANGLING(216), F(6)=>DANGLING(217), F(5)=>DANGLING(218), F(4)=>
      DANGLING(219), F(3)=>DANGLING(220), F(2)=>DANGLING(221), F(1)=>
      DANGLING(222), F(0)=>DANGLING(223));
   loop5_14_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_239, A(14)
      =>FilterToAlu_238, A(13)=>FilterToAlu_237, A(12)=>FilterToAlu_236, 
      A(11)=>FilterToAlu_235, A(10)=>FilterToAlu_234, A(9)=>FilterToAlu_233, 
      A(8)=>FilterToAlu_232, A(7)=>FilterToAlu_231, A(6)=>FilterToAlu_230, 
      A(5)=>FilterToAlu_229, A(4)=>FilterToAlu_228, A(3)=>FilterToAlu_227, 
      A(2)=>FilterToAlu_226, A(1)=>FilterToAlu_225, A(0)=>FilterToAlu_224, 
      B(15)=>OutputImg2(79), B(14)=>OutputImg2(78), B(13)=>OutputImg2(77), 
      B(12)=>OutputImg2(76), B(11)=>OutputImg2(75), B(10)=>OutputImg2(74), 
      B(9)=>OutputImg2(73), B(8)=>OutputImg2(72), B(7)=>OutputImg2(71), B(6)
      =>OutputImg2(70), B(5)=>OutputImg2(69), B(4)=>OutputImg2(68), B(3)=>
      OutputImg2(67), B(2)=>OutputImg2(66), B(1)=>OutputImg2(65), B(0)=>
      OutputImg2(64), F(31)=>DANGLING(224), F(30)=>DANGLING(225), F(29)=>
      DANGLING(226), F(28)=>DANGLING(227), F(27)=>DANGLING(228), F(26)=>
      DANGLING(229), F(25)=>DANGLING(230), F(24)=>MultiplierOut_472, F(23)=>
      MultiplierOut_471, F(22)=>MultiplierOut_470, F(21)=>MultiplierOut_469, 
      F(20)=>MultiplierOut_468, F(19)=>MultiplierOut_467, F(18)=>
      MultiplierOut_466, F(17)=>MultiplierOut_465, F(16)=>MultiplierOut_464, 
      F(15)=>MultiplierOut_463, F(14)=>MultiplierOut_462, F(13)=>
      MultiplierOut_461, F(12)=>MultiplierOut_460, F(11)=>MultiplierOut_459, 
      F(10)=>MultiplierOut_458, F(9)=>MultiplierOut_457, F(8)=>DANGLING(231), 
      F(7)=>DANGLING(232), F(6)=>DANGLING(233), F(5)=>DANGLING(234), F(4)=>
      DANGLING(235), F(3)=>DANGLING(236), F(2)=>DANGLING(237), F(1)=>
      DANGLING(238), F(0)=>DANGLING(239));
   loop5_15_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_255, A(14)
      =>FilterToAlu_254, A(13)=>FilterToAlu_253, A(12)=>FilterToAlu_252, 
      A(11)=>FilterToAlu_251, A(10)=>FilterToAlu_250, A(9)=>FilterToAlu_249, 
      A(8)=>FilterToAlu_248, A(7)=>FilterToAlu_247, A(6)=>FilterToAlu_246, 
      A(5)=>FilterToAlu_245, A(4)=>FilterToAlu_244, A(3)=>FilterToAlu_243, 
      A(2)=>FilterToAlu_242, A(1)=>FilterToAlu_241, A(0)=>FilterToAlu_240, 
      B(15)=>OutputImg3(15), B(14)=>OutputImg3(14), B(13)=>OutputImg3(13), 
      B(12)=>OutputImg3(12), B(11)=>OutputImg3(11), B(10)=>OutputImg3(10), 
      B(9)=>OutputImg3(9), B(8)=>OutputImg3(8), B(7)=>OutputImg3(7), B(6)=>
      OutputImg3(6), B(5)=>OutputImg3(5), B(4)=>OutputImg3(4), B(3)=>
      OutputImg3(3), B(2)=>OutputImg3(2), B(1)=>OutputImg3(1), B(0)=>
      OutputImg3(0), F(31)=>DANGLING(240), F(30)=>DANGLING(241), F(29)=>
      DANGLING(242), F(28)=>DANGLING(243), F(27)=>DANGLING(244), F(26)=>
      DANGLING(245), F(25)=>DANGLING(246), F(24)=>MultiplierOut_504, F(23)=>
      MultiplierOut_503, F(22)=>MultiplierOut_502, F(21)=>MultiplierOut_501, 
      F(20)=>MultiplierOut_500, F(19)=>MultiplierOut_499, F(18)=>
      MultiplierOut_498, F(17)=>MultiplierOut_497, F(16)=>MultiplierOut_496, 
      F(15)=>MultiplierOut_495, F(14)=>MultiplierOut_494, F(13)=>
      MultiplierOut_493, F(12)=>MultiplierOut_492, F(11)=>MultiplierOut_491, 
      F(10)=>MultiplierOut_490, F(9)=>MultiplierOut_489, F(8)=>DANGLING(247), 
      F(7)=>DANGLING(248), F(6)=>DANGLING(249), F(5)=>DANGLING(250), F(4)=>
      DANGLING(251), F(3)=>DANGLING(252), F(2)=>DANGLING(253), F(1)=>
      DANGLING(254), F(0)=>DANGLING(255));
   loop5_16_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_271, A(14)
      =>FilterToAlu_270, A(13)=>FilterToAlu_269, A(12)=>FilterToAlu_268, 
      A(11)=>FilterToAlu_267, A(10)=>FilterToAlu_266, A(9)=>FilterToAlu_265, 
      A(8)=>FilterToAlu_264, A(7)=>FilterToAlu_263, A(6)=>FilterToAlu_262, 
      A(5)=>FilterToAlu_261, A(4)=>FilterToAlu_260, A(3)=>FilterToAlu_259, 
      A(2)=>FilterToAlu_258, A(1)=>FilterToAlu_257, A(0)=>FilterToAlu_256, 
      B(15)=>OutputImg3(31), B(14)=>OutputImg3(30), B(13)=>OutputImg3(29), 
      B(12)=>OutputImg3(28), B(11)=>OutputImg3(27), B(10)=>OutputImg3(26), 
      B(9)=>OutputImg3(25), B(8)=>OutputImg3(24), B(7)=>OutputImg3(23), B(6)
      =>OutputImg3(22), B(5)=>OutputImg3(21), B(4)=>OutputImg3(20), B(3)=>
      OutputImg3(19), B(2)=>OutputImg3(18), B(1)=>OutputImg3(17), B(0)=>
      OutputImg3(16), F(31)=>DANGLING(256), F(30)=>DANGLING(257), F(29)=>
      DANGLING(258), F(28)=>DANGLING(259), F(27)=>DANGLING(260), F(26)=>
      DANGLING(261), F(25)=>DANGLING(262), F(24)=>MultiplierOut_536, F(23)=>
      MultiplierOut_535, F(22)=>MultiplierOut_534, F(21)=>MultiplierOut_533, 
      F(20)=>MultiplierOut_532, F(19)=>MultiplierOut_531, F(18)=>
      MultiplierOut_530, F(17)=>MultiplierOut_529, F(16)=>MultiplierOut_528, 
      F(15)=>MultiplierOut_527, F(14)=>MultiplierOut_526, F(13)=>
      MultiplierOut_525, F(12)=>MultiplierOut_524, F(11)=>MultiplierOut_523, 
      F(10)=>MultiplierOut_522, F(9)=>MultiplierOut_521, F(8)=>DANGLING(263), 
      F(7)=>DANGLING(264), F(6)=>DANGLING(265), F(5)=>DANGLING(266), F(4)=>
      DANGLING(267), F(3)=>DANGLING(268), F(2)=>DANGLING(269), F(1)=>
      DANGLING(270), F(0)=>DANGLING(271));
   loop5_17_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_287, A(14)
      =>FilterToAlu_286, A(13)=>FilterToAlu_285, A(12)=>FilterToAlu_284, 
      A(11)=>FilterToAlu_283, A(10)=>FilterToAlu_282, A(9)=>FilterToAlu_281, 
      A(8)=>FilterToAlu_280, A(7)=>FilterToAlu_279, A(6)=>FilterToAlu_278, 
      A(5)=>FilterToAlu_277, A(4)=>FilterToAlu_276, A(3)=>FilterToAlu_275, 
      A(2)=>FilterToAlu_274, A(1)=>FilterToAlu_273, A(0)=>FilterToAlu_272, 
      B(15)=>OutputImg3(47), B(14)=>OutputImg3(46), B(13)=>OutputImg3(45), 
      B(12)=>OutputImg3(44), B(11)=>OutputImg3(43), B(10)=>OutputImg3(42), 
      B(9)=>OutputImg3(41), B(8)=>OutputImg3(40), B(7)=>OutputImg3(39), B(6)
      =>OutputImg3(38), B(5)=>OutputImg3(37), B(4)=>OutputImg3(36), B(3)=>
      OutputImg3(35), B(2)=>OutputImg3(34), B(1)=>OutputImg3(33), B(0)=>
      OutputImg3(32), F(31)=>DANGLING(272), F(30)=>DANGLING(273), F(29)=>
      DANGLING(274), F(28)=>DANGLING(275), F(27)=>DANGLING(276), F(26)=>
      DANGLING(277), F(25)=>DANGLING(278), F(24)=>MultiplierOut_568, F(23)=>
      MultiplierOut_567, F(22)=>MultiplierOut_566, F(21)=>MultiplierOut_565, 
      F(20)=>MultiplierOut_564, F(19)=>MultiplierOut_563, F(18)=>
      MultiplierOut_562, F(17)=>MultiplierOut_561, F(16)=>MultiplierOut_560, 
      F(15)=>MultiplierOut_559, F(14)=>MultiplierOut_558, F(13)=>
      MultiplierOut_557, F(12)=>MultiplierOut_556, F(11)=>MultiplierOut_555, 
      F(10)=>MultiplierOut_554, F(9)=>MultiplierOut_553, F(8)=>DANGLING(279), 
      F(7)=>DANGLING(280), F(6)=>DANGLING(281), F(5)=>DANGLING(282), F(4)=>
      DANGLING(283), F(3)=>DANGLING(284), F(2)=>DANGLING(285), F(1)=>
      DANGLING(286), F(0)=>DANGLING(287));
   loop5_18_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_303, A(14)
      =>FilterToAlu_302, A(13)=>FilterToAlu_301, A(12)=>FilterToAlu_300, 
      A(11)=>FilterToAlu_299, A(10)=>FilterToAlu_298, A(9)=>FilterToAlu_297, 
      A(8)=>FilterToAlu_296, A(7)=>FilterToAlu_295, A(6)=>FilterToAlu_294, 
      A(5)=>FilterToAlu_293, A(4)=>FilterToAlu_292, A(3)=>FilterToAlu_291, 
      A(2)=>FilterToAlu_290, A(1)=>FilterToAlu_289, A(0)=>FilterToAlu_288, 
      B(15)=>OutputImg3(63), B(14)=>OutputImg3(62), B(13)=>OutputImg3(61), 
      B(12)=>OutputImg3(60), B(11)=>OutputImg3(59), B(10)=>OutputImg3(58), 
      B(9)=>OutputImg3(57), B(8)=>OutputImg3(56), B(7)=>OutputImg3(55), B(6)
      =>OutputImg3(54), B(5)=>OutputImg3(53), B(4)=>OutputImg3(52), B(3)=>
      OutputImg3(51), B(2)=>OutputImg3(50), B(1)=>OutputImg3(49), B(0)=>
      OutputImg3(48), F(31)=>DANGLING(288), F(30)=>DANGLING(289), F(29)=>
      DANGLING(290), F(28)=>DANGLING(291), F(27)=>DANGLING(292), F(26)=>
      DANGLING(293), F(25)=>DANGLING(294), F(24)=>MultiplierOut_600, F(23)=>
      MultiplierOut_599, F(22)=>MultiplierOut_598, F(21)=>MultiplierOut_597, 
      F(20)=>MultiplierOut_596, F(19)=>MultiplierOut_595, F(18)=>
      MultiplierOut_594, F(17)=>MultiplierOut_593, F(16)=>MultiplierOut_592, 
      F(15)=>MultiplierOut_591, F(14)=>MultiplierOut_590, F(13)=>
      MultiplierOut_589, F(12)=>MultiplierOut_588, F(11)=>MultiplierOut_587, 
      F(10)=>MultiplierOut_586, F(9)=>MultiplierOut_585, F(8)=>DANGLING(295), 
      F(7)=>DANGLING(296), F(6)=>DANGLING(297), F(5)=>DANGLING(298), F(4)=>
      DANGLING(299), F(3)=>DANGLING(300), F(2)=>DANGLING(301), F(1)=>
      DANGLING(302), F(0)=>DANGLING(303));
   loop5_19_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_319, A(14)
      =>FilterToAlu_318, A(13)=>FilterToAlu_317, A(12)=>FilterToAlu_316, 
      A(11)=>FilterToAlu_315, A(10)=>FilterToAlu_314, A(9)=>FilterToAlu_313, 
      A(8)=>FilterToAlu_312, A(7)=>FilterToAlu_311, A(6)=>FilterToAlu_310, 
      A(5)=>FilterToAlu_309, A(4)=>FilterToAlu_308, A(3)=>FilterToAlu_307, 
      A(2)=>FilterToAlu_306, A(1)=>FilterToAlu_305, A(0)=>FilterToAlu_304, 
      B(15)=>OutputImg3(79), B(14)=>OutputImg3(78), B(13)=>OutputImg3(77), 
      B(12)=>OutputImg3(76), B(11)=>OutputImg3(75), B(10)=>OutputImg3(74), 
      B(9)=>OutputImg3(73), B(8)=>OutputImg3(72), B(7)=>OutputImg3(71), B(6)
      =>OutputImg3(70), B(5)=>OutputImg3(69), B(4)=>OutputImg3(68), B(3)=>
      OutputImg3(67), B(2)=>OutputImg3(66), B(1)=>OutputImg3(65), B(0)=>
      OutputImg3(64), F(31)=>DANGLING(304), F(30)=>DANGLING(305), F(29)=>
      DANGLING(306), F(28)=>DANGLING(307), F(27)=>DANGLING(308), F(26)=>
      DANGLING(309), F(25)=>DANGLING(310), F(24)=>MultiplierOut_632, F(23)=>
      MultiplierOut_631, F(22)=>MultiplierOut_630, F(21)=>MultiplierOut_629, 
      F(20)=>MultiplierOut_628, F(19)=>MultiplierOut_627, F(18)=>
      MultiplierOut_626, F(17)=>MultiplierOut_625, F(16)=>MultiplierOut_624, 
      F(15)=>MultiplierOut_623, F(14)=>MultiplierOut_622, F(13)=>
      MultiplierOut_621, F(12)=>MultiplierOut_620, F(11)=>MultiplierOut_619, 
      F(10)=>MultiplierOut_618, F(9)=>MultiplierOut_617, F(8)=>DANGLING(311), 
      F(7)=>DANGLING(312), F(6)=>DANGLING(313), F(5)=>DANGLING(314), F(4)=>
      DANGLING(315), F(3)=>DANGLING(316), F(2)=>DANGLING(317), F(1)=>
      DANGLING(318), F(0)=>DANGLING(319));
   loop5_20_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_335, A(14)
      =>FilterToAlu_334, A(13)=>FilterToAlu_333, A(12)=>FilterToAlu_332, 
      A(11)=>FilterToAlu_331, A(10)=>FilterToAlu_330, A(9)=>FilterToAlu_329, 
      A(8)=>FilterToAlu_328, A(7)=>FilterToAlu_327, A(6)=>FilterToAlu_326, 
      A(5)=>FilterToAlu_325, A(4)=>FilterToAlu_324, A(3)=>FilterToAlu_323, 
      A(2)=>FilterToAlu_322, A(1)=>FilterToAlu_321, A(0)=>FilterToAlu_320, 
      B(15)=>OutputImg4(15), B(14)=>OutputImg4(14), B(13)=>OutputImg4(13), 
      B(12)=>OutputImg4(12), B(11)=>OutputImg4(11), B(10)=>OutputImg4(10), 
      B(9)=>OutputImg4(9), B(8)=>OutputImg4(8), B(7)=>OutputImg4(7), B(6)=>
      OutputImg4(6), B(5)=>OutputImg4(5), B(4)=>OutputImg4(4), B(3)=>
      OutputImg4(3), B(2)=>OutputImg4(2), B(1)=>OutputImg4(1), B(0)=>
      OutputImg4(0), F(31)=>DANGLING(320), F(30)=>DANGLING(321), F(29)=>
      DANGLING(322), F(28)=>DANGLING(323), F(27)=>DANGLING(324), F(26)=>
      DANGLING(325), F(25)=>DANGLING(326), F(24)=>MultiplierOut_664, F(23)=>
      MultiplierOut_663, F(22)=>MultiplierOut_662, F(21)=>MultiplierOut_661, 
      F(20)=>MultiplierOut_660, F(19)=>MultiplierOut_659, F(18)=>
      MultiplierOut_658, F(17)=>MultiplierOut_657, F(16)=>MultiplierOut_656, 
      F(15)=>MultiplierOut_655, F(14)=>MultiplierOut_654, F(13)=>
      MultiplierOut_653, F(12)=>MultiplierOut_652, F(11)=>MultiplierOut_651, 
      F(10)=>MultiplierOut_650, F(9)=>MultiplierOut_649, F(8)=>DANGLING(327), 
      F(7)=>DANGLING(328), F(6)=>DANGLING(329), F(5)=>DANGLING(330), F(4)=>
      DANGLING(331), F(3)=>DANGLING(332), F(2)=>DANGLING(333), F(1)=>
      DANGLING(334), F(0)=>DANGLING(335));
   loop5_21_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_351, A(14)
      =>FilterToAlu_350, A(13)=>FilterToAlu_349, A(12)=>FilterToAlu_348, 
      A(11)=>FilterToAlu_347, A(10)=>FilterToAlu_346, A(9)=>FilterToAlu_345, 
      A(8)=>FilterToAlu_344, A(7)=>FilterToAlu_343, A(6)=>FilterToAlu_342, 
      A(5)=>FilterToAlu_341, A(4)=>FilterToAlu_340, A(3)=>FilterToAlu_339, 
      A(2)=>FilterToAlu_338, A(1)=>FilterToAlu_337, A(0)=>FilterToAlu_336, 
      B(15)=>OutputImg4(31), B(14)=>OutputImg4(30), B(13)=>OutputImg4(29), 
      B(12)=>OutputImg4(28), B(11)=>OutputImg4(27), B(10)=>OutputImg4(26), 
      B(9)=>OutputImg4(25), B(8)=>OutputImg4(24), B(7)=>OutputImg4(23), B(6)
      =>OutputImg4(22), B(5)=>OutputImg4(21), B(4)=>OutputImg4(20), B(3)=>
      OutputImg4(19), B(2)=>OutputImg4(18), B(1)=>OutputImg4(17), B(0)=>
      OutputImg4(16), F(31)=>DANGLING(336), F(30)=>DANGLING(337), F(29)=>
      DANGLING(338), F(28)=>DANGLING(339), F(27)=>DANGLING(340), F(26)=>
      DANGLING(341), F(25)=>DANGLING(342), F(24)=>MultiplierOut_696, F(23)=>
      MultiplierOut_695, F(22)=>MultiplierOut_694, F(21)=>MultiplierOut_693, 
      F(20)=>MultiplierOut_692, F(19)=>MultiplierOut_691, F(18)=>
      MultiplierOut_690, F(17)=>MultiplierOut_689, F(16)=>MultiplierOut_688, 
      F(15)=>MultiplierOut_687, F(14)=>MultiplierOut_686, F(13)=>
      MultiplierOut_685, F(12)=>MultiplierOut_684, F(11)=>MultiplierOut_683, 
      F(10)=>MultiplierOut_682, F(9)=>MultiplierOut_681, F(8)=>DANGLING(343), 
      F(7)=>DANGLING(344), F(6)=>DANGLING(345), F(5)=>DANGLING(346), F(4)=>
      DANGLING(347), F(3)=>DANGLING(348), F(2)=>DANGLING(349), F(1)=>
      DANGLING(350), F(0)=>DANGLING(351));
   loop5_22_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_367, A(14)
      =>FilterToAlu_366, A(13)=>FilterToAlu_365, A(12)=>FilterToAlu_364, 
      A(11)=>FilterToAlu_363, A(10)=>FilterToAlu_362, A(9)=>FilterToAlu_361, 
      A(8)=>FilterToAlu_360, A(7)=>FilterToAlu_359, A(6)=>FilterToAlu_358, 
      A(5)=>FilterToAlu_357, A(4)=>FilterToAlu_356, A(3)=>FilterToAlu_355, 
      A(2)=>FilterToAlu_354, A(1)=>FilterToAlu_353, A(0)=>FilterToAlu_352, 
      B(15)=>OutputImg4(47), B(14)=>OutputImg4(46), B(13)=>OutputImg4(45), 
      B(12)=>OutputImg4(44), B(11)=>OutputImg4(43), B(10)=>OutputImg4(42), 
      B(9)=>OutputImg4(41), B(8)=>OutputImg4(40), B(7)=>OutputImg4(39), B(6)
      =>OutputImg4(38), B(5)=>OutputImg4(37), B(4)=>OutputImg4(36), B(3)=>
      OutputImg4(35), B(2)=>OutputImg4(34), B(1)=>OutputImg4(33), B(0)=>
      OutputImg4(32), F(31)=>DANGLING(352), F(30)=>DANGLING(353), F(29)=>
      DANGLING(354), F(28)=>DANGLING(355), F(27)=>DANGLING(356), F(26)=>
      DANGLING(357), F(25)=>DANGLING(358), F(24)=>MultiplierOut_728, F(23)=>
      MultiplierOut_727, F(22)=>MultiplierOut_726, F(21)=>MultiplierOut_725, 
      F(20)=>MultiplierOut_724, F(19)=>MultiplierOut_723, F(18)=>
      MultiplierOut_722, F(17)=>MultiplierOut_721, F(16)=>MultiplierOut_720, 
      F(15)=>MultiplierOut_719, F(14)=>MultiplierOut_718, F(13)=>
      MultiplierOut_717, F(12)=>MultiplierOut_716, F(11)=>MultiplierOut_715, 
      F(10)=>MultiplierOut_714, F(9)=>MultiplierOut_713, F(8)=>DANGLING(359), 
      F(7)=>DANGLING(360), F(6)=>DANGLING(361), F(5)=>DANGLING(362), F(4)=>
      DANGLING(363), F(3)=>DANGLING(364), F(2)=>DANGLING(365), F(1)=>
      DANGLING(366), F(0)=>DANGLING(367));
   loop5_23_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_383, A(14)
      =>FilterToAlu_382, A(13)=>FilterToAlu_381, A(12)=>FilterToAlu_380, 
      A(11)=>FilterToAlu_379, A(10)=>FilterToAlu_378, A(9)=>FilterToAlu_377, 
      A(8)=>FilterToAlu_376, A(7)=>FilterToAlu_375, A(6)=>FilterToAlu_374, 
      A(5)=>FilterToAlu_373, A(4)=>FilterToAlu_372, A(3)=>FilterToAlu_371, 
      A(2)=>FilterToAlu_370, A(1)=>FilterToAlu_369, A(0)=>FilterToAlu_368, 
      B(15)=>OutputImg4(63), B(14)=>OutputImg4(62), B(13)=>OutputImg4(61), 
      B(12)=>OutputImg4(60), B(11)=>OutputImg4(59), B(10)=>OutputImg4(58), 
      B(9)=>OutputImg4(57), B(8)=>OutputImg4(56), B(7)=>OutputImg4(55), B(6)
      =>OutputImg4(54), B(5)=>OutputImg4(53), B(4)=>OutputImg4(52), B(3)=>
      OutputImg4(51), B(2)=>OutputImg4(50), B(1)=>OutputImg4(49), B(0)=>
      OutputImg4(48), F(31)=>DANGLING(368), F(30)=>DANGLING(369), F(29)=>
      DANGLING(370), F(28)=>DANGLING(371), F(27)=>DANGLING(372), F(26)=>
      DANGLING(373), F(25)=>DANGLING(374), F(24)=>MultiplierOut_760, F(23)=>
      MultiplierOut_759, F(22)=>MultiplierOut_758, F(21)=>MultiplierOut_757, 
      F(20)=>MultiplierOut_756, F(19)=>MultiplierOut_755, F(18)=>
      MultiplierOut_754, F(17)=>MultiplierOut_753, F(16)=>MultiplierOut_752, 
      F(15)=>MultiplierOut_751, F(14)=>MultiplierOut_750, F(13)=>
      MultiplierOut_749, F(12)=>MultiplierOut_748, F(11)=>MultiplierOut_747, 
      F(10)=>MultiplierOut_746, F(9)=>MultiplierOut_745, F(8)=>DANGLING(375), 
      F(7)=>DANGLING(376), F(6)=>DANGLING(377), F(5)=>DANGLING(378), F(4)=>
      DANGLING(379), F(3)=>DANGLING(380), F(2)=>DANGLING(381), F(1)=>
      DANGLING(382), F(0)=>DANGLING(383));
   loop5_24_Multip : Multiplier_16 port map ( A(15)=>FilterToAlu_399, A(14)
      =>FilterToAlu_398, A(13)=>FilterToAlu_397, A(12)=>FilterToAlu_396, 
      A(11)=>FilterToAlu_395, A(10)=>FilterToAlu_394, A(9)=>FilterToAlu_393, 
      A(8)=>FilterToAlu_392, A(7)=>FilterToAlu_391, A(6)=>FilterToAlu_390, 
      A(5)=>FilterToAlu_389, A(4)=>FilterToAlu_388, A(3)=>FilterToAlu_387, 
      A(2)=>FilterToAlu_386, A(1)=>FilterToAlu_385, A(0)=>FilterToAlu_384, 
      B(15)=>OutputImg4(79), B(14)=>OutputImg4(78), B(13)=>OutputImg4(77), 
      B(12)=>OutputImg4(76), B(11)=>OutputImg4(75), B(10)=>OutputImg4(74), 
      B(9)=>OutputImg4(73), B(8)=>OutputImg4(72), B(7)=>OutputImg4(71), B(6)
      =>OutputImg4(70), B(5)=>OutputImg4(69), B(4)=>OutputImg4(68), B(3)=>
      OutputImg4(67), B(2)=>OutputImg4(66), B(1)=>OutputImg4(65), B(0)=>
      OutputImg4(64), F(31)=>DANGLING(384), F(30)=>DANGLING(385), F(29)=>
      DANGLING(386), F(28)=>DANGLING(387), F(27)=>DANGLING(388), F(26)=>
      DANGLING(389), F(25)=>DANGLING(390), F(24)=>MultiplierOut_792, F(23)=>
      MultiplierOut_791, F(22)=>MultiplierOut_790, F(21)=>MultiplierOut_789, 
      F(20)=>MultiplierOut_788, F(19)=>MultiplierOut_787, F(18)=>
      MultiplierOut_786, F(17)=>MultiplierOut_785, F(16)=>MultiplierOut_784, 
      F(15)=>MultiplierOut_783, F(14)=>MultiplierOut_782, F(13)=>
      MultiplierOut_781, F(12)=>MultiplierOut_780, F(11)=>MultiplierOut_779, 
      F(10)=>MultiplierOut_778, F(9)=>MultiplierOut_777, F(8)=>DANGLING(391), 
      F(7)=>DANGLING(392), F(6)=>DANGLING(393), F(5)=>DANGLING(394), F(4)=>
      DANGLING(395), F(3)=>DANGLING(396), F(2)=>DANGLING(397), F(1)=>
      DANGLING(398), F(0)=>DANGLING(399));
   adder1 : my_nadder_16 port map ( a(15)=>MultiplierOut_24, a(14)=>
      MultiplierOut_23, a(13)=>MultiplierOut_22, a(12)=>MultiplierOut_21, 
      a(11)=>MultiplierOut_20, a(10)=>MultiplierOut_19, a(9)=>
      MultiplierOut_18, a(8)=>MultiplierOut_17, a(7)=>MultiplierOut_16, a(6)
      =>MultiplierOut_15, a(5)=>MultiplierOut_14, a(4)=>MultiplierOut_13, 
      a(3)=>MultiplierOut_12, a(2)=>MultiplierOut_11, a(1)=>MultiplierOut_10, 
      a(0)=>MultiplierOut_9, b(15)=>MultiplierOut_56, b(14)=>
      MultiplierOut_55, b(13)=>MultiplierOut_54, b(12)=>MultiplierOut_53, 
      b(11)=>MultiplierOut_52, b(10)=>MultiplierOut_51, b(9)=>
      MultiplierOut_50, b(8)=>MultiplierOut_49, b(7)=>MultiplierOut_48, b(6)
      =>MultiplierOut_47, b(5)=>MultiplierOut_46, b(4)=>MultiplierOut_45, 
      b(3)=>MultiplierOut_44, b(2)=>MultiplierOut_43, b(1)=>MultiplierOut_42, 
      b(0)=>MultiplierOut_41, cin=>GND0, s(15)=>AddOutputLvL1_15, s(14)=>
      AddOutputLvL1_14, s(13)=>AddOutputLvL1_13, s(12)=>AddOutputLvL1_12, 
      s(11)=>AddOutputLvL1_11, s(10)=>AddOutputLvL1_10, s(9)=>
      AddOutputLvL1_9, s(8)=>AddOutputLvL1_8, s(7)=>AddOutputLvL1_7, s(6)=>
      AddOutputLvL1_6, s(5)=>AddOutputLvL1_5, s(4)=>AddOutputLvL1_4, s(3)=>
      AddOutputLvL1_3, s(2)=>AddOutputLvL1_2, s(1)=>AddOutputLvL1_1, s(0)=>
      AddOutputLvL1_0, cout=>DANGLING(400));
   adder2 : my_nadder_16 port map ( a(15)=>MultiplierOut_88, a(14)=>
      MultiplierOut_87, a(13)=>MultiplierOut_86, a(12)=>MultiplierOut_85, 
      a(11)=>MultiplierOut_84, a(10)=>MultiplierOut_83, a(9)=>
      MultiplierOut_82, a(8)=>MultiplierOut_81, a(7)=>MultiplierOut_80, a(6)
      =>MultiplierOut_79, a(5)=>MultiplierOut_78, a(4)=>MultiplierOut_77, 
      a(3)=>MultiplierOut_76, a(2)=>MultiplierOut_75, a(1)=>MultiplierOut_74, 
      a(0)=>MultiplierOut_73, b(15)=>MultiplierOut_120, b(14)=>
      MultiplierOut_119, b(13)=>MultiplierOut_118, b(12)=>MultiplierOut_117, 
      b(11)=>MultiplierOut_116, b(10)=>MultiplierOut_115, b(9)=>
      MultiplierOut_114, b(8)=>MultiplierOut_113, b(7)=>MultiplierOut_112, 
      b(6)=>MultiplierOut_111, b(5)=>MultiplierOut_110, b(4)=>
      MultiplierOut_109, b(3)=>MultiplierOut_108, b(2)=>MultiplierOut_107, 
      b(1)=>MultiplierOut_106, b(0)=>MultiplierOut_105, cin=>GND0, s(15)=>
      AddOutputLvL1_31, s(14)=>AddOutputLvL1_30, s(13)=>AddOutputLvL1_29, 
      s(12)=>AddOutputLvL1_28, s(11)=>AddOutputLvL1_27, s(10)=>
      AddOutputLvL1_26, s(9)=>AddOutputLvL1_25, s(8)=>AddOutputLvL1_24, s(7)
      =>AddOutputLvL1_23, s(6)=>AddOutputLvL1_22, s(5)=>AddOutputLvL1_21, 
      s(4)=>AddOutputLvL1_20, s(3)=>AddOutputLvL1_19, s(2)=>AddOutputLvL1_18, 
      s(1)=>AddOutputLvL1_17, s(0)=>AddOutputLvL1_16, cout=>DANGLING(401));
   adder3 : my_nadder_16 port map ( a(15)=>MultiplierOut_152, a(14)=>
      MultiplierOut_151, a(13)=>MultiplierOut_150, a(12)=>MultiplierOut_149, 
      a(11)=>MultiplierOut_148, a(10)=>MultiplierOut_147, a(9)=>
      MultiplierOut_146, a(8)=>MultiplierOut_145, a(7)=>MultiplierOut_144, 
      a(6)=>MultiplierOut_143, a(5)=>MultiplierOut_142, a(4)=>
      MultiplierOut_141, a(3)=>MultiplierOut_140, a(2)=>MultiplierOut_139, 
      a(1)=>MultiplierOut_138, a(0)=>MultiplierOut_137, b(15)=>
      MultiplierOut_184, b(14)=>MultiplierOut_183, b(13)=>MultiplierOut_182, 
      b(12)=>MultiplierOut_181, b(11)=>MultiplierOut_180, b(10)=>
      MultiplierOut_179, b(9)=>MultiplierOut_178, b(8)=>MultiplierOut_177, 
      b(7)=>MultiplierOut_176, b(6)=>MultiplierOut_175, b(5)=>
      MultiplierOut_174, b(4)=>MultiplierOut_173, b(3)=>MultiplierOut_172, 
      b(2)=>MultiplierOut_171, b(1)=>MultiplierOut_170, b(0)=>
      MultiplierOut_169, cin=>GND0, s(15)=>AddOutputLvL1_47, s(14)=>
      AddOutputLvL1_46, s(13)=>AddOutputLvL1_45, s(12)=>AddOutputLvL1_44, 
      s(11)=>AddOutputLvL1_43, s(10)=>AddOutputLvL1_42, s(9)=>
      AddOutputLvL1_41, s(8)=>AddOutputLvL1_40, s(7)=>AddOutputLvL1_39, s(6)
      =>AddOutputLvL1_38, s(5)=>AddOutputLvL1_37, s(4)=>AddOutputLvL1_36, 
      s(3)=>AddOutputLvL1_35, s(2)=>AddOutputLvL1_34, s(1)=>AddOutputLvL1_33, 
      s(0)=>AddOutputLvL1_32, cout=>DANGLING(402));
   adder4 : my_nadder_16 port map ( a(15)=>MultiplierOut_216, a(14)=>
      MultiplierOut_215, a(13)=>MultiplierOut_214, a(12)=>MultiplierOut_213, 
      a(11)=>MultiplierOut_212, a(10)=>MultiplierOut_211, a(9)=>
      MultiplierOut_210, a(8)=>MultiplierOut_209, a(7)=>MultiplierOut_208, 
      a(6)=>MultiplierOut_207, a(5)=>MultiplierOut_206, a(4)=>
      MultiplierOut_205, a(3)=>MultiplierOut_204, a(2)=>MultiplierOut_203, 
      a(1)=>MultiplierOut_202, a(0)=>MultiplierOut_201, b(15)=>
      MultiplierOut_248, b(14)=>MultiplierOut_247, b(13)=>MultiplierOut_246, 
      b(12)=>MultiplierOut_245, b(11)=>MultiplierOut_244, b(10)=>
      MultiplierOut_243, b(9)=>MultiplierOut_242, b(8)=>MultiplierOut_241, 
      b(7)=>MultiplierOut_240, b(6)=>MultiplierOut_239, b(5)=>
      MultiplierOut_238, b(4)=>MultiplierOut_237, b(3)=>MultiplierOut_236, 
      b(2)=>MultiplierOut_235, b(1)=>MultiplierOut_234, b(0)=>
      MultiplierOut_233, cin=>GND0, s(15)=>AddOutputLvL1_63, s(14)=>
      AddOutputLvL1_62, s(13)=>AddOutputLvL1_61, s(12)=>AddOutputLvL1_60, 
      s(11)=>AddOutputLvL1_59, s(10)=>AddOutputLvL1_58, s(9)=>
      AddOutputLvL1_57, s(8)=>AddOutputLvL1_56, s(7)=>AddOutputLvL1_55, s(6)
      =>AddOutputLvL1_54, s(5)=>AddOutputLvL1_53, s(4)=>AddOutputLvL1_52, 
      s(3)=>AddOutputLvL1_51, s(2)=>AddOutputLvL1_50, s(1)=>AddOutputLvL1_49, 
      s(0)=>AddOutputLvL1_48, cout=>DANGLING(403));
   adder12 : my_nadder_16 port map ( a(15)=>AddOutputLvL1_15, a(14)=>
      AddOutputLvL1_14, a(13)=>AddOutputLvL1_13, a(12)=>AddOutputLvL1_12, 
      a(11)=>AddOutputLvL1_11, a(10)=>AddOutputLvL1_10, a(9)=>
      AddOutputLvL1_9, a(8)=>AddOutputLvL1_8, a(7)=>AddOutputLvL1_7, a(6)=>
      AddOutputLvL1_6, a(5)=>AddOutputLvL1_5, a(4)=>AddOutputLvL1_4, a(3)=>
      AddOutputLvL1_3, a(2)=>AddOutputLvL1_2, a(1)=>AddOutputLvL1_1, a(0)=>
      AddOutputLvL1_0, b(15)=>AddOutputLvL1_31, b(14)=>AddOutputLvL1_30, 
      b(13)=>AddOutputLvL1_29, b(12)=>AddOutputLvL1_28, b(11)=>
      AddOutputLvL1_27, b(10)=>AddOutputLvL1_26, b(9)=>AddOutputLvL1_25, 
      b(8)=>AddOutputLvL1_24, b(7)=>AddOutputLvL1_23, b(6)=>AddOutputLvL1_22, 
      b(5)=>AddOutputLvL1_21, b(4)=>AddOutputLvL1_20, b(3)=>AddOutputLvL1_19, 
      b(2)=>AddOutputLvL1_18, b(1)=>AddOutputLvL1_17, b(0)=>AddOutputLvL1_16, 
      cin=>GND0, s(15)=>AddOutputLvL2_15, s(14)=>AddOutputLvL2_14, s(13)=>
      AddOutputLvL2_13, s(12)=>AddOutputLvL2_12, s(11)=>AddOutputLvL2_11, 
      s(10)=>AddOutputLvL2_10, s(9)=>AddOutputLvL2_9, s(8)=>AddOutputLvL2_8, 
      s(7)=>AddOutputLvL2_7, s(6)=>AddOutputLvL2_6, s(5)=>AddOutputLvL2_5, 
      s(4)=>AddOutputLvL2_4, s(3)=>AddOutputLvL2_3, s(2)=>AddOutputLvL2_2, 
      s(1)=>AddOutputLvL2_1, s(0)=>AddOutputLvL2_0, cout=>DANGLING(404));
   adder13 : my_nadder_16 port map ( a(15)=>AddOutputLvL1_47, a(14)=>
      AddOutputLvL1_46, a(13)=>AddOutputLvL1_45, a(12)=>AddOutputLvL1_44, 
      a(11)=>AddOutputLvL1_43, a(10)=>AddOutputLvL1_42, a(9)=>
      AddOutputLvL1_41, a(8)=>AddOutputLvL1_40, a(7)=>AddOutputLvL1_39, a(6)
      =>AddOutputLvL1_38, a(5)=>AddOutputLvL1_37, a(4)=>AddOutputLvL1_36, 
      a(3)=>AddOutputLvL1_35, a(2)=>AddOutputLvL1_34, a(1)=>AddOutputLvL1_33, 
      a(0)=>AddOutputLvL1_32, b(15)=>AddOutputLvL1_63, b(14)=>
      AddOutputLvL1_62, b(13)=>AddOutputLvL1_61, b(12)=>AddOutputLvL1_60, 
      b(11)=>AddOutputLvL1_59, b(10)=>AddOutputLvL1_58, b(9)=>
      AddOutputLvL1_57, b(8)=>AddOutputLvL1_56, b(7)=>AddOutputLvL1_55, b(6)
      =>AddOutputLvL1_54, b(5)=>AddOutputLvL1_53, b(4)=>AddOutputLvL1_52, 
      b(3)=>AddOutputLvL1_51, b(2)=>AddOutputLvL1_50, b(1)=>AddOutputLvL1_49, 
      b(0)=>AddOutputLvL1_48, cin=>GND0, s(15)=>AddOutputLvL2_31, s(14)=>
      AddOutputLvL2_30, s(13)=>AddOutputLvL2_29, s(12)=>AddOutputLvL2_28, 
      s(11)=>AddOutputLvL2_27, s(10)=>AddOutputLvL2_26, s(9)=>
      AddOutputLvL2_25, s(8)=>AddOutputLvL2_24, s(7)=>AddOutputLvL2_23, s(6)
      =>AddOutputLvL2_22, s(5)=>AddOutputLvL2_21, s(4)=>AddOutputLvL2_20, 
      s(3)=>AddOutputLvL2_19, s(2)=>AddOutputLvL2_18, s(1)=>AddOutputLvL2_17, 
      s(0)=>AddOutputLvL2_16, cout=>DANGLING(405));
   adder18 : my_nadder_16 port map ( a(15)=>AddOutputLvL2_15, a(14)=>
      AddOutputLvL2_14, a(13)=>AddOutputLvL2_13, a(12)=>AddOutputLvL2_12, 
      a(11)=>AddOutputLvL2_11, a(10)=>AddOutputLvL2_10, a(9)=>
      AddOutputLvL2_9, a(8)=>AddOutputLvL2_8, a(7)=>AddOutputLvL2_7, a(6)=>
      AddOutputLvL2_6, a(5)=>AddOutputLvL2_5, a(4)=>AddOutputLvL2_4, a(3)=>
      AddOutputLvL2_3, a(2)=>AddOutputLvL2_2, a(1)=>AddOutputLvL2_1, a(0)=>
      AddOutputLvL2_0, b(15)=>AddOutputLvL2_31, b(14)=>AddOutputLvL2_30, 
      b(13)=>AddOutputLvL2_29, b(12)=>AddOutputLvL2_28, b(11)=>
      AddOutputLvL2_27, b(10)=>AddOutputLvL2_26, b(9)=>AddOutputLvL2_25, 
      b(8)=>AddOutputLvL2_24, b(7)=>AddOutputLvL2_23, b(6)=>AddOutputLvL2_22, 
      b(5)=>AddOutputLvL2_21, b(4)=>AddOutputLvL2_20, b(3)=>AddOutputLvL2_19, 
      b(2)=>AddOutputLvL2_18, b(1)=>AddOutputLvL2_17, b(0)=>AddOutputLvL2_16, 
      cin=>GND0, s(15)=>AddOutputLvL3_15, s(14)=>AddOutputLvL3_14, s(13)=>
      AddOutputLvL3_13, s(12)=>AddOutputLvL3_12, s(11)=>AddOutputLvL3_11, 
      s(10)=>AddOutputLvL3_10, s(9)=>AddOutputLvL3_9, s(8)=>AddOutputLvL3_8, 
      s(7)=>AddOutputLvL3_7, s(6)=>AddOutputLvL3_6, s(5)=>AddOutputLvL3_5, 
      s(4)=>AddOutputLvL3_4, s(3)=>AddOutputLvL3_3, s(2)=>AddOutputLvL3_2, 
      s(1)=>AddOutputLvL3_1, s(0)=>AddOutputLvL3_0, cout=>DANGLING(406));
   adder21 : my_nadder_16 port map ( a(15)=>AddOutputLvL3_15, a(14)=>
      AddOutputLvL3_14, a(13)=>AddOutputLvL3_13, a(12)=>AddOutputLvL3_12, 
      a(11)=>AddOutputLvL3_11, a(10)=>AddOutputLvL3_10, a(9)=>
      AddOutputLvL3_9, a(8)=>AddOutputLvL3_8, a(7)=>AddOutputLvL3_7, a(6)=>
      AddOutputLvL3_6, a(5)=>AddOutputLvL3_5, a(4)=>AddOutputLvL3_4, a(3)=>
      AddOutputLvL3_3, a(2)=>AddOutputLvL3_2, a(1)=>AddOutputLvL3_1, a(0)=>
      AddOutputLvL3_0, b(15)=>MultiplierOut_280, b(14)=>MultiplierOut_279, 
      b(13)=>MultiplierOut_278, b(12)=>MultiplierOut_277, b(11)=>
      MultiplierOut_276, b(10)=>MultiplierOut_275, b(9)=>MultiplierOut_274, 
      b(8)=>MultiplierOut_273, b(7)=>MultiplierOut_272, b(6)=>
      MultiplierOut_271, b(5)=>MultiplierOut_270, b(4)=>MultiplierOut_269, 
      b(3)=>MultiplierOut_268, b(2)=>MultiplierOut_267, b(1)=>
      MultiplierOut_266, b(0)=>MultiplierOut_265, cin=>GND0, s(15)=>
      AddOut33_15, s(14)=>AddOut33_14, s(13)=>AddOut33_13, s(12)=>
      AddOut33_12, s(11)=>AddOut33_11, s(10)=>AddOut33_10, s(9)=>AddOut33_9, 
      s(8)=>AddOut33_8, s(7)=>AddOut33_7, s(6)=>AddOut33_6, s(5)=>AddOut33_5, 
      s(4)=>AddOut33_4, s(3)=>AddOut33_3, s(2)=>AddOut33_2, s(1)=>AddOut33_1, 
      s(0)=>AddOut33_0, cout=>DANGLING(407));
   adder5 : my_nadder_16 port map ( a(15)=>MultiplierOut_312, a(14)=>
      MultiplierOut_311, a(13)=>MultiplierOut_310, a(12)=>MultiplierOut_309, 
      a(11)=>MultiplierOut_308, a(10)=>MultiplierOut_307, a(9)=>
      MultiplierOut_306, a(8)=>MultiplierOut_305, a(7)=>MultiplierOut_304, 
      a(6)=>MultiplierOut_303, a(5)=>MultiplierOut_302, a(4)=>
      MultiplierOut_301, a(3)=>MultiplierOut_300, a(2)=>MultiplierOut_299, 
      a(1)=>MultiplierOut_298, a(0)=>MultiplierOut_297, b(15)=>
      MultiplierOut_344, b(14)=>MultiplierOut_343, b(13)=>MultiplierOut_342, 
      b(12)=>MultiplierOut_341, b(11)=>MultiplierOut_340, b(10)=>
      MultiplierOut_339, b(9)=>MultiplierOut_338, b(8)=>MultiplierOut_337, 
      b(7)=>MultiplierOut_336, b(6)=>MultiplierOut_335, b(5)=>
      MultiplierOut_334, b(4)=>MultiplierOut_333, b(3)=>MultiplierOut_332, 
      b(2)=>MultiplierOut_331, b(1)=>MultiplierOut_330, b(0)=>
      MultiplierOut_329, cin=>GND0, s(15)=>AddOutputLvL1_79, s(14)=>
      AddOutputLvL1_78, s(13)=>AddOutputLvL1_77, s(12)=>AddOutputLvL1_76, 
      s(11)=>AddOutputLvL1_75, s(10)=>AddOutputLvL1_74, s(9)=>
      AddOutputLvL1_73, s(8)=>AddOutputLvL1_72, s(7)=>AddOutputLvL1_71, s(6)
      =>AddOutputLvL1_70, s(5)=>AddOutputLvL1_69, s(4)=>AddOutputLvL1_68, 
      s(3)=>AddOutputLvL1_67, s(2)=>AddOutputLvL1_66, s(1)=>AddOutputLvL1_65, 
      s(0)=>AddOutputLvL1_64, cout=>DANGLING(408));
   adder6 : my_nadder_16 port map ( a(15)=>MultiplierOut_376, a(14)=>
      MultiplierOut_375, a(13)=>MultiplierOut_374, a(12)=>MultiplierOut_373, 
      a(11)=>MultiplierOut_372, a(10)=>MultiplierOut_371, a(9)=>
      MultiplierOut_370, a(8)=>MultiplierOut_369, a(7)=>MultiplierOut_368, 
      a(6)=>MultiplierOut_367, a(5)=>MultiplierOut_366, a(4)=>
      MultiplierOut_365, a(3)=>MultiplierOut_364, a(2)=>MultiplierOut_363, 
      a(1)=>MultiplierOut_362, a(0)=>MultiplierOut_361, b(15)=>
      MultiplierOut_408, b(14)=>MultiplierOut_407, b(13)=>MultiplierOut_406, 
      b(12)=>MultiplierOut_405, b(11)=>MultiplierOut_404, b(10)=>
      MultiplierOut_403, b(9)=>MultiplierOut_402, b(8)=>MultiplierOut_401, 
      b(7)=>MultiplierOut_400, b(6)=>MultiplierOut_399, b(5)=>
      MultiplierOut_398, b(4)=>MultiplierOut_397, b(3)=>MultiplierOut_396, 
      b(2)=>MultiplierOut_395, b(1)=>MultiplierOut_394, b(0)=>
      MultiplierOut_393, cin=>GND0, s(15)=>AddOutputLvL1_95, s(14)=>
      AddOutputLvL1_94, s(13)=>AddOutputLvL1_93, s(12)=>AddOutputLvL1_92, 
      s(11)=>AddOutputLvL1_91, s(10)=>AddOutputLvL1_90, s(9)=>
      AddOutputLvL1_89, s(8)=>AddOutputLvL1_88, s(7)=>AddOutputLvL1_87, s(6)
      =>AddOutputLvL1_86, s(5)=>AddOutputLvL1_85, s(4)=>AddOutputLvL1_84, 
      s(3)=>AddOutputLvL1_83, s(2)=>AddOutputLvL1_82, s(1)=>AddOutputLvL1_81, 
      s(0)=>AddOutputLvL1_80, cout=>DANGLING(409));
   adder7 : my_nadder_16 port map ( a(15)=>MultiplierOut_440, a(14)=>
      MultiplierOut_439, a(13)=>MultiplierOut_438, a(12)=>MultiplierOut_437, 
      a(11)=>MultiplierOut_436, a(10)=>MultiplierOut_435, a(9)=>
      MultiplierOut_434, a(8)=>MultiplierOut_433, a(7)=>MultiplierOut_432, 
      a(6)=>MultiplierOut_431, a(5)=>MultiplierOut_430, a(4)=>
      MultiplierOut_429, a(3)=>MultiplierOut_428, a(2)=>MultiplierOut_427, 
      a(1)=>MultiplierOut_426, a(0)=>MultiplierOut_425, b(15)=>
      MultiplierOut_472, b(14)=>MultiplierOut_471, b(13)=>MultiplierOut_470, 
      b(12)=>MultiplierOut_469, b(11)=>MultiplierOut_468, b(10)=>
      MultiplierOut_467, b(9)=>MultiplierOut_466, b(8)=>MultiplierOut_465, 
      b(7)=>MultiplierOut_464, b(6)=>MultiplierOut_463, b(5)=>
      MultiplierOut_462, b(4)=>MultiplierOut_461, b(3)=>MultiplierOut_460, 
      b(2)=>MultiplierOut_459, b(1)=>MultiplierOut_458, b(0)=>
      MultiplierOut_457, cin=>GND0, s(15)=>AddOutputLvL1_111, s(14)=>
      AddOutputLvL1_110, s(13)=>AddOutputLvL1_109, s(12)=>AddOutputLvL1_108, 
      s(11)=>AddOutputLvL1_107, s(10)=>AddOutputLvL1_106, s(9)=>
      AddOutputLvL1_105, s(8)=>AddOutputLvL1_104, s(7)=>AddOutputLvL1_103, 
      s(6)=>AddOutputLvL1_102, s(5)=>AddOutputLvL1_101, s(4)=>
      AddOutputLvL1_100, s(3)=>AddOutputLvL1_99, s(2)=>AddOutputLvL1_98, 
      s(1)=>AddOutputLvL1_97, s(0)=>AddOutputLvL1_96, cout=>DANGLING(410));
   adder8 : my_nadder_16 port map ( a(15)=>MultiplierOut_504, a(14)=>
      MultiplierOut_503, a(13)=>MultiplierOut_502, a(12)=>MultiplierOut_501, 
      a(11)=>MultiplierOut_500, a(10)=>MultiplierOut_499, a(9)=>
      MultiplierOut_498, a(8)=>MultiplierOut_497, a(7)=>MultiplierOut_496, 
      a(6)=>MultiplierOut_495, a(5)=>MultiplierOut_494, a(4)=>
      MultiplierOut_493, a(3)=>MultiplierOut_492, a(2)=>MultiplierOut_491, 
      a(1)=>MultiplierOut_490, a(0)=>MultiplierOut_489, b(15)=>
      MultiplierOut_536, b(14)=>MultiplierOut_535, b(13)=>MultiplierOut_534, 
      b(12)=>MultiplierOut_533, b(11)=>MultiplierOut_532, b(10)=>
      MultiplierOut_531, b(9)=>MultiplierOut_530, b(8)=>MultiplierOut_529, 
      b(7)=>MultiplierOut_528, b(6)=>MultiplierOut_527, b(5)=>
      MultiplierOut_526, b(4)=>MultiplierOut_525, b(3)=>MultiplierOut_524, 
      b(2)=>MultiplierOut_523, b(1)=>MultiplierOut_522, b(0)=>
      MultiplierOut_521, cin=>GND0, s(15)=>AddOutputLvL1_127, s(14)=>
      AddOutputLvL1_126, s(13)=>AddOutputLvL1_125, s(12)=>AddOutputLvL1_124, 
      s(11)=>AddOutputLvL1_123, s(10)=>AddOutputLvL1_122, s(9)=>
      AddOutputLvL1_121, s(8)=>AddOutputLvL1_120, s(7)=>AddOutputLvL1_119, 
      s(6)=>AddOutputLvL1_118, s(5)=>AddOutputLvL1_117, s(4)=>
      AddOutputLvL1_116, s(3)=>AddOutputLvL1_115, s(2)=>AddOutputLvL1_114, 
      s(1)=>AddOutputLvL1_113, s(0)=>AddOutputLvL1_112, cout=>DANGLING(411)
   );
   adder9 : my_nadder_16 port map ( a(15)=>MultiplierOut_568, a(14)=>
      MultiplierOut_567, a(13)=>MultiplierOut_566, a(12)=>MultiplierOut_565, 
      a(11)=>MultiplierOut_564, a(10)=>MultiplierOut_563, a(9)=>
      MultiplierOut_562, a(8)=>MultiplierOut_561, a(7)=>MultiplierOut_560, 
      a(6)=>MultiplierOut_559, a(5)=>MultiplierOut_558, a(4)=>
      MultiplierOut_557, a(3)=>MultiplierOut_556, a(2)=>MultiplierOut_555, 
      a(1)=>MultiplierOut_554, a(0)=>MultiplierOut_553, b(15)=>
      MultiplierOut_600, b(14)=>MultiplierOut_599, b(13)=>MultiplierOut_598, 
      b(12)=>MultiplierOut_597, b(11)=>MultiplierOut_596, b(10)=>
      MultiplierOut_595, b(9)=>MultiplierOut_594, b(8)=>MultiplierOut_593, 
      b(7)=>MultiplierOut_592, b(6)=>MultiplierOut_591, b(5)=>
      MultiplierOut_590, b(4)=>MultiplierOut_589, b(3)=>MultiplierOut_588, 
      b(2)=>MultiplierOut_587, b(1)=>MultiplierOut_586, b(0)=>
      MultiplierOut_585, cin=>GND0, s(15)=>AddOutputLvL1_143, s(14)=>
      AddOutputLvL1_142, s(13)=>AddOutputLvL1_141, s(12)=>AddOutputLvL1_140, 
      s(11)=>AddOutputLvL1_139, s(10)=>AddOutputLvL1_138, s(9)=>
      AddOutputLvL1_137, s(8)=>AddOutputLvL1_136, s(7)=>AddOutputLvL1_135, 
      s(6)=>AddOutputLvL1_134, s(5)=>AddOutputLvL1_133, s(4)=>
      AddOutputLvL1_132, s(3)=>AddOutputLvL1_131, s(2)=>AddOutputLvL1_130, 
      s(1)=>AddOutputLvL1_129, s(0)=>AddOutputLvL1_128, cout=>DANGLING(412)
   );
   adder10 : my_nadder_16 port map ( a(15)=>MultiplierOut_632, a(14)=>
      MultiplierOut_631, a(13)=>MultiplierOut_630, a(12)=>MultiplierOut_629, 
      a(11)=>MultiplierOut_628, a(10)=>MultiplierOut_627, a(9)=>
      MultiplierOut_626, a(8)=>MultiplierOut_625, a(7)=>MultiplierOut_624, 
      a(6)=>MultiplierOut_623, a(5)=>MultiplierOut_622, a(4)=>
      MultiplierOut_621, a(3)=>MultiplierOut_620, a(2)=>MultiplierOut_619, 
      a(1)=>MultiplierOut_618, a(0)=>MultiplierOut_617, b(15)=>
      MultiplierOut_664, b(14)=>MultiplierOut_663, b(13)=>MultiplierOut_662, 
      b(12)=>MultiplierOut_661, b(11)=>MultiplierOut_660, b(10)=>
      MultiplierOut_659, b(9)=>MultiplierOut_658, b(8)=>MultiplierOut_657, 
      b(7)=>MultiplierOut_656, b(6)=>MultiplierOut_655, b(5)=>
      MultiplierOut_654, b(4)=>MultiplierOut_653, b(3)=>MultiplierOut_652, 
      b(2)=>MultiplierOut_651, b(1)=>MultiplierOut_650, b(0)=>
      MultiplierOut_649, cin=>GND0, s(15)=>AddOutputLvL1_159, s(14)=>
      AddOutputLvL1_158, s(13)=>AddOutputLvL1_157, s(12)=>AddOutputLvL1_156, 
      s(11)=>AddOutputLvL1_155, s(10)=>AddOutputLvL1_154, s(9)=>
      AddOutputLvL1_153, s(8)=>AddOutputLvL1_152, s(7)=>AddOutputLvL1_151, 
      s(6)=>AddOutputLvL1_150, s(5)=>AddOutputLvL1_149, s(4)=>
      AddOutputLvL1_148, s(3)=>AddOutputLvL1_147, s(2)=>AddOutputLvL1_146, 
      s(1)=>AddOutputLvL1_145, s(0)=>AddOutputLvL1_144, cout=>DANGLING(413)
   );
   adder11 : my_nadder_16 port map ( a(15)=>MultiplierOut_696, a(14)=>
      MultiplierOut_695, a(13)=>MultiplierOut_694, a(12)=>MultiplierOut_693, 
      a(11)=>MultiplierOut_692, a(10)=>MultiplierOut_691, a(9)=>
      MultiplierOut_690, a(8)=>MultiplierOut_689, a(7)=>MultiplierOut_688, 
      a(6)=>MultiplierOut_687, a(5)=>MultiplierOut_686, a(4)=>
      MultiplierOut_685, a(3)=>MultiplierOut_684, a(2)=>MultiplierOut_683, 
      a(1)=>MultiplierOut_682, a(0)=>MultiplierOut_681, b(15)=>
      MultiplierOut_728, b(14)=>MultiplierOut_727, b(13)=>MultiplierOut_726, 
      b(12)=>MultiplierOut_725, b(11)=>MultiplierOut_724, b(10)=>
      MultiplierOut_723, b(9)=>MultiplierOut_722, b(8)=>MultiplierOut_721, 
      b(7)=>MultiplierOut_720, b(6)=>MultiplierOut_719, b(5)=>
      MultiplierOut_718, b(4)=>MultiplierOut_717, b(3)=>MultiplierOut_716, 
      b(2)=>MultiplierOut_715, b(1)=>MultiplierOut_714, b(0)=>
      MultiplierOut_713, cin=>GND0, s(15)=>AddOutputLvL1_175, s(14)=>
      AddOutputLvL1_174, s(13)=>AddOutputLvL1_173, s(12)=>AddOutputLvL1_172, 
      s(11)=>AddOutputLvL1_171, s(10)=>AddOutputLvL1_170, s(9)=>
      AddOutputLvL1_169, s(8)=>AddOutputLvL1_168, s(7)=>AddOutputLvL1_167, 
      s(6)=>AddOutputLvL1_166, s(5)=>AddOutputLvL1_165, s(4)=>
      AddOutputLvL1_164, s(3)=>AddOutputLvL1_163, s(2)=>AddOutputLvL1_162, 
      s(1)=>AddOutputLvL1_161, s(0)=>AddOutputLvL1_160, cout=>DANGLING(414)
   );
   adder0 : my_nadder_16 port map ( a(15)=>MultiplierOut_760, a(14)=>
      MultiplierOut_759, a(13)=>MultiplierOut_758, a(12)=>MultiplierOut_757, 
      a(11)=>MultiplierOut_756, a(10)=>MultiplierOut_755, a(9)=>
      MultiplierOut_754, a(8)=>MultiplierOut_753, a(7)=>MultiplierOut_752, 
      a(6)=>MultiplierOut_751, a(5)=>MultiplierOut_750, a(4)=>
      MultiplierOut_749, a(3)=>MultiplierOut_748, a(2)=>MultiplierOut_747, 
      a(1)=>MultiplierOut_746, a(0)=>MultiplierOut_745, b(15)=>
      MultiplierOut_792, b(14)=>MultiplierOut_791, b(13)=>MultiplierOut_790, 
      b(12)=>MultiplierOut_789, b(11)=>MultiplierOut_788, b(10)=>
      MultiplierOut_787, b(9)=>MultiplierOut_786, b(8)=>MultiplierOut_785, 
      b(7)=>MultiplierOut_784, b(6)=>MultiplierOut_783, b(5)=>
      MultiplierOut_782, b(4)=>MultiplierOut_781, b(3)=>MultiplierOut_780, 
      b(2)=>MultiplierOut_779, b(1)=>MultiplierOut_778, b(0)=>
      MultiplierOut_777, cin=>GND0, s(15)=>AddOutputLvL1_191, s(14)=>
      AddOutputLvL1_190, s(13)=>AddOutputLvL1_189, s(12)=>AddOutputLvL1_188, 
      s(11)=>AddOutputLvL1_187, s(10)=>AddOutputLvL1_186, s(9)=>
      AddOutputLvL1_185, s(8)=>AddOutputLvL1_184, s(7)=>AddOutputLvL1_183, 
      s(6)=>AddOutputLvL1_182, s(5)=>AddOutputLvL1_181, s(4)=>
      AddOutputLvL1_180, s(3)=>AddOutputLvL1_179, s(2)=>AddOutputLvL1_178, 
      s(1)=>AddOutputLvL1_177, s(0)=>AddOutputLvL1_176, cout=>DANGLING(415)
   );
   adder14 : my_nadder_16 port map ( a(15)=>AddOutputLvL1_79, a(14)=>
      AddOutputLvL1_78, a(13)=>AddOutputLvL1_77, a(12)=>AddOutputLvL1_76, 
      a(11)=>AddOutputLvL1_75, a(10)=>AddOutputLvL1_74, a(9)=>
      AddOutputLvL1_73, a(8)=>AddOutputLvL1_72, a(7)=>AddOutputLvL1_71, a(6)
      =>AddOutputLvL1_70, a(5)=>AddOutputLvL1_69, a(4)=>AddOutputLvL1_68, 
      a(3)=>AddOutputLvL1_67, a(2)=>AddOutputLvL1_66, a(1)=>AddOutputLvL1_65, 
      a(0)=>AddOutputLvL1_64, b(15)=>AddOutputLvL1_95, b(14)=>
      AddOutputLvL1_94, b(13)=>AddOutputLvL1_93, b(12)=>AddOutputLvL1_92, 
      b(11)=>AddOutputLvL1_91, b(10)=>AddOutputLvL1_90, b(9)=>
      AddOutputLvL1_89, b(8)=>AddOutputLvL1_88, b(7)=>AddOutputLvL1_87, b(6)
      =>AddOutputLvL1_86, b(5)=>AddOutputLvL1_85, b(4)=>AddOutputLvL1_84, 
      b(3)=>AddOutputLvL1_83, b(2)=>AddOutputLvL1_82, b(1)=>AddOutputLvL1_81, 
      b(0)=>AddOutputLvL1_80, cin=>GND0, s(15)=>AddOutputLvL2_47, s(14)=>
      AddOutputLvL2_46, s(13)=>AddOutputLvL2_45, s(12)=>AddOutputLvL2_44, 
      s(11)=>AddOutputLvL2_43, s(10)=>AddOutputLvL2_42, s(9)=>
      AddOutputLvL2_41, s(8)=>AddOutputLvL2_40, s(7)=>AddOutputLvL2_39, s(6)
      =>AddOutputLvL2_38, s(5)=>AddOutputLvL2_37, s(4)=>AddOutputLvL2_36, 
      s(3)=>AddOutputLvL2_35, s(2)=>AddOutputLvL2_34, s(1)=>AddOutputLvL2_33, 
      s(0)=>AddOutputLvL2_32, cout=>DANGLING(416));
   adder15 : my_nadder_16 port map ( a(15)=>AddOutputLvL1_111, a(14)=>
      AddOutputLvL1_110, a(13)=>AddOutputLvL1_109, a(12)=>AddOutputLvL1_108, 
      a(11)=>AddOutputLvL1_107, a(10)=>AddOutputLvL1_106, a(9)=>
      AddOutputLvL1_105, a(8)=>AddOutputLvL1_104, a(7)=>AddOutputLvL1_103, 
      a(6)=>AddOutputLvL1_102, a(5)=>AddOutputLvL1_101, a(4)=>
      AddOutputLvL1_100, a(3)=>AddOutputLvL1_99, a(2)=>AddOutputLvL1_98, 
      a(1)=>AddOutputLvL1_97, a(0)=>AddOutputLvL1_96, b(15)=>
      AddOutputLvL1_127, b(14)=>AddOutputLvL1_126, b(13)=>AddOutputLvL1_125, 
      b(12)=>AddOutputLvL1_124, b(11)=>AddOutputLvL1_123, b(10)=>
      AddOutputLvL1_122, b(9)=>AddOutputLvL1_121, b(8)=>AddOutputLvL1_120, 
      b(7)=>AddOutputLvL1_119, b(6)=>AddOutputLvL1_118, b(5)=>
      AddOutputLvL1_117, b(4)=>AddOutputLvL1_116, b(3)=>AddOutputLvL1_115, 
      b(2)=>AddOutputLvL1_114, b(1)=>AddOutputLvL1_113, b(0)=>
      AddOutputLvL1_112, cin=>GND0, s(15)=>AddOutputLvL2_63, s(14)=>
      AddOutputLvL2_62, s(13)=>AddOutputLvL2_61, s(12)=>AddOutputLvL2_60, 
      s(11)=>AddOutputLvL2_59, s(10)=>AddOutputLvL2_58, s(9)=>
      AddOutputLvL2_57, s(8)=>AddOutputLvL2_56, s(7)=>AddOutputLvL2_55, s(6)
      =>AddOutputLvL2_54, s(5)=>AddOutputLvL2_53, s(4)=>AddOutputLvL2_52, 
      s(3)=>AddOutputLvL2_51, s(2)=>AddOutputLvL2_50, s(1)=>AddOutputLvL2_49, 
      s(0)=>AddOutputLvL2_48, cout=>DANGLING(417));
   adder16 : my_nadder_16 port map ( a(15)=>AddOutputLvL1_143, a(14)=>
      AddOutputLvL1_142, a(13)=>AddOutputLvL1_141, a(12)=>AddOutputLvL1_140, 
      a(11)=>AddOutputLvL1_139, a(10)=>AddOutputLvL1_138, a(9)=>
      AddOutputLvL1_137, a(8)=>AddOutputLvL1_136, a(7)=>AddOutputLvL1_135, 
      a(6)=>AddOutputLvL1_134, a(5)=>AddOutputLvL1_133, a(4)=>
      AddOutputLvL1_132, a(3)=>AddOutputLvL1_131, a(2)=>AddOutputLvL1_130, 
      a(1)=>AddOutputLvL1_129, a(0)=>AddOutputLvL1_128, b(15)=>
      AddOutputLvL1_159, b(14)=>AddOutputLvL1_158, b(13)=>AddOutputLvL1_157, 
      b(12)=>AddOutputLvL1_156, b(11)=>AddOutputLvL1_155, b(10)=>
      AddOutputLvL1_154, b(9)=>AddOutputLvL1_153, b(8)=>AddOutputLvL1_152, 
      b(7)=>AddOutputLvL1_151, b(6)=>AddOutputLvL1_150, b(5)=>
      AddOutputLvL1_149, b(4)=>AddOutputLvL1_148, b(3)=>AddOutputLvL1_147, 
      b(2)=>AddOutputLvL1_146, b(1)=>AddOutputLvL1_145, b(0)=>
      AddOutputLvL1_144, cin=>GND0, s(15)=>AddOutputLvL2_79, s(14)=>
      AddOutputLvL2_78, s(13)=>AddOutputLvL2_77, s(12)=>AddOutputLvL2_76, 
      s(11)=>AddOutputLvL2_75, s(10)=>AddOutputLvL2_74, s(9)=>
      AddOutputLvL2_73, s(8)=>AddOutputLvL2_72, s(7)=>AddOutputLvL2_71, s(6)
      =>AddOutputLvL2_70, s(5)=>AddOutputLvL2_69, s(4)=>AddOutputLvL2_68, 
      s(3)=>AddOutputLvL2_67, s(2)=>AddOutputLvL2_66, s(1)=>AddOutputLvL2_65, 
      s(0)=>AddOutputLvL2_64, cout=>DANGLING(418));
   adder17 : my_nadder_16 port map ( a(15)=>AddOutputLvL1_175, a(14)=>
      AddOutputLvL1_174, a(13)=>AddOutputLvL1_173, a(12)=>AddOutputLvL1_172, 
      a(11)=>AddOutputLvL1_171, a(10)=>AddOutputLvL1_170, a(9)=>
      AddOutputLvL1_169, a(8)=>AddOutputLvL1_168, a(7)=>AddOutputLvL1_167, 
      a(6)=>AddOutputLvL1_166, a(5)=>AddOutputLvL1_165, a(4)=>
      AddOutputLvL1_164, a(3)=>AddOutputLvL1_163, a(2)=>AddOutputLvL1_162, 
      a(1)=>AddOutputLvL1_161, a(0)=>AddOutputLvL1_160, b(15)=>
      AddOutputLvL1_191, b(14)=>AddOutputLvL1_190, b(13)=>AddOutputLvL1_189, 
      b(12)=>AddOutputLvL1_188, b(11)=>AddOutputLvL1_187, b(10)=>
      AddOutputLvL1_186, b(9)=>AddOutputLvL1_185, b(8)=>AddOutputLvL1_184, 
      b(7)=>AddOutputLvL1_183, b(6)=>AddOutputLvL1_182, b(5)=>
      AddOutputLvL1_181, b(4)=>AddOutputLvL1_180, b(3)=>AddOutputLvL1_179, 
      b(2)=>AddOutputLvL1_178, b(1)=>AddOutputLvL1_177, b(0)=>
      AddOutputLvL1_176, cin=>GND0, s(15)=>AddOutputLvL2_95, s(14)=>
      AddOutputLvL2_94, s(13)=>AddOutputLvL2_93, s(12)=>AddOutputLvL2_92, 
      s(11)=>AddOutputLvL2_91, s(10)=>AddOutputLvL2_90, s(9)=>
      AddOutputLvL2_89, s(8)=>AddOutputLvL2_88, s(7)=>AddOutputLvL2_87, s(6)
      =>AddOutputLvL2_86, s(5)=>AddOutputLvL2_85, s(4)=>AddOutputLvL2_84, 
      s(3)=>AddOutputLvL2_83, s(2)=>AddOutputLvL2_82, s(1)=>AddOutputLvL2_81, 
      s(0)=>AddOutputLvL2_80, cout=>DANGLING(419));
   adder19 : my_nadder_16 port map ( a(15)=>AddOutputLvL2_47, a(14)=>
      AddOutputLvL2_46, a(13)=>AddOutputLvL2_45, a(12)=>AddOutputLvL2_44, 
      a(11)=>AddOutputLvL2_43, a(10)=>AddOutputLvL2_42, a(9)=>
      AddOutputLvL2_41, a(8)=>AddOutputLvL2_40, a(7)=>AddOutputLvL2_39, a(6)
      =>AddOutputLvL2_38, a(5)=>AddOutputLvL2_37, a(4)=>AddOutputLvL2_36, 
      a(3)=>AddOutputLvL2_35, a(2)=>AddOutputLvL2_34, a(1)=>AddOutputLvL2_33, 
      a(0)=>AddOutputLvL2_32, b(15)=>AddOutputLvL2_63, b(14)=>
      AddOutputLvL2_62, b(13)=>AddOutputLvL2_61, b(12)=>AddOutputLvL2_60, 
      b(11)=>AddOutputLvL2_59, b(10)=>AddOutputLvL2_58, b(9)=>
      AddOutputLvL2_57, b(8)=>AddOutputLvL2_56, b(7)=>AddOutputLvL2_55, b(6)
      =>AddOutputLvL2_54, b(5)=>AddOutputLvL2_53, b(4)=>AddOutputLvL2_52, 
      b(3)=>AddOutputLvL2_51, b(2)=>AddOutputLvL2_50, b(1)=>AddOutputLvL2_49, 
      b(0)=>AddOutputLvL2_48, cin=>GND0, s(15)=>AddOutputLvL3_31, s(14)=>
      AddOutputLvL3_30, s(13)=>AddOutputLvL3_29, s(12)=>AddOutputLvL3_28, 
      s(11)=>AddOutputLvL3_27, s(10)=>AddOutputLvL3_26, s(9)=>
      AddOutputLvL3_25, s(8)=>AddOutputLvL3_24, s(7)=>AddOutputLvL3_23, s(6)
      =>AddOutputLvL3_22, s(5)=>AddOutputLvL3_21, s(4)=>AddOutputLvL3_20, 
      s(3)=>AddOutputLvL3_19, s(2)=>AddOutputLvL3_18, s(1)=>AddOutputLvL3_17, 
      s(0)=>AddOutputLvL3_16, cout=>DANGLING(420));
   adder20 : my_nadder_16 port map ( a(15)=>AddOutputLvL2_79, a(14)=>
      AddOutputLvL2_78, a(13)=>AddOutputLvL2_77, a(12)=>AddOutputLvL2_76, 
      a(11)=>AddOutputLvL2_75, a(10)=>AddOutputLvL2_74, a(9)=>
      AddOutputLvL2_73, a(8)=>AddOutputLvL2_72, a(7)=>AddOutputLvL2_71, a(6)
      =>AddOutputLvL2_70, a(5)=>AddOutputLvL2_69, a(4)=>AddOutputLvL2_68, 
      a(3)=>AddOutputLvL2_67, a(2)=>AddOutputLvL2_66, a(1)=>AddOutputLvL2_65, 
      a(0)=>AddOutputLvL2_64, b(15)=>AddOutputLvL2_95, b(14)=>
      AddOutputLvL2_94, b(13)=>AddOutputLvL2_93, b(12)=>AddOutputLvL2_92, 
      b(11)=>AddOutputLvL2_91, b(10)=>AddOutputLvL2_90, b(9)=>
      AddOutputLvL2_89, b(8)=>AddOutputLvL2_88, b(7)=>AddOutputLvL2_87, b(6)
      =>AddOutputLvL2_86, b(5)=>AddOutputLvL2_85, b(4)=>AddOutputLvL2_84, 
      b(3)=>AddOutputLvL2_83, b(2)=>AddOutputLvL2_82, b(1)=>AddOutputLvL2_81, 
      b(0)=>AddOutputLvL2_80, cin=>GND0, s(15)=>AddOutputLvL3_47, s(14)=>
      AddOutputLvL3_46, s(13)=>AddOutputLvL3_45, s(12)=>AddOutputLvL3_44, 
      s(11)=>AddOutputLvL3_43, s(10)=>AddOutputLvL3_42, s(9)=>
      AddOutputLvL3_41, s(8)=>AddOutputLvL3_40, s(7)=>AddOutputLvL3_39, s(6)
      =>AddOutputLvL3_38, s(5)=>AddOutputLvL3_37, s(4)=>AddOutputLvL3_36, 
      s(3)=>AddOutputLvL3_35, s(2)=>AddOutputLvL3_34, s(1)=>AddOutputLvL3_33, 
      s(0)=>AddOutputLvL3_32, cout=>DANGLING(421));
   adder22 : my_nadder_16 port map ( a(15)=>AddOutputLvL3_31, a(14)=>
      AddOutputLvL3_30, a(13)=>AddOutputLvL3_29, a(12)=>AddOutputLvL3_28, 
      a(11)=>AddOutputLvL3_27, a(10)=>AddOutputLvL3_26, a(9)=>
      AddOutputLvL3_25, a(8)=>AddOutputLvL3_24, a(7)=>AddOutputLvL3_23, a(6)
      =>AddOutputLvL3_22, a(5)=>AddOutputLvL3_21, a(4)=>AddOutputLvL3_20, 
      a(3)=>AddOutputLvL3_19, a(2)=>AddOutputLvL3_18, a(1)=>AddOutputLvL3_17, 
      a(0)=>AddOutputLvL3_16, b(15)=>AddOutputLvL3_47, b(14)=>
      AddOutputLvL3_46, b(13)=>AddOutputLvL3_45, b(12)=>AddOutputLvL3_44, 
      b(11)=>AddOutputLvL3_43, b(10)=>AddOutputLvL3_42, b(9)=>
      AddOutputLvL3_41, b(8)=>AddOutputLvL3_40, b(7)=>AddOutputLvL3_39, b(6)
      =>AddOutputLvL3_38, b(5)=>AddOutputLvL3_37, b(4)=>AddOutputLvL3_36, 
      b(3)=>AddOutputLvL3_35, b(2)=>AddOutputLvL3_34, b(1)=>AddOutputLvL3_33, 
      b(0)=>AddOutputLvL3_32, cin=>GND0, s(15)=>AddOut55_15, s(14)=>
      AddOut55_14, s(13)=>AddOut55_13, s(12)=>AddOut55_12, s(11)=>
      AddOut55_11, s(10)=>AddOut55_10, s(9)=>AddOut55_9, s(8)=>AddOut55_8, 
      s(7)=>AddOut55_7, s(6)=>AddOut55_6, s(5)=>AddOut55_5, s(4)=>AddOut55_4, 
      s(3)=>AddOut55_3, s(2)=>AddOut55_2, s(1)=>AddOut55_1, s(0)=>AddOut55_0, 
      cout=>DANGLING(422));
   adder23 : my_nadder_16 port map ( a(15)=>AddOut55_15, a(14)=>AddOut55_14, 
      a(13)=>AddOut55_13, a(12)=>AddOut55_12, a(11)=>AddOut55_11, a(10)=>
      AddOut55_10, a(9)=>AddOut55_9, a(8)=>AddOut55_8, a(7)=>AddOut55_7, 
      a(6)=>AddOut55_6, a(5)=>AddOut55_5, a(4)=>AddOut55_4, a(3)=>AddOut55_3, 
      a(2)=>AddOut55_2, a(1)=>AddOut55_1, a(0)=>AddOut55_0, b(15)=>
      AddOut33_15, b(14)=>AddOut33_14, b(13)=>AddOut33_13, b(12)=>
      AddOut33_12, b(11)=>AddOut33_11, b(10)=>AddOut33_10, b(9)=>AddOut33_9, 
      b(8)=>AddOut33_8, b(7)=>AddOut33_7, b(6)=>AddOut33_6, b(5)=>AddOut33_5, 
      b(4)=>AddOut33_4, b(3)=>AddOut33_3, b(2)=>AddOut33_2, b(1)=>AddOut33_1, 
      b(0)=>AddOut33_0, cin=>GND0, s(15)=>Final55_15, s(14)=>Final55_14, 
      s(13)=>Final55_13, s(12)=>Final55_12, s(11)=>Final55_11, s(10)=>
      Final55_10, s(9)=>Final55_9, s(8)=>Final55_8, s(7)=>Final55_7, s(6)=>
      Final55_6, s(5)=>Final55_5, s(4)=>Final55_4, s(3)=>Final55_3, s(2)=>
      Final55_2, s(1)=>Final55_1, s(0)=>Final55_0, cout=>DANGLING(423));
   EndCounter : Counter_3 port map ( enable=>CountereEN, reset=>CountereRST, 
      clk=>CLK, load=>GND0, output(2)=>CounterOut_2, output(1)=>CounterOut_1, 
      output(0)=>CounterOut_0, input(2)=>GND0, input(1)=>GND0, input(0)=>
      GND0);
   ix6941 : fake_gnd port map ( Y=>GND0);
   ix3555 : or02 port map ( Y=>CountereRST, A0=>nx3552, A1=>RST);
   ix3553 : nor03_2x port map ( Y=>nx3552, A0=>CounterOut_0, A1=>nx7936, A2
      =>CounterOut_1);
   ix7937 : inv01 port map ( Y=>nx7936, A=>CounterOut_2);
   ix3571 : nor02ii port map ( Y=>CountereEN, A0=>ACK_EXMPLR, A1=>
      current_state(7));
   reg_ACKC_dup_1 : dffs_ni port map ( Q=>ACK_EXMPLR, QB=>OPEN, D=>GND0, CLK
      =>CLK, S=>nx3562);
   ix3563 : and03 port map ( Y=>nx3562, A0=>CounterOut_0, A1=>nx7936, A2=>
      CounterOut_1);
   ix3425 : mux21_ni port map ( Y=>SecondInputToMult_48, A0=>OutputImg1(0), 
      A1=>OutputImg0(48), S0=>nx8858);
   ix3433 : mux21_ni port map ( Y=>SecondInputToMult_49, A0=>OutputImg1(1), 
      A1=>OutputImg0(49), S0=>nx8858);
   ix3441 : mux21_ni port map ( Y=>SecondInputToMult_50, A0=>OutputImg1(2), 
      A1=>OutputImg0(50), S0=>nx8858);
   ix3449 : mux21_ni port map ( Y=>SecondInputToMult_51, A0=>OutputImg1(3), 
      A1=>OutputImg0(51), S0=>nx8858);
   ix3457 : mux21_ni port map ( Y=>SecondInputToMult_52, A0=>OutputImg1(4), 
      A1=>OutputImg0(52), S0=>nx8858);
   ix3465 : mux21_ni port map ( Y=>SecondInputToMult_53, A0=>OutputImg1(5), 
      A1=>OutputImg0(53), S0=>nx8858);
   ix3473 : mux21_ni port map ( Y=>SecondInputToMult_54, A0=>OutputImg1(6), 
      A1=>OutputImg0(54), S0=>nx8858);
   ix3481 : mux21_ni port map ( Y=>SecondInputToMult_55, A0=>OutputImg1(7), 
      A1=>OutputImg0(55), S0=>nx8860);
   ix3489 : mux21_ni port map ( Y=>SecondInputToMult_56, A0=>OutputImg1(8), 
      A1=>OutputImg0(56), S0=>nx8860);
   ix3497 : mux21_ni port map ( Y=>SecondInputToMult_57, A0=>OutputImg1(9), 
      A1=>OutputImg0(57), S0=>nx8860);
   ix3505 : mux21_ni port map ( Y=>SecondInputToMult_58, A0=>OutputImg1(10), 
      A1=>OutputImg0(58), S0=>nx8860);
   ix3513 : mux21_ni port map ( Y=>SecondInputToMult_59, A0=>OutputImg1(11), 
      A1=>OutputImg0(59), S0=>nx8860);
   ix3521 : mux21_ni port map ( Y=>SecondInputToMult_60, A0=>OutputImg1(12), 
      A1=>OutputImg0(60), S0=>nx8860);
   ix3529 : mux21_ni port map ( Y=>SecondInputToMult_61, A0=>OutputImg1(13), 
      A1=>OutputImg0(61), S0=>nx8860);
   ix3537 : mux21_ni port map ( Y=>SecondInputToMult_62, A0=>OutputImg1(14), 
      A1=>OutputImg0(62), S0=>nx8862);
   ix3545 : mux21_ni port map ( Y=>SecondInputToMult_63, A0=>OutputImg1(15), 
      A1=>OutputImg0(63), S0=>nx8862);
   ix3297 : mux21_ni port map ( Y=>SecondInputToMult_64, A0=>OutputImg1(16), 
      A1=>OutputImg0(64), S0=>nx8862);
   ix3305 : mux21_ni port map ( Y=>SecondInputToMult_65, A0=>OutputImg1(17), 
      A1=>OutputImg0(65), S0=>nx8862);
   ix3313 : mux21_ni port map ( Y=>SecondInputToMult_66, A0=>OutputImg1(18), 
      A1=>OutputImg0(66), S0=>nx8862);
   ix3321 : mux21_ni port map ( Y=>SecondInputToMult_67, A0=>OutputImg1(19), 
      A1=>OutputImg0(67), S0=>nx8862);
   ix3329 : mux21_ni port map ( Y=>SecondInputToMult_68, A0=>OutputImg1(20), 
      A1=>OutputImg0(68), S0=>nx8862);
   ix3337 : mux21_ni port map ( Y=>SecondInputToMult_69, A0=>OutputImg1(21), 
      A1=>OutputImg0(69), S0=>nx8864);
   ix3345 : mux21_ni port map ( Y=>SecondInputToMult_70, A0=>OutputImg1(22), 
      A1=>OutputImg0(70), S0=>nx8864);
   ix3353 : mux21_ni port map ( Y=>SecondInputToMult_71, A0=>OutputImg1(23), 
      A1=>OutputImg0(71), S0=>nx8864);
   ix3361 : mux21_ni port map ( Y=>SecondInputToMult_72, A0=>OutputImg1(24), 
      A1=>OutputImg0(72), S0=>nx8864);
   ix3369 : mux21_ni port map ( Y=>SecondInputToMult_73, A0=>OutputImg1(25), 
      A1=>OutputImg0(73), S0=>nx8864);
   ix3377 : mux21_ni port map ( Y=>SecondInputToMult_74, A0=>OutputImg1(26), 
      A1=>OutputImg0(74), S0=>nx8864);
   ix3385 : mux21_ni port map ( Y=>SecondInputToMult_75, A0=>OutputImg1(27), 
      A1=>OutputImg0(75), S0=>nx8864);
   ix3393 : mux21_ni port map ( Y=>SecondInputToMult_76, A0=>OutputImg1(28), 
      A1=>OutputImg0(76), S0=>nx8866);
   ix3401 : mux21_ni port map ( Y=>SecondInputToMult_77, A0=>OutputImg1(29), 
      A1=>OutputImg0(77), S0=>nx8866);
   ix3409 : mux21_ni port map ( Y=>SecondInputToMult_78, A0=>OutputImg1(30), 
      A1=>OutputImg0(78), S0=>nx8866);
   ix3417 : mux21_ni port map ( Y=>SecondInputToMult_79, A0=>OutputImg1(31), 
      A1=>OutputImg0(79), S0=>nx8866);
   ix3169 : mux21_ni port map ( Y=>SecondInputToMult_80, A0=>OutputImg1(32), 
      A1=>OutputImg1(0), S0=>nx8866);
   ix3177 : mux21_ni port map ( Y=>SecondInputToMult_81, A0=>OutputImg1(33), 
      A1=>OutputImg1(1), S0=>nx8866);
   ix3185 : mux21_ni port map ( Y=>SecondInputToMult_82, A0=>OutputImg1(34), 
      A1=>OutputImg1(2), S0=>nx8866);
   ix3193 : mux21_ni port map ( Y=>SecondInputToMult_83, A0=>OutputImg1(35), 
      A1=>OutputImg1(3), S0=>nx8868);
   ix3201 : mux21_ni port map ( Y=>SecondInputToMult_84, A0=>OutputImg1(36), 
      A1=>OutputImg1(4), S0=>nx8868);
   ix3209 : mux21_ni port map ( Y=>SecondInputToMult_85, A0=>OutputImg1(37), 
      A1=>OutputImg1(5), S0=>nx8868);
   ix3217 : mux21_ni port map ( Y=>SecondInputToMult_86, A0=>OutputImg1(38), 
      A1=>OutputImg1(6), S0=>nx8868);
   ix3225 : mux21_ni port map ( Y=>SecondInputToMult_87, A0=>OutputImg1(39), 
      A1=>OutputImg1(7), S0=>nx8868);
   ix3233 : mux21_ni port map ( Y=>SecondInputToMult_88, A0=>OutputImg1(40), 
      A1=>OutputImg1(8), S0=>nx8868);
   ix3241 : mux21_ni port map ( Y=>SecondInputToMult_89, A0=>OutputImg1(41), 
      A1=>OutputImg1(9), S0=>nx8868);
   ix3249 : mux21_ni port map ( Y=>SecondInputToMult_90, A0=>OutputImg1(42), 
      A1=>OutputImg1(10), S0=>nx8870);
   ix3257 : mux21_ni port map ( Y=>SecondInputToMult_91, A0=>OutputImg1(43), 
      A1=>OutputImg1(11), S0=>nx8870);
   ix3265 : mux21_ni port map ( Y=>SecondInputToMult_92, A0=>OutputImg1(44), 
      A1=>OutputImg1(12), S0=>nx8870);
   ix3273 : mux21_ni port map ( Y=>SecondInputToMult_93, A0=>OutputImg1(45), 
      A1=>OutputImg1(13), S0=>nx8870);
   ix3281 : mux21_ni port map ( Y=>SecondInputToMult_94, A0=>OutputImg1(46), 
      A1=>OutputImg1(14), S0=>nx8870);
   ix3289 : mux21_ni port map ( Y=>SecondInputToMult_95, A0=>OutputImg1(47), 
      A1=>OutputImg1(15), S0=>nx8870);
   ix3041 : mux21_ni port map ( Y=>SecondInputToMult_96, A0=>OutputImg2(0), 
      A1=>OutputImg1(16), S0=>nx8870);
   ix3049 : mux21_ni port map ( Y=>SecondInputToMult_97, A0=>OutputImg2(1), 
      A1=>OutputImg1(17), S0=>nx8872);
   ix3057 : mux21_ni port map ( Y=>SecondInputToMult_98, A0=>OutputImg2(2), 
      A1=>OutputImg1(18), S0=>nx8872);
   ix3065 : mux21_ni port map ( Y=>SecondInputToMult_99, A0=>OutputImg2(3), 
      A1=>OutputImg1(19), S0=>nx8872);
   ix3073 : mux21_ni port map ( Y=>SecondInputToMult_100, A0=>OutputImg2(4), 
      A1=>OutputImg1(20), S0=>nx8872);
   ix3081 : mux21_ni port map ( Y=>SecondInputToMult_101, A0=>OutputImg2(5), 
      A1=>OutputImg1(21), S0=>nx8872);
   ix3089 : mux21_ni port map ( Y=>SecondInputToMult_102, A0=>OutputImg2(6), 
      A1=>OutputImg1(22), S0=>nx8872);
   ix3097 : mux21_ni port map ( Y=>SecondInputToMult_103, A0=>OutputImg2(7), 
      A1=>OutputImg1(23), S0=>nx8872);
   ix3105 : mux21_ni port map ( Y=>SecondInputToMult_104, A0=>OutputImg2(8), 
      A1=>OutputImg1(24), S0=>nx8874);
   ix3113 : mux21_ni port map ( Y=>SecondInputToMult_105, A0=>OutputImg2(9), 
      A1=>OutputImg1(25), S0=>nx8874);
   ix3121 : mux21_ni port map ( Y=>SecondInputToMult_106, A0=>OutputImg2(10), 
      A1=>OutputImg1(26), S0=>nx8874);
   ix3129 : mux21_ni port map ( Y=>SecondInputToMult_107, A0=>OutputImg2(11), 
      A1=>OutputImg1(27), S0=>nx8874);
   ix3137 : mux21_ni port map ( Y=>SecondInputToMult_108, A0=>OutputImg2(12), 
      A1=>OutputImg1(28), S0=>nx8874);
   ix3145 : mux21_ni port map ( Y=>SecondInputToMult_109, A0=>OutputImg2(13), 
      A1=>OutputImg1(29), S0=>nx8874);
   ix3153 : mux21_ni port map ( Y=>SecondInputToMult_110, A0=>OutputImg2(14), 
      A1=>OutputImg1(30), S0=>nx8874);
   ix3161 : mux21_ni port map ( Y=>SecondInputToMult_111, A0=>OutputImg2(15), 
      A1=>OutputImg1(31), S0=>nx8876);
   ix2913 : mux21_ni port map ( Y=>SecondInputToMult_112, A0=>OutputImg2(16), 
      A1=>OutputImg1(32), S0=>nx8876);
   ix2921 : mux21_ni port map ( Y=>SecondInputToMult_113, A0=>OutputImg2(17), 
      A1=>OutputImg1(33), S0=>nx8876);
   ix2929 : mux21_ni port map ( Y=>SecondInputToMult_114, A0=>OutputImg2(18), 
      A1=>OutputImg1(34), S0=>nx8876);
   ix2937 : mux21_ni port map ( Y=>SecondInputToMult_115, A0=>OutputImg2(19), 
      A1=>OutputImg1(35), S0=>nx8876);
   ix2945 : mux21_ni port map ( Y=>SecondInputToMult_116, A0=>OutputImg2(20), 
      A1=>OutputImg1(36), S0=>nx8876);
   ix2953 : mux21_ni port map ( Y=>SecondInputToMult_117, A0=>OutputImg2(21), 
      A1=>OutputImg1(37), S0=>nx8876);
   ix2961 : mux21_ni port map ( Y=>SecondInputToMult_118, A0=>OutputImg2(22), 
      A1=>OutputImg1(38), S0=>nx8878);
   ix2969 : mux21_ni port map ( Y=>SecondInputToMult_119, A0=>OutputImg2(23), 
      A1=>OutputImg1(39), S0=>nx8878);
   ix2977 : mux21_ni port map ( Y=>SecondInputToMult_120, A0=>OutputImg2(24), 
      A1=>OutputImg1(40), S0=>nx8878);
   ix2985 : mux21_ni port map ( Y=>SecondInputToMult_121, A0=>OutputImg2(25), 
      A1=>OutputImg1(41), S0=>nx8878);
   ix2993 : mux21_ni port map ( Y=>SecondInputToMult_122, A0=>OutputImg2(26), 
      A1=>OutputImg1(42), S0=>nx8878);
   ix3001 : mux21_ni port map ( Y=>SecondInputToMult_123, A0=>OutputImg2(27), 
      A1=>OutputImg1(43), S0=>nx8878);
   ix3009 : mux21_ni port map ( Y=>SecondInputToMult_124, A0=>OutputImg2(28), 
      A1=>OutputImg1(44), S0=>nx8878);
   ix3017 : mux21_ni port map ( Y=>SecondInputToMult_125, A0=>OutputImg2(29), 
      A1=>OutputImg1(45), S0=>nx8880);
   ix3025 : mux21_ni port map ( Y=>SecondInputToMult_126, A0=>OutputImg2(30), 
      A1=>OutputImg1(46), S0=>nx8880);
   ix3033 : mux21_ni port map ( Y=>SecondInputToMult_127, A0=>OutputImg2(31), 
      A1=>OutputImg1(47), S0=>nx8880);
   ix2785 : mux21_ni port map ( Y=>SecondInputToMult_128, A0=>OutputImg2(32), 
      A1=>OutputImg1(48), S0=>nx8880);
   ix2793 : mux21_ni port map ( Y=>SecondInputToMult_129, A0=>OutputImg2(33), 
      A1=>OutputImg1(49), S0=>nx8880);
   ix2801 : mux21_ni port map ( Y=>SecondInputToMult_130, A0=>OutputImg2(34), 
      A1=>OutputImg1(50), S0=>nx8880);
   ix2809 : mux21_ni port map ( Y=>SecondInputToMult_131, A0=>OutputImg2(35), 
      A1=>OutputImg1(51), S0=>nx8880);
   ix2817 : mux21_ni port map ( Y=>SecondInputToMult_132, A0=>OutputImg2(36), 
      A1=>OutputImg1(52), S0=>nx8882);
   ix2825 : mux21_ni port map ( Y=>SecondInputToMult_133, A0=>OutputImg2(37), 
      A1=>OutputImg1(53), S0=>nx8882);
   ix2833 : mux21_ni port map ( Y=>SecondInputToMult_134, A0=>OutputImg2(38), 
      A1=>OutputImg1(54), S0=>nx8882);
   ix2841 : mux21_ni port map ( Y=>SecondInputToMult_135, A0=>OutputImg2(39), 
      A1=>OutputImg1(55), S0=>nx8882);
   ix2849 : mux21_ni port map ( Y=>SecondInputToMult_136, A0=>OutputImg2(40), 
      A1=>OutputImg1(56), S0=>nx8882);
   ix2857 : mux21_ni port map ( Y=>SecondInputToMult_137, A0=>OutputImg2(41), 
      A1=>OutputImg1(57), S0=>nx8882);
   ix2865 : mux21_ni port map ( Y=>SecondInputToMult_138, A0=>OutputImg2(42), 
      A1=>OutputImg1(58), S0=>nx8882);
   ix2873 : mux21_ni port map ( Y=>SecondInputToMult_139, A0=>OutputImg2(43), 
      A1=>OutputImg1(59), S0=>nx8884);
   ix2881 : mux21_ni port map ( Y=>SecondInputToMult_140, A0=>OutputImg2(44), 
      A1=>OutputImg1(60), S0=>nx8884);
   ix2889 : mux21_ni port map ( Y=>SecondInputToMult_141, A0=>OutputImg2(45), 
      A1=>OutputImg1(61), S0=>nx8884);
   ix2897 : mux21_ni port map ( Y=>SecondInputToMult_142, A0=>OutputImg2(46), 
      A1=>OutputImg1(62), S0=>nx8884);
   ix2905 : mux21_ni port map ( Y=>SecondInputToMult_143, A0=>OutputImg2(47), 
      A1=>OutputImg1(63), S0=>nx8884);
   ix2681 : ao22 port map ( Y=>FilterToAlu_0, A0=>outFilter0(0), A1=>nx8586, 
      B0=>outFilter1(0), B1=>nx8696);
   ix511 : nor02_2x port map ( Y=>nx510, A0=>nx8896, A1=>nx8852);
   ix2687 : ao22 port map ( Y=>FilterToAlu_1, A0=>outFilter0(1), A1=>nx8586, 
      B0=>outFilter1(1), B1=>nx8696);
   ix2693 : ao22 port map ( Y=>FilterToAlu_2, A0=>outFilter0(2), A1=>nx8586, 
      B0=>outFilter1(2), B1=>nx8696);
   ix2699 : ao22 port map ( Y=>FilterToAlu_3, A0=>outFilter0(3), A1=>nx8586, 
      B0=>outFilter1(3), B1=>nx8696);
   ix2705 : ao22 port map ( Y=>FilterToAlu_4, A0=>outFilter0(4), A1=>nx8586, 
      B0=>outFilter1(4), B1=>nx8696);
   ix2711 : ao22 port map ( Y=>FilterToAlu_5, A0=>outFilter0(5), A1=>nx8586, 
      B0=>outFilter1(5), B1=>nx8696);
   ix2717 : ao22 port map ( Y=>FilterToAlu_6, A0=>outFilter0(6), A1=>nx8586, 
      B0=>outFilter1(6), B1=>nx8696);
   ix2723 : ao22 port map ( Y=>FilterToAlu_7, A0=>outFilter0(7), A1=>nx8588, 
      B0=>outFilter1(7), B1=>nx8698);
   ix2729 : ao22 port map ( Y=>FilterToAlu_8, A0=>outFilter0(8), A1=>nx8588, 
      B0=>outFilter1(8), B1=>nx8698);
   ix505 : nand02 port map ( Y=>FilterToAlu_9, A0=>nx8052, A1=>nx8924);
   ix8053 : mux21 port map ( Y=>nx8052, A0=>outFilter0(9), A1=>outFilter1(9), 
      S0=>nx8896);
   ix2735 : ao22 port map ( Y=>FilterToAlu_10, A0=>outFilter0(10), A1=>
      nx8588, B0=>outFilter1(10), B1=>nx8698);
   ix2741 : ao22 port map ( Y=>FilterToAlu_11, A0=>outFilter0(11), A1=>
      nx8588, B0=>outFilter1(11), B1=>nx8698);
   ix2747 : ao22 port map ( Y=>FilterToAlu_12, A0=>outFilter0(12), A1=>
      nx8588, B0=>outFilter1(12), B1=>nx8698);
   ix2753 : ao22 port map ( Y=>FilterToAlu_13, A0=>outFilter0(13), A1=>
      nx8588, B0=>outFilter1(13), B1=>nx8698);
   ix2759 : ao22 port map ( Y=>FilterToAlu_14, A0=>outFilter0(14), A1=>
      nx8588, B0=>outFilter1(14), B1=>nx8698);
   ix2765 : ao22 port map ( Y=>FilterToAlu_15, A0=>outFilter0(15), A1=>
      nx8590, B0=>outFilter1(15), B1=>nx8700);
   ix2591 : ao22 port map ( Y=>FilterToAlu_16, A0=>outFilter0(16), A1=>
      nx8590, B0=>outFilter1(16), B1=>nx8700);
   ix2597 : ao22 port map ( Y=>FilterToAlu_17, A0=>outFilter0(17), A1=>
      nx8590, B0=>outFilter1(17), B1=>nx8700);
   ix2603 : ao22 port map ( Y=>FilterToAlu_18, A0=>outFilter0(18), A1=>
      nx8590, B0=>outFilter1(18), B1=>nx8700);
   ix2609 : ao22 port map ( Y=>FilterToAlu_19, A0=>outFilter0(19), A1=>
      nx8590, B0=>outFilter1(19), B1=>nx8700);
   ix2615 : ao22 port map ( Y=>FilterToAlu_20, A0=>outFilter0(20), A1=>
      nx8590, B0=>outFilter1(20), B1=>nx8700);
   ix2621 : ao22 port map ( Y=>FilterToAlu_21, A0=>outFilter0(21), A1=>
      nx8590, B0=>outFilter1(21), B1=>nx8700);
   ix2627 : ao22 port map ( Y=>FilterToAlu_22, A0=>outFilter0(22), A1=>
      nx8592, B0=>outFilter1(22), B1=>nx8702);
   ix2633 : ao22 port map ( Y=>FilterToAlu_23, A0=>outFilter0(23), A1=>
      nx8592, B0=>outFilter1(23), B1=>nx8702);
   ix2639 : ao22 port map ( Y=>FilterToAlu_24, A0=>outFilter0(24), A1=>
      nx8592, B0=>outFilter1(24), B1=>nx8702);
   ix495 : nand02 port map ( Y=>FilterToAlu_25, A0=>nx8072, A1=>nx8924);
   ix8073 : mux21 port map ( Y=>nx8072, A0=>outFilter0(25), A1=>
      outFilter1(25), S0=>nx8896);
   ix2645 : ao22 port map ( Y=>FilterToAlu_26, A0=>outFilter0(26), A1=>
      nx8592, B0=>outFilter1(26), B1=>nx8702);
   ix2651 : ao22 port map ( Y=>FilterToAlu_27, A0=>outFilter0(27), A1=>
      nx8592, B0=>outFilter1(27), B1=>nx8702);
   ix2657 : ao22 port map ( Y=>FilterToAlu_28, A0=>outFilter0(28), A1=>
      nx8592, B0=>outFilter1(28), B1=>nx8702);
   ix2663 : ao22 port map ( Y=>FilterToAlu_29, A0=>outFilter0(29), A1=>
      nx8592, B0=>outFilter1(29), B1=>nx8702);
   ix2669 : ao22 port map ( Y=>FilterToAlu_30, A0=>outFilter0(30), A1=>
      nx8594, B0=>outFilter1(30), B1=>nx8704);
   ix2675 : ao22 port map ( Y=>FilterToAlu_31, A0=>outFilter0(31), A1=>
      nx8594, B0=>outFilter1(31), B1=>nx8704);
   ix2501 : ao22 port map ( Y=>FilterToAlu_32, A0=>outFilter0(32), A1=>
      nx8594, B0=>outFilter1(32), B1=>nx8704);
   ix2507 : ao22 port map ( Y=>FilterToAlu_33, A0=>outFilter0(33), A1=>
      nx8594, B0=>outFilter1(33), B1=>nx8704);
   ix2513 : ao22 port map ( Y=>FilterToAlu_34, A0=>outFilter0(34), A1=>
      nx8594, B0=>outFilter1(34), B1=>nx8704);
   ix2519 : ao22 port map ( Y=>FilterToAlu_35, A0=>outFilter0(35), A1=>
      nx8594, B0=>outFilter1(35), B1=>nx8704);
   ix2525 : ao22 port map ( Y=>FilterToAlu_36, A0=>outFilter0(36), A1=>
      nx8594, B0=>outFilter1(36), B1=>nx8704);
   ix2531 : ao22 port map ( Y=>FilterToAlu_37, A0=>outFilter0(37), A1=>
      nx8596, B0=>outFilter1(37), B1=>nx8706);
   ix2537 : ao22 port map ( Y=>FilterToAlu_38, A0=>outFilter0(38), A1=>
      nx8596, B0=>outFilter1(38), B1=>nx8706);
   ix2543 : ao22 port map ( Y=>FilterToAlu_39, A0=>outFilter0(39), A1=>
      nx8596, B0=>outFilter1(39), B1=>nx8706);
   ix2549 : ao22 port map ( Y=>FilterToAlu_40, A0=>outFilter0(40), A1=>
      nx8596, B0=>outFilter1(40), B1=>nx8706);
   ix485 : nand02 port map ( Y=>FilterToAlu_41, A0=>nx8090, A1=>nx8924);
   ix8091 : mux21 port map ( Y=>nx8090, A0=>outFilter0(41), A1=>
      outFilter1(41), S0=>nx8896);
   ix2555 : ao22 port map ( Y=>FilterToAlu_42, A0=>outFilter0(42), A1=>
      nx8596, B0=>outFilter1(42), B1=>nx8706);
   ix2561 : ao22 port map ( Y=>FilterToAlu_43, A0=>outFilter0(43), A1=>
      nx8596, B0=>outFilter1(43), B1=>nx8706);
   ix2567 : ao22 port map ( Y=>FilterToAlu_44, A0=>outFilter0(44), A1=>
      nx8596, B0=>outFilter1(44), B1=>nx8706);
   ix2573 : ao22 port map ( Y=>FilterToAlu_45, A0=>outFilter0(45), A1=>
      nx8598, B0=>outFilter1(45), B1=>nx8708);
   ix2579 : ao22 port map ( Y=>FilterToAlu_46, A0=>outFilter0(46), A1=>
      nx8598, B0=>outFilter1(46), B1=>nx8708);
   ix2585 : ao22 port map ( Y=>FilterToAlu_47, A0=>outFilter0(47), A1=>
      nx8598, B0=>outFilter1(47), B1=>nx8708);
   ix2411 : ao22 port map ( Y=>FilterToAlu_48, A0=>outFilter0(48), A1=>
      nx8598, B0=>outFilter1(48), B1=>nx8708);
   ix2417 : ao22 port map ( Y=>FilterToAlu_49, A0=>outFilter0(49), A1=>
      nx8598, B0=>outFilter1(49), B1=>nx8708);
   ix2423 : ao22 port map ( Y=>FilterToAlu_50, A0=>outFilter0(50), A1=>
      nx8598, B0=>outFilter1(50), B1=>nx8708);
   ix2429 : ao22 port map ( Y=>FilterToAlu_51, A0=>outFilter0(51), A1=>
      nx8598, B0=>outFilter1(51), B1=>nx8708);
   ix2435 : ao22 port map ( Y=>FilterToAlu_52, A0=>outFilter0(52), A1=>
      nx8600, B0=>outFilter1(52), B1=>nx8710);
   ix2441 : ao22 port map ( Y=>FilterToAlu_53, A0=>outFilter0(53), A1=>
      nx8600, B0=>outFilter1(53), B1=>nx8710);
   ix2447 : ao22 port map ( Y=>FilterToAlu_54, A0=>outFilter0(54), A1=>
      nx8600, B0=>outFilter1(54), B1=>nx8710);
   ix2453 : ao22 port map ( Y=>FilterToAlu_55, A0=>outFilter0(55), A1=>
      nx8600, B0=>outFilter1(55), B1=>nx8710);
   ix2459 : ao22 port map ( Y=>FilterToAlu_56, A0=>outFilter0(56), A1=>
      nx8600, B0=>outFilter1(56), B1=>nx8710);
   ix475 : nand02 port map ( Y=>FilterToAlu_57, A0=>nx8108, A1=>nx8924);
   ix8109 : mux21 port map ( Y=>nx8108, A0=>outFilter0(57), A1=>
      outFilter1(57), S0=>nx8896);
   ix2465 : ao22 port map ( Y=>FilterToAlu_58, A0=>outFilter0(58), A1=>
      nx8600, B0=>outFilter1(58), B1=>nx8710);
   ix2471 : ao22 port map ( Y=>FilterToAlu_59, A0=>outFilter0(59), A1=>
      nx8600, B0=>outFilter1(59), B1=>nx8710);
   ix2477 : ao22 port map ( Y=>FilterToAlu_60, A0=>outFilter0(60), A1=>
      nx8602, B0=>outFilter1(60), B1=>nx8712);
   ix2483 : ao22 port map ( Y=>FilterToAlu_61, A0=>outFilter0(61), A1=>
      nx8602, B0=>outFilter1(61), B1=>nx8712);
   ix2489 : ao22 port map ( Y=>FilterToAlu_62, A0=>outFilter0(62), A1=>
      nx8602, B0=>outFilter1(62), B1=>nx8712);
   ix2495 : ao22 port map ( Y=>FilterToAlu_63, A0=>outFilter0(63), A1=>
      nx8602, B0=>outFilter1(63), B1=>nx8712);
   ix2321 : ao22 port map ( Y=>FilterToAlu_64, A0=>outFilter0(64), A1=>
      nx8602, B0=>outFilter1(64), B1=>nx8712);
   ix2327 : ao22 port map ( Y=>FilterToAlu_65, A0=>outFilter0(65), A1=>
      nx8602, B0=>outFilter1(65), B1=>nx8712);
   ix2333 : ao22 port map ( Y=>FilterToAlu_66, A0=>outFilter0(66), A1=>
      nx8602, B0=>outFilter1(66), B1=>nx8712);
   ix2339 : ao22 port map ( Y=>FilterToAlu_67, A0=>outFilter0(67), A1=>
      nx8604, B0=>outFilter1(67), B1=>nx8714);
   ix2345 : ao22 port map ( Y=>FilterToAlu_68, A0=>outFilter0(68), A1=>
      nx8604, B0=>outFilter1(68), B1=>nx8714);
   ix2351 : ao22 port map ( Y=>FilterToAlu_69, A0=>outFilter0(69), A1=>
      nx8604, B0=>outFilter1(69), B1=>nx8714);
   ix2357 : ao22 port map ( Y=>FilterToAlu_70, A0=>outFilter0(70), A1=>
      nx8604, B0=>outFilter1(70), B1=>nx8714);
   ix2363 : ao22 port map ( Y=>FilterToAlu_71, A0=>outFilter0(71), A1=>
      nx8604, B0=>outFilter1(71), B1=>nx8714);
   ix2369 : ao22 port map ( Y=>FilterToAlu_72, A0=>outFilter0(72), A1=>
      nx8604, B0=>outFilter1(72), B1=>nx8714);
   ix465 : nand02 port map ( Y=>FilterToAlu_73, A0=>nx8126, A1=>nx8924);
   ix8127 : mux21 port map ( Y=>nx8126, A0=>outFilter0(73), A1=>
      outFilter1(73), S0=>nx8896);
   ix2375 : ao22 port map ( Y=>FilterToAlu_74, A0=>outFilter0(74), A1=>
      nx8604, B0=>outFilter1(74), B1=>nx8714);
   ix2381 : ao22 port map ( Y=>FilterToAlu_75, A0=>outFilter0(75), A1=>
      nx8606, B0=>outFilter1(75), B1=>nx8716);
   ix2387 : ao22 port map ( Y=>FilterToAlu_76, A0=>outFilter0(76), A1=>
      nx8606, B0=>outFilter1(76), B1=>nx8716);
   ix2393 : ao22 port map ( Y=>FilterToAlu_77, A0=>outFilter0(77), A1=>
      nx8606, B0=>outFilter1(77), B1=>nx8716);
   ix2399 : ao22 port map ( Y=>FilterToAlu_78, A0=>outFilter0(78), A1=>
      nx8606, B0=>outFilter1(78), B1=>nx8716);
   ix2405 : ao22 port map ( Y=>FilterToAlu_79, A0=>outFilter0(79), A1=>
      nx8606, B0=>outFilter1(79), B1=>nx8716);
   ix2231 : ao22 port map ( Y=>FilterToAlu_80, A0=>outFilter0(80), A1=>
      nx8606, B0=>outFilter1(80), B1=>nx8716);
   ix2237 : ao22 port map ( Y=>FilterToAlu_81, A0=>outFilter0(81), A1=>
      nx8606, B0=>outFilter1(81), B1=>nx8716);
   ix2243 : ao22 port map ( Y=>FilterToAlu_82, A0=>outFilter0(82), A1=>
      nx8608, B0=>outFilter1(82), B1=>nx8718);
   ix2249 : ao22 port map ( Y=>FilterToAlu_83, A0=>outFilter0(83), A1=>
      nx8608, B0=>outFilter1(83), B1=>nx8718);
   ix2255 : ao22 port map ( Y=>FilterToAlu_84, A0=>outFilter0(84), A1=>
      nx8608, B0=>outFilter1(84), B1=>nx8718);
   ix2261 : ao22 port map ( Y=>FilterToAlu_85, A0=>outFilter0(85), A1=>
      nx8608, B0=>outFilter1(85), B1=>nx8718);
   ix2267 : ao22 port map ( Y=>FilterToAlu_86, A0=>outFilter0(86), A1=>
      nx8608, B0=>outFilter1(86), B1=>nx8718);
   ix2273 : ao22 port map ( Y=>FilterToAlu_87, A0=>outFilter0(87), A1=>
      nx8608, B0=>outFilter1(87), B1=>nx8718);
   ix2279 : ao22 port map ( Y=>FilterToAlu_88, A0=>outFilter0(88), A1=>
      nx8608, B0=>outFilter1(88), B1=>nx8718);
   ix455 : nand02 port map ( Y=>FilterToAlu_89, A0=>nx8144, A1=>nx8924);
   ix8145 : mux21 port map ( Y=>nx8144, A0=>outFilter0(89), A1=>
      outFilter1(89), S0=>nx8896);
   ix2285 : ao22 port map ( Y=>FilterToAlu_90, A0=>outFilter0(90), A1=>
      nx8610, B0=>outFilter1(90), B1=>nx8720);
   ix2291 : ao22 port map ( Y=>FilterToAlu_91, A0=>outFilter0(91), A1=>
      nx8610, B0=>outFilter1(91), B1=>nx8720);
   ix2297 : ao22 port map ( Y=>FilterToAlu_92, A0=>outFilter0(92), A1=>
      nx8610, B0=>outFilter1(92), B1=>nx8720);
   ix2303 : ao22 port map ( Y=>FilterToAlu_93, A0=>outFilter0(93), A1=>
      nx8610, B0=>outFilter1(93), B1=>nx8720);
   ix2309 : ao22 port map ( Y=>FilterToAlu_94, A0=>outFilter0(94), A1=>
      nx8610, B0=>outFilter1(94), B1=>nx8720);
   ix2315 : ao22 port map ( Y=>FilterToAlu_95, A0=>outFilter0(95), A1=>
      nx8610, B0=>outFilter1(95), B1=>nx8720);
   ix2141 : ao22 port map ( Y=>FilterToAlu_96, A0=>outFilter0(96), A1=>
      nx8610, B0=>outFilter1(96), B1=>nx8720);
   ix2147 : ao22 port map ( Y=>FilterToAlu_97, A0=>outFilter0(97), A1=>
      nx8612, B0=>outFilter1(97), B1=>nx8722);
   ix2153 : ao22 port map ( Y=>FilterToAlu_98, A0=>outFilter0(98), A1=>
      nx8612, B0=>outFilter1(98), B1=>nx8722);
   ix2159 : ao22 port map ( Y=>FilterToAlu_99, A0=>outFilter0(99), A1=>
      nx8612, B0=>outFilter1(99), B1=>nx8722);
   ix2165 : ao22 port map ( Y=>FilterToAlu_100, A0=>outFilter0(100), A1=>
      nx8612, B0=>outFilter1(100), B1=>nx8722);
   ix2171 : ao22 port map ( Y=>FilterToAlu_101, A0=>outFilter0(101), A1=>
      nx8612, B0=>outFilter1(101), B1=>nx8722);
   ix2177 : ao22 port map ( Y=>FilterToAlu_102, A0=>outFilter0(102), A1=>
      nx8612, B0=>outFilter1(102), B1=>nx8722);
   ix2183 : ao22 port map ( Y=>FilterToAlu_103, A0=>outFilter0(103), A1=>
      nx8612, B0=>outFilter1(103), B1=>nx8722);
   ix2189 : ao22 port map ( Y=>FilterToAlu_104, A0=>outFilter0(104), A1=>
      nx8614, B0=>outFilter1(104), B1=>nx8724);
   ix445 : nand02 port map ( Y=>FilterToAlu_105, A0=>nx8162, A1=>nx8924);
   ix8163 : mux21 port map ( Y=>nx8162, A0=>outFilter0(105), A1=>
      outFilter1(105), S0=>nx8898);
   ix2195 : ao22 port map ( Y=>FilterToAlu_106, A0=>outFilter0(106), A1=>
      nx8614, B0=>outFilter1(106), B1=>nx8724);
   ix2201 : ao22 port map ( Y=>FilterToAlu_107, A0=>outFilter0(107), A1=>
      nx8614, B0=>outFilter1(107), B1=>nx8724);
   ix2207 : ao22 port map ( Y=>FilterToAlu_108, A0=>outFilter0(108), A1=>
      nx8614, B0=>outFilter1(108), B1=>nx8724);
   ix2213 : ao22 port map ( Y=>FilterToAlu_109, A0=>outFilter0(109), A1=>
      nx8614, B0=>outFilter1(109), B1=>nx8724);
   ix2219 : ao22 port map ( Y=>FilterToAlu_110, A0=>outFilter0(110), A1=>
      nx8614, B0=>outFilter1(110), B1=>nx8724);
   ix2225 : ao22 port map ( Y=>FilterToAlu_111, A0=>outFilter0(111), A1=>
      nx8614, B0=>outFilter1(111), B1=>nx8724);
   ix2051 : ao22 port map ( Y=>FilterToAlu_112, A0=>outFilter0(112), A1=>
      nx8616, B0=>outFilter1(112), B1=>nx8726);
   ix2057 : ao22 port map ( Y=>FilterToAlu_113, A0=>outFilter0(113), A1=>
      nx8616, B0=>outFilter1(113), B1=>nx8726);
   ix2063 : ao22 port map ( Y=>FilterToAlu_114, A0=>outFilter0(114), A1=>
      nx8616, B0=>outFilter1(114), B1=>nx8726);
   ix2069 : ao22 port map ( Y=>FilterToAlu_115, A0=>outFilter0(115), A1=>
      nx8616, B0=>outFilter1(115), B1=>nx8726);
   ix2075 : ao22 port map ( Y=>FilterToAlu_116, A0=>outFilter0(116), A1=>
      nx8616, B0=>outFilter1(116), B1=>nx8726);
   ix2081 : ao22 port map ( Y=>FilterToAlu_117, A0=>outFilter0(117), A1=>
      nx8616, B0=>outFilter1(117), B1=>nx8726);
   ix2087 : ao22 port map ( Y=>FilterToAlu_118, A0=>outFilter0(118), A1=>
      nx8616, B0=>outFilter1(118), B1=>nx8726);
   ix2093 : ao22 port map ( Y=>FilterToAlu_119, A0=>outFilter0(119), A1=>
      nx8618, B0=>outFilter1(119), B1=>nx8728);
   ix2099 : ao22 port map ( Y=>FilterToAlu_120, A0=>outFilter0(120), A1=>
      nx8618, B0=>outFilter1(120), B1=>nx8728);
   ix435 : nand02 port map ( Y=>FilterToAlu_121, A0=>nx8180, A1=>nx8806);
   ix8181 : mux21 port map ( Y=>nx8180, A0=>outFilter0(121), A1=>
      outFilter1(121), S0=>nx8898);
   ix2105 : ao22 port map ( Y=>FilterToAlu_122, A0=>outFilter0(122), A1=>
      nx8618, B0=>outFilter1(122), B1=>nx8728);
   ix2111 : ao22 port map ( Y=>FilterToAlu_123, A0=>outFilter0(123), A1=>
      nx8618, B0=>outFilter1(123), B1=>nx8728);
   ix2117 : ao22 port map ( Y=>FilterToAlu_124, A0=>outFilter0(124), A1=>
      nx8618, B0=>outFilter1(124), B1=>nx8728);
   ix2123 : ao22 port map ( Y=>FilterToAlu_125, A0=>outFilter0(125), A1=>
      nx8618, B0=>outFilter1(125), B1=>nx8728);
   ix2129 : ao22 port map ( Y=>FilterToAlu_126, A0=>outFilter0(126), A1=>
      nx8618, B0=>outFilter1(126), B1=>nx8728);
   ix2135 : ao22 port map ( Y=>FilterToAlu_127, A0=>outFilter0(127), A1=>
      nx8620, B0=>outFilter1(127), B1=>nx8730);
   ix1961 : ao22 port map ( Y=>FilterToAlu_128, A0=>outFilter0(128), A1=>
      nx8620, B0=>outFilter1(128), B1=>nx8730);
   ix1967 : ao22 port map ( Y=>FilterToAlu_129, A0=>outFilter0(129), A1=>
      nx8620, B0=>outFilter1(129), B1=>nx8730);
   ix1973 : ao22 port map ( Y=>FilterToAlu_130, A0=>outFilter0(130), A1=>
      nx8620, B0=>outFilter1(130), B1=>nx8730);
   ix1979 : ao22 port map ( Y=>FilterToAlu_131, A0=>outFilter0(131), A1=>
      nx8620, B0=>outFilter1(131), B1=>nx8730);
   ix1985 : ao22 port map ( Y=>FilterToAlu_132, A0=>outFilter0(132), A1=>
      nx8620, B0=>outFilter1(132), B1=>nx8730);
   ix1991 : ao22 port map ( Y=>FilterToAlu_133, A0=>outFilter0(133), A1=>
      nx8620, B0=>outFilter1(133), B1=>nx8730);
   ix1997 : ao22 port map ( Y=>FilterToAlu_134, A0=>outFilter0(134), A1=>
      nx8622, B0=>outFilter1(134), B1=>nx8732);
   ix2003 : ao22 port map ( Y=>FilterToAlu_135, A0=>outFilter0(135), A1=>
      nx8622, B0=>outFilter1(135), B1=>nx8732);
   ix2009 : ao22 port map ( Y=>FilterToAlu_136, A0=>outFilter0(136), A1=>
      nx8622, B0=>outFilter1(136), B1=>nx8732);
   ix425 : nand02 port map ( Y=>FilterToAlu_137, A0=>nx8198, A1=>nx8806);
   ix8199 : mux21 port map ( Y=>nx8198, A0=>outFilter0(137), A1=>
      outFilter1(137), S0=>nx8898);
   ix2015 : ao22 port map ( Y=>FilterToAlu_138, A0=>outFilter0(138), A1=>
      nx8622, B0=>outFilter1(138), B1=>nx8732);
   ix2021 : ao22 port map ( Y=>FilterToAlu_139, A0=>outFilter0(139), A1=>
      nx8622, B0=>outFilter1(139), B1=>nx8732);
   ix2027 : ao22 port map ( Y=>FilterToAlu_140, A0=>outFilter0(140), A1=>
      nx8622, B0=>outFilter1(140), B1=>nx8732);
   ix2033 : ao22 port map ( Y=>FilterToAlu_141, A0=>outFilter0(141), A1=>
      nx8622, B0=>outFilter1(141), B1=>nx8732);
   ix2039 : ao22 port map ( Y=>FilterToAlu_142, A0=>outFilter0(142), A1=>
      nx8624, B0=>outFilter1(142), B1=>nx8734);
   ix2045 : ao22 port map ( Y=>FilterToAlu_143, A0=>outFilter0(143), A1=>
      nx8624, B0=>outFilter1(143), B1=>nx8734);
   ix1871 : ao22 port map ( Y=>FilterToAlu_144, A0=>outFilter0(144), A1=>
      nx8624, B0=>outFilter1(144), B1=>nx8734);
   ix1877 : ao22 port map ( Y=>FilterToAlu_145, A0=>outFilter0(145), A1=>
      nx8624, B0=>outFilter1(145), B1=>nx8734);
   ix1883 : ao22 port map ( Y=>FilterToAlu_146, A0=>outFilter0(146), A1=>
      nx8624, B0=>outFilter1(146), B1=>nx8734);
   ix1889 : ao22 port map ( Y=>FilterToAlu_147, A0=>outFilter0(147), A1=>
      nx8624, B0=>outFilter1(147), B1=>nx8734);
   ix1895 : ao22 port map ( Y=>FilterToAlu_148, A0=>outFilter0(148), A1=>
      nx8624, B0=>outFilter1(148), B1=>nx8734);
   ix1901 : ao22 port map ( Y=>FilterToAlu_149, A0=>outFilter0(149), A1=>
      nx8626, B0=>outFilter1(149), B1=>nx8736);
   ix1907 : ao22 port map ( Y=>FilterToAlu_150, A0=>outFilter0(150), A1=>
      nx8626, B0=>outFilter1(150), B1=>nx8736);
   ix1913 : ao22 port map ( Y=>FilterToAlu_151, A0=>outFilter0(151), A1=>
      nx8626, B0=>outFilter1(151), B1=>nx8736);
   ix1919 : ao22 port map ( Y=>FilterToAlu_152, A0=>outFilter0(152), A1=>
      nx8626, B0=>outFilter1(152), B1=>nx8736);
   ix415 : nand02 port map ( Y=>FilterToAlu_153, A0=>nx8216, A1=>nx8806);
   ix8217 : mux21 port map ( Y=>nx8216, A0=>outFilter0(153), A1=>
      outFilter1(153), S0=>nx8898);
   ix1925 : ao22 port map ( Y=>FilterToAlu_154, A0=>outFilter0(154), A1=>
      nx8626, B0=>outFilter1(154), B1=>nx8736);
   ix1931 : ao22 port map ( Y=>FilterToAlu_155, A0=>outFilter0(155), A1=>
      nx8626, B0=>outFilter1(155), B1=>nx8736);
   ix1937 : ao22 port map ( Y=>FilterToAlu_156, A0=>outFilter0(156), A1=>
      nx8626, B0=>outFilter1(156), B1=>nx8736);
   ix1943 : ao22 port map ( Y=>FilterToAlu_157, A0=>outFilter0(157), A1=>
      nx8628, B0=>outFilter1(157), B1=>nx8738);
   ix1949 : ao22 port map ( Y=>FilterToAlu_158, A0=>outFilter0(158), A1=>
      nx8628, B0=>outFilter1(158), B1=>nx8738);
   ix1955 : ao22 port map ( Y=>FilterToAlu_159, A0=>outFilter0(159), A1=>
      nx8628, B0=>outFilter1(159), B1=>nx8738);
   ix1781 : ao22 port map ( Y=>FilterToAlu_160, A0=>outFilter0(160), A1=>
      nx8628, B0=>outFilter1(160), B1=>nx8738);
   ix1787 : ao22 port map ( Y=>FilterToAlu_161, A0=>outFilter0(161), A1=>
      nx8628, B0=>outFilter1(161), B1=>nx8738);
   ix1793 : ao22 port map ( Y=>FilterToAlu_162, A0=>outFilter0(162), A1=>
      nx8628, B0=>outFilter1(162), B1=>nx8738);
   ix1799 : ao22 port map ( Y=>FilterToAlu_163, A0=>outFilter0(163), A1=>
      nx8628, B0=>outFilter1(163), B1=>nx8738);
   ix1805 : ao22 port map ( Y=>FilterToAlu_164, A0=>outFilter0(164), A1=>
      nx8630, B0=>outFilter1(164), B1=>nx8740);
   ix1811 : ao22 port map ( Y=>FilterToAlu_165, A0=>outFilter0(165), A1=>
      nx8630, B0=>outFilter1(165), B1=>nx8740);
   ix1817 : ao22 port map ( Y=>FilterToAlu_166, A0=>outFilter0(166), A1=>
      nx8630, B0=>outFilter1(166), B1=>nx8740);
   ix1823 : ao22 port map ( Y=>FilterToAlu_167, A0=>outFilter0(167), A1=>
      nx8630, B0=>outFilter1(167), B1=>nx8740);
   ix1829 : ao22 port map ( Y=>FilterToAlu_168, A0=>outFilter0(168), A1=>
      nx8630, B0=>outFilter1(168), B1=>nx8740);
   ix405 : nand02 port map ( Y=>FilterToAlu_169, A0=>nx8234, A1=>nx8806);
   ix8235 : mux21 port map ( Y=>nx8234, A0=>outFilter0(169), A1=>
      outFilter1(169), S0=>nx8898);
   ix1835 : ao22 port map ( Y=>FilterToAlu_170, A0=>outFilter0(170), A1=>
      nx8630, B0=>outFilter1(170), B1=>nx8740);
   ix1841 : ao22 port map ( Y=>FilterToAlu_171, A0=>outFilter0(171), A1=>
      nx8630, B0=>outFilter1(171), B1=>nx8740);
   ix1847 : ao22 port map ( Y=>FilterToAlu_172, A0=>outFilter0(172), A1=>
      nx8632, B0=>outFilter1(172), B1=>nx8742);
   ix1853 : ao22 port map ( Y=>FilterToAlu_173, A0=>outFilter0(173), A1=>
      nx8632, B0=>outFilter1(173), B1=>nx8742);
   ix1859 : ao22 port map ( Y=>FilterToAlu_174, A0=>outFilter0(174), A1=>
      nx8632, B0=>outFilter1(174), B1=>nx8742);
   ix1865 : ao22 port map ( Y=>FilterToAlu_175, A0=>outFilter0(175), A1=>
      nx8632, B0=>outFilter1(175), B1=>nx8742);
   ix1691 : ao22 port map ( Y=>FilterToAlu_176, A0=>outFilter0(176), A1=>
      nx8632, B0=>outFilter1(176), B1=>nx8742);
   ix1697 : ao22 port map ( Y=>FilterToAlu_177, A0=>outFilter0(177), A1=>
      nx8632, B0=>outFilter1(177), B1=>nx8742);
   ix1703 : ao22 port map ( Y=>FilterToAlu_178, A0=>outFilter0(178), A1=>
      nx8632, B0=>outFilter1(178), B1=>nx8742);
   ix1709 : ao22 port map ( Y=>FilterToAlu_179, A0=>outFilter0(179), A1=>
      nx8634, B0=>outFilter1(179), B1=>nx8744);
   ix1715 : ao22 port map ( Y=>FilterToAlu_180, A0=>outFilter0(180), A1=>
      nx8634, B0=>outFilter1(180), B1=>nx8744);
   ix1721 : ao22 port map ( Y=>FilterToAlu_181, A0=>outFilter0(181), A1=>
      nx8634, B0=>outFilter1(181), B1=>nx8744);
   ix1727 : ao22 port map ( Y=>FilterToAlu_182, A0=>outFilter0(182), A1=>
      nx8634, B0=>outFilter1(182), B1=>nx8744);
   ix1733 : ao22 port map ( Y=>FilterToAlu_183, A0=>outFilter0(183), A1=>
      nx8634, B0=>outFilter1(183), B1=>nx8744);
   ix1739 : ao22 port map ( Y=>FilterToAlu_184, A0=>outFilter0(184), A1=>
      nx8634, B0=>outFilter1(184), B1=>nx8744);
   ix395 : nand02 port map ( Y=>FilterToAlu_185, A0=>nx8252, A1=>nx8806);
   ix8253 : mux21 port map ( Y=>nx8252, A0=>outFilter0(185), A1=>
      outFilter1(185), S0=>nx8898);
   ix1745 : ao22 port map ( Y=>FilterToAlu_186, A0=>outFilter0(186), A1=>
      nx8634, B0=>outFilter1(186), B1=>nx8744);
   ix1751 : ao22 port map ( Y=>FilterToAlu_187, A0=>outFilter0(187), A1=>
      nx8636, B0=>outFilter1(187), B1=>nx8746);
   ix1757 : ao22 port map ( Y=>FilterToAlu_188, A0=>outFilter0(188), A1=>
      nx8636, B0=>outFilter1(188), B1=>nx8746);
   ix1763 : ao22 port map ( Y=>FilterToAlu_189, A0=>outFilter0(189), A1=>
      nx8636, B0=>outFilter1(189), B1=>nx8746);
   ix1769 : ao22 port map ( Y=>FilterToAlu_190, A0=>outFilter0(190), A1=>
      nx8636, B0=>outFilter1(190), B1=>nx8746);
   ix1775 : ao22 port map ( Y=>FilterToAlu_191, A0=>outFilter0(191), A1=>
      nx8636, B0=>outFilter1(191), B1=>nx8746);
   ix1601 : ao22 port map ( Y=>FilterToAlu_192, A0=>outFilter0(192), A1=>
      nx8636, B0=>outFilter1(192), B1=>nx8746);
   ix1607 : ao22 port map ( Y=>FilterToAlu_193, A0=>outFilter0(193), A1=>
      nx8636, B0=>outFilter1(193), B1=>nx8746);
   ix1613 : ao22 port map ( Y=>FilterToAlu_194, A0=>outFilter0(194), A1=>
      nx8638, B0=>outFilter1(194), B1=>nx8748);
   ix1619 : ao22 port map ( Y=>FilterToAlu_195, A0=>outFilter0(195), A1=>
      nx8638, B0=>outFilter1(195), B1=>nx8748);
   ix1625 : ao22 port map ( Y=>FilterToAlu_196, A0=>outFilter0(196), A1=>
      nx8638, B0=>outFilter1(196), B1=>nx8748);
   ix1631 : ao22 port map ( Y=>FilterToAlu_197, A0=>outFilter0(197), A1=>
      nx8638, B0=>outFilter1(197), B1=>nx8748);
   ix1637 : ao22 port map ( Y=>FilterToAlu_198, A0=>outFilter0(198), A1=>
      nx8638, B0=>outFilter1(198), B1=>nx8748);
   ix1643 : ao22 port map ( Y=>FilterToAlu_199, A0=>outFilter0(199), A1=>
      nx8638, B0=>outFilter1(199), B1=>nx8748);
   ix1649 : ao22 port map ( Y=>FilterToAlu_200, A0=>outFilter0(200), A1=>
      nx8638, B0=>outFilter1(200), B1=>nx8748);
   ix385 : nand02 port map ( Y=>FilterToAlu_201, A0=>nx8270, A1=>nx8806);
   ix8271 : mux21 port map ( Y=>nx8270, A0=>outFilter0(201), A1=>
      outFilter1(201), S0=>nx8898);
   ix1655 : ao22 port map ( Y=>FilterToAlu_202, A0=>outFilter0(202), A1=>
      nx8640, B0=>outFilter1(202), B1=>nx8750);
   ix1661 : ao22 port map ( Y=>FilterToAlu_203, A0=>outFilter0(203), A1=>
      nx8640, B0=>outFilter1(203), B1=>nx8750);
   ix1667 : ao22 port map ( Y=>FilterToAlu_204, A0=>outFilter0(204), A1=>
      nx8640, B0=>outFilter1(204), B1=>nx8750);
   ix1673 : ao22 port map ( Y=>FilterToAlu_205, A0=>outFilter0(205), A1=>
      nx8640, B0=>outFilter1(205), B1=>nx8750);
   ix1679 : ao22 port map ( Y=>FilterToAlu_206, A0=>outFilter0(206), A1=>
      nx8640, B0=>outFilter1(206), B1=>nx8750);
   ix1685 : ao22 port map ( Y=>FilterToAlu_207, A0=>outFilter0(207), A1=>
      nx8640, B0=>outFilter1(207), B1=>nx8750);
   ix1511 : ao22 port map ( Y=>FilterToAlu_208, A0=>outFilter0(208), A1=>
      nx8640, B0=>outFilter1(208), B1=>nx8750);
   ix1517 : ao22 port map ( Y=>FilterToAlu_209, A0=>outFilter0(209), A1=>
      nx8642, B0=>outFilter1(209), B1=>nx8752);
   ix1523 : ao22 port map ( Y=>FilterToAlu_210, A0=>outFilter0(210), A1=>
      nx8642, B0=>outFilter1(210), B1=>nx8752);
   ix1529 : ao22 port map ( Y=>FilterToAlu_211, A0=>outFilter0(211), A1=>
      nx8642, B0=>outFilter1(211), B1=>nx8752);
   ix1535 : ao22 port map ( Y=>FilterToAlu_212, A0=>outFilter0(212), A1=>
      nx8642, B0=>outFilter1(212), B1=>nx8752);
   ix1541 : ao22 port map ( Y=>FilterToAlu_213, A0=>outFilter0(213), A1=>
      nx8642, B0=>outFilter1(213), B1=>nx8752);
   ix1547 : ao22 port map ( Y=>FilterToAlu_214, A0=>outFilter0(214), A1=>
      nx8642, B0=>outFilter1(214), B1=>nx8752);
   ix1553 : ao22 port map ( Y=>FilterToAlu_215, A0=>outFilter0(215), A1=>
      nx8642, B0=>outFilter1(215), B1=>nx8752);
   ix1559 : ao22 port map ( Y=>FilterToAlu_216, A0=>outFilter0(216), A1=>
      nx8644, B0=>outFilter1(216), B1=>nx8754);
   ix375 : nand02 port map ( Y=>FilterToAlu_217, A0=>nx8288, A1=>nx8806);
   ix8289 : mux21 port map ( Y=>nx8288, A0=>outFilter0(217), A1=>
      outFilter1(217), S0=>nx8900);
   ix1565 : ao22 port map ( Y=>FilterToAlu_218, A0=>outFilter0(218), A1=>
      nx8644, B0=>outFilter1(218), B1=>nx8754);
   ix1571 : ao22 port map ( Y=>FilterToAlu_219, A0=>outFilter0(219), A1=>
      nx8644, B0=>outFilter1(219), B1=>nx8754);
   ix1577 : ao22 port map ( Y=>FilterToAlu_220, A0=>outFilter0(220), A1=>
      nx8644, B0=>outFilter1(220), B1=>nx8754);
   ix1583 : ao22 port map ( Y=>FilterToAlu_221, A0=>outFilter0(221), A1=>
      nx8644, B0=>outFilter1(221), B1=>nx8754);
   ix1589 : ao22 port map ( Y=>FilterToAlu_222, A0=>outFilter0(222), A1=>
      nx8644, B0=>outFilter1(222), B1=>nx8754);
   ix1595 : ao22 port map ( Y=>FilterToAlu_223, A0=>outFilter0(223), A1=>
      nx8644, B0=>outFilter1(223), B1=>nx8754);
   ix1421 : ao22 port map ( Y=>FilterToAlu_224, A0=>outFilter0(224), A1=>
      nx8646, B0=>outFilter1(224), B1=>nx8756);
   ix1427 : ao22 port map ( Y=>FilterToAlu_225, A0=>outFilter0(225), A1=>
      nx8646, B0=>outFilter1(225), B1=>nx8756);
   ix1433 : ao22 port map ( Y=>FilterToAlu_226, A0=>outFilter0(226), A1=>
      nx8646, B0=>outFilter1(226), B1=>nx8756);
   ix1439 : ao22 port map ( Y=>FilterToAlu_227, A0=>outFilter0(227), A1=>
      nx8646, B0=>outFilter1(227), B1=>nx8756);
   ix1445 : ao22 port map ( Y=>FilterToAlu_228, A0=>outFilter0(228), A1=>
      nx8646, B0=>outFilter1(228), B1=>nx8756);
   ix1451 : ao22 port map ( Y=>FilterToAlu_229, A0=>outFilter0(229), A1=>
      nx8646, B0=>outFilter1(229), B1=>nx8756);
   ix1457 : ao22 port map ( Y=>FilterToAlu_230, A0=>outFilter0(230), A1=>
      nx8646, B0=>outFilter1(230), B1=>nx8756);
   ix1463 : ao22 port map ( Y=>FilterToAlu_231, A0=>outFilter0(231), A1=>
      nx8648, B0=>outFilter1(231), B1=>nx8758);
   ix1469 : ao22 port map ( Y=>FilterToAlu_232, A0=>outFilter0(232), A1=>
      nx8648, B0=>outFilter1(232), B1=>nx8758);
   ix365 : nand02 port map ( Y=>FilterToAlu_233, A0=>nx8306, A1=>nx8808);
   ix8307 : mux21 port map ( Y=>nx8306, A0=>outFilter0(233), A1=>
      outFilter1(233), S0=>nx8900);
   ix1475 : ao22 port map ( Y=>FilterToAlu_234, A0=>outFilter0(234), A1=>
      nx8648, B0=>outFilter1(234), B1=>nx8758);
   ix1481 : ao22 port map ( Y=>FilterToAlu_235, A0=>outFilter0(235), A1=>
      nx8648, B0=>outFilter1(235), B1=>nx8758);
   ix1487 : ao22 port map ( Y=>FilterToAlu_236, A0=>outFilter0(236), A1=>
      nx8648, B0=>outFilter1(236), B1=>nx8758);
   ix1493 : ao22 port map ( Y=>FilterToAlu_237, A0=>outFilter0(237), A1=>
      nx8648, B0=>outFilter1(237), B1=>nx8758);
   ix1499 : ao22 port map ( Y=>FilterToAlu_238, A0=>outFilter0(238), A1=>
      nx8648, B0=>outFilter1(238), B1=>nx8758);
   ix1505 : ao22 port map ( Y=>FilterToAlu_239, A0=>outFilter0(239), A1=>
      nx8650, B0=>outFilter1(239), B1=>nx8760);
   ix1331 : ao22 port map ( Y=>FilterToAlu_240, A0=>outFilter0(240), A1=>
      nx8650, B0=>outFilter1(240), B1=>nx8760);
   ix1337 : ao22 port map ( Y=>FilterToAlu_241, A0=>outFilter0(241), A1=>
      nx8650, B0=>outFilter1(241), B1=>nx8760);
   ix1343 : ao22 port map ( Y=>FilterToAlu_242, A0=>outFilter0(242), A1=>
      nx8650, B0=>outFilter1(242), B1=>nx8760);
   ix1349 : ao22 port map ( Y=>FilterToAlu_243, A0=>outFilter0(243), A1=>
      nx8650, B0=>outFilter1(243), B1=>nx8760);
   ix1355 : ao22 port map ( Y=>FilterToAlu_244, A0=>outFilter0(244), A1=>
      nx8650, B0=>outFilter1(244), B1=>nx8760);
   ix1361 : ao22 port map ( Y=>FilterToAlu_245, A0=>outFilter0(245), A1=>
      nx8650, B0=>outFilter1(245), B1=>nx8760);
   ix1367 : ao22 port map ( Y=>FilterToAlu_246, A0=>outFilter0(246), A1=>
      nx8652, B0=>outFilter1(246), B1=>nx8762);
   ix1373 : ao22 port map ( Y=>FilterToAlu_247, A0=>outFilter0(247), A1=>
      nx8652, B0=>outFilter1(247), B1=>nx8762);
   ix1379 : ao22 port map ( Y=>FilterToAlu_248, A0=>outFilter0(248), A1=>
      nx8652, B0=>outFilter1(248), B1=>nx8762);
   ix355 : nand02 port map ( Y=>FilterToAlu_249, A0=>nx8324, A1=>nx8808);
   ix8325 : mux21 port map ( Y=>nx8324, A0=>outFilter0(249), A1=>
      outFilter1(249), S0=>nx8900);
   ix1385 : ao22 port map ( Y=>FilterToAlu_250, A0=>outFilter0(250), A1=>
      nx8652, B0=>outFilter1(250), B1=>nx8762);
   ix1391 : ao22 port map ( Y=>FilterToAlu_251, A0=>outFilter0(251), A1=>
      nx8652, B0=>outFilter1(251), B1=>nx8762);
   ix1397 : ao22 port map ( Y=>FilterToAlu_252, A0=>outFilter0(252), A1=>
      nx8652, B0=>outFilter1(252), B1=>nx8762);
   ix1403 : ao22 port map ( Y=>FilterToAlu_253, A0=>outFilter0(253), A1=>
      nx8652, B0=>outFilter1(253), B1=>nx8762);
   ix1409 : ao22 port map ( Y=>FilterToAlu_254, A0=>outFilter0(254), A1=>
      nx8654, B0=>outFilter1(254), B1=>nx8764);
   ix1415 : ao22 port map ( Y=>FilterToAlu_255, A0=>outFilter0(255), A1=>
      nx8654, B0=>outFilter1(255), B1=>nx8764);
   ix1241 : ao22 port map ( Y=>FilterToAlu_256, A0=>outFilter0(256), A1=>
      nx8654, B0=>outFilter1(256), B1=>nx8764);
   ix1247 : ao22 port map ( Y=>FilterToAlu_257, A0=>outFilter0(257), A1=>
      nx8654, B0=>outFilter1(257), B1=>nx8764);
   ix1253 : ao22 port map ( Y=>FilterToAlu_258, A0=>outFilter0(258), A1=>
      nx8654, B0=>outFilter1(258), B1=>nx8764);
   ix1259 : ao22 port map ( Y=>FilterToAlu_259, A0=>outFilter0(259), A1=>
      nx8654, B0=>outFilter1(259), B1=>nx8764);
   ix1265 : ao22 port map ( Y=>FilterToAlu_260, A0=>outFilter0(260), A1=>
      nx8654, B0=>outFilter1(260), B1=>nx8764);
   ix1271 : ao22 port map ( Y=>FilterToAlu_261, A0=>outFilter0(261), A1=>
      nx8656, B0=>outFilter1(261), B1=>nx8766);
   ix1277 : ao22 port map ( Y=>FilterToAlu_262, A0=>outFilter0(262), A1=>
      nx8656, B0=>outFilter1(262), B1=>nx8766);
   ix1283 : ao22 port map ( Y=>FilterToAlu_263, A0=>outFilter0(263), A1=>
      nx8656, B0=>outFilter1(263), B1=>nx8766);
   ix1289 : ao22 port map ( Y=>FilterToAlu_264, A0=>outFilter0(264), A1=>
      nx8656, B0=>outFilter1(264), B1=>nx8766);
   ix345 : nand02 port map ( Y=>FilterToAlu_265, A0=>nx8342, A1=>nx8808);
   ix8343 : mux21 port map ( Y=>nx8342, A0=>outFilter0(265), A1=>
      outFilter1(265), S0=>nx8900);
   ix1295 : ao22 port map ( Y=>FilterToAlu_266, A0=>outFilter0(266), A1=>
      nx8656, B0=>outFilter1(266), B1=>nx8766);
   ix1301 : ao22 port map ( Y=>FilterToAlu_267, A0=>outFilter0(267), A1=>
      nx8656, B0=>outFilter1(267), B1=>nx8766);
   ix1307 : ao22 port map ( Y=>FilterToAlu_268, A0=>outFilter0(268), A1=>
      nx8656, B0=>outFilter1(268), B1=>nx8766);
   ix1313 : ao22 port map ( Y=>FilterToAlu_269, A0=>outFilter0(269), A1=>
      nx8658, B0=>outFilter1(269), B1=>nx8768);
   ix1319 : ao22 port map ( Y=>FilterToAlu_270, A0=>outFilter0(270), A1=>
      nx8658, B0=>outFilter1(270), B1=>nx8768);
   ix1325 : ao22 port map ( Y=>FilterToAlu_271, A0=>outFilter0(271), A1=>
      nx8658, B0=>outFilter1(271), B1=>nx8768);
   ix1151 : ao22 port map ( Y=>FilterToAlu_272, A0=>outFilter0(272), A1=>
      nx8658, B0=>outFilter1(272), B1=>nx8768);
   ix1157 : ao22 port map ( Y=>FilterToAlu_273, A0=>outFilter0(273), A1=>
      nx8658, B0=>outFilter1(273), B1=>nx8768);
   ix1163 : ao22 port map ( Y=>FilterToAlu_274, A0=>outFilter0(274), A1=>
      nx8658, B0=>outFilter1(274), B1=>nx8768);
   ix1169 : ao22 port map ( Y=>FilterToAlu_275, A0=>outFilter0(275), A1=>
      nx8658, B0=>outFilter1(275), B1=>nx8768);
   ix1175 : ao22 port map ( Y=>FilterToAlu_276, A0=>outFilter0(276), A1=>
      nx8660, B0=>outFilter1(276), B1=>nx8770);
   ix1181 : ao22 port map ( Y=>FilterToAlu_277, A0=>outFilter0(277), A1=>
      nx8660, B0=>outFilter1(277), B1=>nx8770);
   ix1187 : ao22 port map ( Y=>FilterToAlu_278, A0=>outFilter0(278), A1=>
      nx8660, B0=>outFilter1(278), B1=>nx8770);
   ix1193 : ao22 port map ( Y=>FilterToAlu_279, A0=>outFilter0(279), A1=>
      nx8660, B0=>outFilter1(279), B1=>nx8770);
   ix1199 : ao22 port map ( Y=>FilterToAlu_280, A0=>outFilter0(280), A1=>
      nx8660, B0=>outFilter1(280), B1=>nx8770);
   ix335 : nand02 port map ( Y=>FilterToAlu_281, A0=>nx8360, A1=>nx8808);
   ix8361 : mux21 port map ( Y=>nx8360, A0=>outFilter0(281), A1=>
      outFilter1(281), S0=>nx8900);
   ix1205 : ao22 port map ( Y=>FilterToAlu_282, A0=>outFilter0(282), A1=>
      nx8660, B0=>outFilter1(282), B1=>nx8770);
   ix1211 : ao22 port map ( Y=>FilterToAlu_283, A0=>outFilter0(283), A1=>
      nx8660, B0=>outFilter1(283), B1=>nx8770);
   ix1217 : ao22 port map ( Y=>FilterToAlu_284, A0=>outFilter0(284), A1=>
      nx8662, B0=>outFilter1(284), B1=>nx8772);
   ix1223 : ao22 port map ( Y=>FilterToAlu_285, A0=>outFilter0(285), A1=>
      nx8662, B0=>outFilter1(285), B1=>nx8772);
   ix1229 : ao22 port map ( Y=>FilterToAlu_286, A0=>outFilter0(286), A1=>
      nx8662, B0=>outFilter1(286), B1=>nx8772);
   ix1235 : ao22 port map ( Y=>FilterToAlu_287, A0=>outFilter0(287), A1=>
      nx8662, B0=>outFilter1(287), B1=>nx8772);
   ix1061 : ao22 port map ( Y=>FilterToAlu_288, A0=>outFilter0(288), A1=>
      nx8662, B0=>outFilter1(288), B1=>nx8772);
   ix1067 : ao22 port map ( Y=>FilterToAlu_289, A0=>outFilter0(289), A1=>
      nx8662, B0=>outFilter1(289), B1=>nx8772);
   ix1073 : ao22 port map ( Y=>FilterToAlu_290, A0=>outFilter0(290), A1=>
      nx8662, B0=>outFilter1(290), B1=>nx8772);
   ix1079 : ao22 port map ( Y=>FilterToAlu_291, A0=>outFilter0(291), A1=>
      nx8664, B0=>outFilter1(291), B1=>nx8774);
   ix1085 : ao22 port map ( Y=>FilterToAlu_292, A0=>outFilter0(292), A1=>
      nx8664, B0=>outFilter1(292), B1=>nx8774);
   ix1091 : ao22 port map ( Y=>FilterToAlu_293, A0=>outFilter0(293), A1=>
      nx8664, B0=>outFilter1(293), B1=>nx8774);
   ix1097 : ao22 port map ( Y=>FilterToAlu_294, A0=>outFilter0(294), A1=>
      nx8664, B0=>outFilter1(294), B1=>nx8774);
   ix1103 : ao22 port map ( Y=>FilterToAlu_295, A0=>outFilter0(295), A1=>
      nx8664, B0=>outFilter1(295), B1=>nx8774);
   ix1109 : ao22 port map ( Y=>FilterToAlu_296, A0=>outFilter0(296), A1=>
      nx8664, B0=>outFilter1(296), B1=>nx8774);
   ix325 : nand02 port map ( Y=>FilterToAlu_297, A0=>nx8378, A1=>nx8808);
   ix8379 : mux21 port map ( Y=>nx8378, A0=>outFilter0(297), A1=>
      outFilter1(297), S0=>nx8900);
   ix1115 : ao22 port map ( Y=>FilterToAlu_298, A0=>outFilter0(298), A1=>
      nx8664, B0=>outFilter1(298), B1=>nx8774);
   ix1121 : ao22 port map ( Y=>FilterToAlu_299, A0=>outFilter0(299), A1=>
      nx8666, B0=>outFilter1(299), B1=>nx8776);
   ix1127 : ao22 port map ( Y=>FilterToAlu_300, A0=>outFilter0(300), A1=>
      nx8666, B0=>outFilter1(300), B1=>nx8776);
   ix1133 : ao22 port map ( Y=>FilterToAlu_301, A0=>outFilter0(301), A1=>
      nx8666, B0=>outFilter1(301), B1=>nx8776);
   ix1139 : ao22 port map ( Y=>FilterToAlu_302, A0=>outFilter0(302), A1=>
      nx8666, B0=>outFilter1(302), B1=>nx8776);
   ix1145 : ao22 port map ( Y=>FilterToAlu_303, A0=>outFilter0(303), A1=>
      nx8666, B0=>outFilter1(303), B1=>nx8776);
   ix971 : ao22 port map ( Y=>FilterToAlu_304, A0=>outFilter0(304), A1=>
      nx8666, B0=>outFilter1(304), B1=>nx8776);
   ix977 : ao22 port map ( Y=>FilterToAlu_305, A0=>outFilter0(305), A1=>
      nx8666, B0=>outFilter1(305), B1=>nx8776);
   ix983 : ao22 port map ( Y=>FilterToAlu_306, A0=>outFilter0(306), A1=>
      nx8668, B0=>outFilter1(306), B1=>nx8778);
   ix989 : ao22 port map ( Y=>FilterToAlu_307, A0=>outFilter0(307), A1=>
      nx8668, B0=>outFilter1(307), B1=>nx8778);
   ix995 : ao22 port map ( Y=>FilterToAlu_308, A0=>outFilter0(308), A1=>
      nx8668, B0=>outFilter1(308), B1=>nx8778);
   ix1001 : ao22 port map ( Y=>FilterToAlu_309, A0=>outFilter0(309), A1=>
      nx8668, B0=>outFilter1(309), B1=>nx8778);
   ix1007 : ao22 port map ( Y=>FilterToAlu_310, A0=>outFilter0(310), A1=>
      nx8668, B0=>outFilter1(310), B1=>nx8778);
   ix1013 : ao22 port map ( Y=>FilterToAlu_311, A0=>outFilter0(311), A1=>
      nx8668, B0=>outFilter1(311), B1=>nx8778);
   ix1019 : ao22 port map ( Y=>FilterToAlu_312, A0=>outFilter0(312), A1=>
      nx8668, B0=>outFilter1(312), B1=>nx8778);
   ix315 : nand02 port map ( Y=>FilterToAlu_313, A0=>nx8396, A1=>nx8808);
   ix8397 : mux21 port map ( Y=>nx8396, A0=>outFilter0(313), A1=>
      outFilter1(313), S0=>nx8900);
   ix1025 : ao22 port map ( Y=>FilterToAlu_314, A0=>outFilter0(314), A1=>
      nx8670, B0=>outFilter1(314), B1=>nx8780);
   ix1031 : ao22 port map ( Y=>FilterToAlu_315, A0=>outFilter0(315), A1=>
      nx8670, B0=>outFilter1(315), B1=>nx8780);
   ix1037 : ao22 port map ( Y=>FilterToAlu_316, A0=>outFilter0(316), A1=>
      nx8670, B0=>outFilter1(316), B1=>nx8780);
   ix1043 : ao22 port map ( Y=>FilterToAlu_317, A0=>outFilter0(317), A1=>
      nx8670, B0=>outFilter1(317), B1=>nx8780);
   ix1049 : ao22 port map ( Y=>FilterToAlu_318, A0=>outFilter0(318), A1=>
      nx8670, B0=>outFilter1(318), B1=>nx8780);
   ix1055 : ao22 port map ( Y=>FilterToAlu_319, A0=>outFilter0(319), A1=>
      nx8670, B0=>outFilter1(319), B1=>nx8780);
   ix881 : ao22 port map ( Y=>FilterToAlu_320, A0=>outFilter0(320), A1=>
      nx8670, B0=>outFilter1(320), B1=>nx8780);
   ix887 : ao22 port map ( Y=>FilterToAlu_321, A0=>outFilter0(321), A1=>
      nx8672, B0=>outFilter1(321), B1=>nx8782);
   ix893 : ao22 port map ( Y=>FilterToAlu_322, A0=>outFilter0(322), A1=>
      nx8672, B0=>outFilter1(322), B1=>nx8782);
   ix899 : ao22 port map ( Y=>FilterToAlu_323, A0=>outFilter0(323), A1=>
      nx8672, B0=>outFilter1(323), B1=>nx8782);
   ix905 : ao22 port map ( Y=>FilterToAlu_324, A0=>outFilter0(324), A1=>
      nx8672, B0=>outFilter1(324), B1=>nx8782);
   ix911 : ao22 port map ( Y=>FilterToAlu_325, A0=>outFilter0(325), A1=>
      nx8672, B0=>outFilter1(325), B1=>nx8782);
   ix917 : ao22 port map ( Y=>FilterToAlu_326, A0=>outFilter0(326), A1=>
      nx8672, B0=>outFilter1(326), B1=>nx8782);
   ix923 : ao22 port map ( Y=>FilterToAlu_327, A0=>outFilter0(327), A1=>
      nx8672, B0=>outFilter1(327), B1=>nx8782);
   ix929 : ao22 port map ( Y=>FilterToAlu_328, A0=>outFilter0(328), A1=>
      nx8674, B0=>outFilter1(328), B1=>nx8784);
   ix305 : nand02 port map ( Y=>FilterToAlu_329, A0=>nx8414, A1=>nx8808);
   ix8415 : mux21 port map ( Y=>nx8414, A0=>outFilter0(329), A1=>
      outFilter1(329), S0=>nx8902);
   ix935 : ao22 port map ( Y=>FilterToAlu_330, A0=>outFilter0(330), A1=>
      nx8674, B0=>outFilter1(330), B1=>nx8784);
   ix941 : ao22 port map ( Y=>FilterToAlu_331, A0=>outFilter0(331), A1=>
      nx8674, B0=>outFilter1(331), B1=>nx8784);
   ix947 : ao22 port map ( Y=>FilterToAlu_332, A0=>outFilter0(332), A1=>
      nx8674, B0=>outFilter1(332), B1=>nx8784);
   ix953 : ao22 port map ( Y=>FilterToAlu_333, A0=>outFilter0(333), A1=>
      nx8674, B0=>outFilter1(333), B1=>nx8784);
   ix959 : ao22 port map ( Y=>FilterToAlu_334, A0=>outFilter0(334), A1=>
      nx8674, B0=>outFilter1(334), B1=>nx8784);
   ix965 : ao22 port map ( Y=>FilterToAlu_335, A0=>outFilter0(335), A1=>
      nx8674, B0=>outFilter1(335), B1=>nx8784);
   ix791 : ao22 port map ( Y=>FilterToAlu_336, A0=>outFilter0(336), A1=>
      nx8676, B0=>outFilter1(336), B1=>nx8786);
   ix797 : ao22 port map ( Y=>FilterToAlu_337, A0=>outFilter0(337), A1=>
      nx8676, B0=>outFilter1(337), B1=>nx8786);
   ix803 : ao22 port map ( Y=>FilterToAlu_338, A0=>outFilter0(338), A1=>
      nx8676, B0=>outFilter1(338), B1=>nx8786);
   ix809 : ao22 port map ( Y=>FilterToAlu_339, A0=>outFilter0(339), A1=>
      nx8676, B0=>outFilter1(339), B1=>nx8786);
   ix815 : ao22 port map ( Y=>FilterToAlu_340, A0=>outFilter0(340), A1=>
      nx8676, B0=>outFilter1(340), B1=>nx8786);
   ix821 : ao22 port map ( Y=>FilterToAlu_341, A0=>outFilter0(341), A1=>
      nx8676, B0=>outFilter1(341), B1=>nx8786);
   ix827 : ao22 port map ( Y=>FilterToAlu_342, A0=>outFilter0(342), A1=>
      nx8676, B0=>outFilter1(342), B1=>nx8786);
   ix833 : ao22 port map ( Y=>FilterToAlu_343, A0=>outFilter0(343), A1=>
      nx8678, B0=>outFilter1(343), B1=>nx8788);
   ix839 : ao22 port map ( Y=>FilterToAlu_344, A0=>outFilter0(344), A1=>
      nx8678, B0=>outFilter1(344), B1=>nx8788);
   ix295 : nand02 port map ( Y=>FilterToAlu_345, A0=>nx8432, A1=>nx8810);
   ix8433 : mux21 port map ( Y=>nx8432, A0=>outFilter0(345), A1=>
      outFilter1(345), S0=>nx8902);
   ix845 : ao22 port map ( Y=>FilterToAlu_346, A0=>outFilter0(346), A1=>
      nx8678, B0=>outFilter1(346), B1=>nx8788);
   ix851 : ao22 port map ( Y=>FilterToAlu_347, A0=>outFilter0(347), A1=>
      nx8678, B0=>outFilter1(347), B1=>nx8788);
   ix857 : ao22 port map ( Y=>FilterToAlu_348, A0=>outFilter0(348), A1=>
      nx8678, B0=>outFilter1(348), B1=>nx8788);
   ix863 : ao22 port map ( Y=>FilterToAlu_349, A0=>outFilter0(349), A1=>
      nx8678, B0=>outFilter1(349), B1=>nx8788);
   ix869 : ao22 port map ( Y=>FilterToAlu_350, A0=>outFilter0(350), A1=>
      nx8678, B0=>outFilter1(350), B1=>nx8788);
   ix875 : ao22 port map ( Y=>FilterToAlu_351, A0=>outFilter0(351), A1=>
      nx8680, B0=>outFilter1(351), B1=>nx8790);
   ix701 : ao22 port map ( Y=>FilterToAlu_352, A0=>outFilter0(352), A1=>
      nx8680, B0=>outFilter1(352), B1=>nx8790);
   ix707 : ao22 port map ( Y=>FilterToAlu_353, A0=>outFilter0(353), A1=>
      nx8680, B0=>outFilter1(353), B1=>nx8790);
   ix713 : ao22 port map ( Y=>FilterToAlu_354, A0=>outFilter0(354), A1=>
      nx8680, B0=>outFilter1(354), B1=>nx8790);
   ix719 : ao22 port map ( Y=>FilterToAlu_355, A0=>outFilter0(355), A1=>
      nx8680, B0=>outFilter1(355), B1=>nx8790);
   ix725 : ao22 port map ( Y=>FilterToAlu_356, A0=>outFilter0(356), A1=>
      nx8680, B0=>outFilter1(356), B1=>nx8790);
   ix731 : ao22 port map ( Y=>FilterToAlu_357, A0=>outFilter0(357), A1=>
      nx8680, B0=>outFilter1(357), B1=>nx8790);
   ix737 : ao22 port map ( Y=>FilterToAlu_358, A0=>outFilter0(358), A1=>
      nx8682, B0=>outFilter1(358), B1=>nx8792);
   ix743 : ao22 port map ( Y=>FilterToAlu_359, A0=>outFilter0(359), A1=>
      nx8682, B0=>outFilter1(359), B1=>nx8792);
   ix749 : ao22 port map ( Y=>FilterToAlu_360, A0=>outFilter0(360), A1=>
      nx8682, B0=>outFilter1(360), B1=>nx8792);
   ix285 : nand02 port map ( Y=>FilterToAlu_361, A0=>nx8450, A1=>nx8810);
   ix8451 : mux21 port map ( Y=>nx8450, A0=>outFilter0(361), A1=>
      outFilter1(361), S0=>nx8902);
   ix755 : ao22 port map ( Y=>FilterToAlu_362, A0=>outFilter0(362), A1=>
      nx8682, B0=>outFilter1(362), B1=>nx8792);
   ix761 : ao22 port map ( Y=>FilterToAlu_363, A0=>outFilter0(363), A1=>
      nx8682, B0=>outFilter1(363), B1=>nx8792);
   ix767 : ao22 port map ( Y=>FilterToAlu_364, A0=>outFilter0(364), A1=>
      nx8682, B0=>outFilter1(364), B1=>nx8792);
   ix773 : ao22 port map ( Y=>FilterToAlu_365, A0=>outFilter0(365), A1=>
      nx8682, B0=>outFilter1(365), B1=>nx8792);
   ix779 : ao22 port map ( Y=>FilterToAlu_366, A0=>outFilter0(366), A1=>
      nx8684, B0=>outFilter1(366), B1=>nx8794);
   ix785 : ao22 port map ( Y=>FilterToAlu_367, A0=>outFilter0(367), A1=>
      nx8684, B0=>outFilter1(367), B1=>nx8794);
   ix611 : ao22 port map ( Y=>FilterToAlu_368, A0=>outFilter0(368), A1=>
      nx8684, B0=>outFilter1(368), B1=>nx8794);
   ix617 : ao22 port map ( Y=>FilterToAlu_369, A0=>outFilter0(369), A1=>
      nx8684, B0=>outFilter1(369), B1=>nx8794);
   ix623 : ao22 port map ( Y=>FilterToAlu_370, A0=>outFilter0(370), A1=>
      nx8684, B0=>outFilter1(370), B1=>nx8794);
   ix629 : ao22 port map ( Y=>FilterToAlu_371, A0=>outFilter0(371), A1=>
      nx8684, B0=>outFilter1(371), B1=>nx8794);
   ix635 : ao22 port map ( Y=>FilterToAlu_372, A0=>outFilter0(372), A1=>
      nx8684, B0=>outFilter1(372), B1=>nx8794);
   ix641 : ao22 port map ( Y=>FilterToAlu_373, A0=>outFilter0(373), A1=>
      nx8686, B0=>outFilter1(373), B1=>nx8796);
   ix647 : ao22 port map ( Y=>FilterToAlu_374, A0=>outFilter0(374), A1=>
      nx8686, B0=>outFilter1(374), B1=>nx8796);
   ix653 : ao22 port map ( Y=>FilterToAlu_375, A0=>outFilter0(375), A1=>
      nx8686, B0=>outFilter1(375), B1=>nx8796);
   ix659 : ao22 port map ( Y=>FilterToAlu_376, A0=>outFilter0(376), A1=>
      nx8686, B0=>outFilter1(376), B1=>nx8796);
   ix275 : nand02 port map ( Y=>FilterToAlu_377, A0=>nx8468, A1=>nx8810);
   ix8469 : mux21 port map ( Y=>nx8468, A0=>outFilter0(377), A1=>
      outFilter1(377), S0=>nx8902);
   ix665 : ao22 port map ( Y=>FilterToAlu_378, A0=>outFilter0(378), A1=>
      nx8686, B0=>outFilter1(378), B1=>nx8796);
   ix671 : ao22 port map ( Y=>FilterToAlu_379, A0=>outFilter0(379), A1=>
      nx8686, B0=>outFilter1(379), B1=>nx8796);
   ix677 : ao22 port map ( Y=>FilterToAlu_380, A0=>outFilter0(380), A1=>
      nx8686, B0=>outFilter1(380), B1=>nx8796);
   ix683 : ao22 port map ( Y=>FilterToAlu_381, A0=>outFilter0(381), A1=>
      nx8688, B0=>outFilter1(381), B1=>nx8798);
   ix689 : ao22 port map ( Y=>FilterToAlu_382, A0=>outFilter0(382), A1=>
      nx8688, B0=>outFilter1(382), B1=>nx8798);
   ix695 : ao22 port map ( Y=>FilterToAlu_383, A0=>outFilter0(383), A1=>
      nx8688, B0=>outFilter1(383), B1=>nx8798);
   ix521 : ao22 port map ( Y=>FilterToAlu_384, A0=>outFilter0(384), A1=>
      nx8688, B0=>outFilter1(384), B1=>nx8798);
   ix527 : ao22 port map ( Y=>FilterToAlu_385, A0=>outFilter0(385), A1=>
      nx8688, B0=>outFilter1(385), B1=>nx8798);
   ix533 : ao22 port map ( Y=>FilterToAlu_386, A0=>outFilter0(386), A1=>
      nx8688, B0=>outFilter1(386), B1=>nx8798);
   ix539 : ao22 port map ( Y=>FilterToAlu_387, A0=>outFilter0(387), A1=>
      nx8688, B0=>outFilter1(387), B1=>nx8798);
   ix545 : ao22 port map ( Y=>FilterToAlu_388, A0=>outFilter0(388), A1=>
      nx8690, B0=>outFilter1(388), B1=>nx8800);
   ix551 : ao22 port map ( Y=>FilterToAlu_389, A0=>outFilter0(389), A1=>
      nx8690, B0=>outFilter1(389), B1=>nx8800);
   ix557 : ao22 port map ( Y=>FilterToAlu_390, A0=>outFilter0(390), A1=>
      nx8690, B0=>outFilter1(390), B1=>nx8800);
   ix563 : ao22 port map ( Y=>FilterToAlu_391, A0=>outFilter0(391), A1=>
      nx8690, B0=>outFilter1(391), B1=>nx8800);
   ix569 : ao22 port map ( Y=>FilterToAlu_392, A0=>outFilter0(392), A1=>
      nx8690, B0=>outFilter1(392), B1=>nx8800);
   ix265 : nand02 port map ( Y=>FilterToAlu_393, A0=>nx8486, A1=>nx8810);
   ix8487 : mux21 port map ( Y=>nx8486, A0=>outFilter0(393), A1=>
      outFilter1(393), S0=>nx8902);
   ix575 : ao22 port map ( Y=>FilterToAlu_394, A0=>outFilter0(394), A1=>
      nx8690, B0=>outFilter1(394), B1=>nx8800);
   ix581 : ao22 port map ( Y=>FilterToAlu_395, A0=>outFilter0(395), A1=>
      nx8690, B0=>outFilter1(395), B1=>nx8800);
   ix587 : ao22 port map ( Y=>FilterToAlu_396, A0=>outFilter0(396), A1=>
      nx8692, B0=>outFilter1(396), B1=>nx8802);
   ix593 : ao22 port map ( Y=>FilterToAlu_397, A0=>outFilter0(397), A1=>
      nx8692, B0=>outFilter1(397), B1=>nx8802);
   ix599 : ao22 port map ( Y=>FilterToAlu_398, A0=>outFilter0(398), A1=>
      nx8692, B0=>outFilter1(398), B1=>nx8802);
   ix605 : ao22 port map ( Y=>FilterToAlu_399, A0=>outFilter0(399), A1=>
      nx8692, B0=>outFilter1(399), B1=>nx8802);
   ix55 : nand02 port map ( Y=>ConvOuput(0), A0=>nx8495, A1=>nx8501);
   ix8496 : aoi32 port map ( Y=>nx8495, A0=>nx8916, A1=>AddOut33_3, A2=>
      nx8852, B0=>nx32, B1=>nx34);
   ix33 : mux21_ni port map ( Y=>nx32, A0=>AddOut33_5, A1=>Final55_5, S0=>
      nx8884);
   ix8502 : aoi32 port map ( Y=>nx8501, A0=>Final55_0, A1=>nx8884, A2=>
      nx8904, B0=>AddOut33_0, B1=>nx20);
   ix13 : nor02_2x port map ( Y=>nx12, A0=>nx8852, A1=>nx6);
   ix7 : mux21_ni port map ( Y=>nx6, A0=>AddOut33_15, A1=>Final55_15, S0=>
      nx8886);
   ix85 : nand02 port map ( Y=>ConvOuput(1), A0=>nx8511, A1=>nx8514);
   ix8512 : aoi32 port map ( Y=>nx8511, A0=>nx8916, A1=>AddOut33_4, A2=>
      nx8852, B0=>nx68, B1=>nx34);
   ix69 : mux21_ni port map ( Y=>nx68, A0=>AddOut33_6, A1=>Final55_6, S0=>
      nx8886);
   ix8515 : aoi32 port map ( Y=>nx8514, A0=>Final55_1, A1=>nx8886, A2=>
      nx8904, B0=>AddOut33_1, B1=>nx20);
   ix107 : nand02 port map ( Y=>ConvOuput(2), A0=>nx8517, A1=>nx8520);
   ix8518 : aoi32 port map ( Y=>nx8517, A0=>Final55_7, A1=>nx8886, A2=>
      nx8852, B0=>nx32, B1=>nx8908);
   ix8521 : aoi32 port map ( Y=>nx8520, A0=>Final55_2, A1=>nx8886, A2=>
      nx8904, B0=>AddOut33_2, B1=>nx20);
   ix125 : oai21 port map ( Y=>ConvOuput(3), A0=>nx8523, A1=>nx8812, B0=>
      nx8525);
   ix8524 : mux21 port map ( Y=>nx8523, A0=>AddOut33_3, A1=>Final55_3, S0=>
      nx8886);
   ix8526 : aoi32 port map ( Y=>nx8525, A0=>Final55_8, A1=>nx8886, A2=>
      nx8852, B0=>nx68, B1=>nx8908);
   ix143 : oai21 port map ( Y=>ConvOuput(4), A0=>nx8528, A1=>nx8812, B0=>
      nx8530);
   ix8529 : mux21 port map ( Y=>nx8528, A0=>AddOut33_4, A1=>Final55_4, S0=>
      nx8888);
   ix8531 : aoi32 port map ( Y=>nx8530, A0=>Final55_9, A1=>nx8888, A2=>
      nx8852, B0=>nx98, B1=>nx8908);
   ix99 : mux21_ni port map ( Y=>nx98, A0=>AddOut33_7, A1=>Final55_7, S0=>
      nx8888);
   ix161 : oai21 port map ( Y=>ConvOuput(5), A0=>nx8534, A1=>nx8812, B0=>
      nx8536);
   ix8537 : aoi32 port map ( Y=>nx8536, A0=>Final55_10, A1=>nx8888, A2=>
      nx8854, B0=>nx116, B1=>nx8908);
   ix117 : mux21_ni port map ( Y=>nx116, A0=>AddOut33_8, A1=>Final55_8, S0=>
      nx8888);
   ix179 : oai21 port map ( Y=>ConvOuput(6), A0=>nx8540, A1=>nx8812, B0=>
      nx8542);
   ix8543 : aoi32 port map ( Y=>nx8542, A0=>Final55_11, A1=>nx8888, A2=>
      nx8854, B0=>nx134, B1=>nx8908);
   ix135 : mux21_ni port map ( Y=>nx134, A0=>AddOut33_9, A1=>Final55_9, S0=>
      nx8888);
   ix197 : oai21 port map ( Y=>ConvOuput(7), A0=>nx8546, A1=>nx8812, B0=>
      nx8548);
   ix8549 : aoi32 port map ( Y=>nx8548, A0=>Final55_12, A1=>nx8890, A2=>
      nx8854, B0=>nx152, B1=>nx8908);
   ix153 : mux21_ni port map ( Y=>nx152, A0=>AddOut33_10, A1=>Final55_10, S0
      =>nx8890);
   ix215 : oai21 port map ( Y=>ConvOuput(8), A0=>nx8552, A1=>nx8812, B0=>
      nx8554);
   ix8555 : aoi32 port map ( Y=>nx8554, A0=>Final55_13, A1=>nx8890, A2=>
      nx8854, B0=>nx170, B1=>nx8908);
   ix171 : mux21_ni port map ( Y=>nx170, A0=>AddOut33_11, A1=>Final55_11, S0
      =>nx8890);
   ix233 : oai21 port map ( Y=>ConvOuput(9), A0=>nx8558, A1=>nx8814, B0=>
      nx8560);
   ix8561 : aoi32 port map ( Y=>nx8560, A0=>Final55_14, A1=>nx8890, A2=>
      nx8854, B0=>nx188, B1=>nx8910);
   ix189 : mux21_ni port map ( Y=>nx188, A0=>AddOut33_12, A1=>Final55_12, S0
      =>nx8890);
   ix243 : oai21 port map ( Y=>ConvOuput(10), A0=>nx8564, A1=>nx8814, B0=>
      nx8566);
   ix8567 : aoi32 port map ( Y=>nx8566, A0=>nx8916, A1=>AddOut33_13, A2=>
      nx8854, B0=>nx6, B1=>nx34);
   ix253 : oai21 port map ( Y=>ConvOuput(11), A0=>nx8569, A1=>nx8814, B0=>
      nx8571);
   ix8572 : aoi32 port map ( Y=>nx8571, A0=>nx8916, A1=>AddOut33_14, A2=>
      nx8854, B0=>nx6, B1=>nx34);
   ix2769 : ao21 port map ( Y=>ConvOuput(12), A0=>nx188, A1=>nx8904, B0=>
      ConvOuput_15_EXMPLR);
   ix2773 : ao21 port map ( Y=>ConvOuput(13), A0=>nx206, A1=>nx8904, B0=>
      ConvOuput_15_EXMPLR);
   ix207 : mux21_ni port map ( Y=>nx206, A0=>AddOut33_13, A1=>Final55_13, S0
      =>nx8890);
   ix2777 : ao21 port map ( Y=>ConvOuput(14), A0=>nx224, A1=>nx8904, B0=>
      ConvOuput_15_EXMPLR);
   ix225 : mux21_ni port map ( Y=>nx224, A0=>AddOut33_14, A1=>Final55_14, S0
      =>nx8892);
   ix8570 : inv01 port map ( Y=>nx8569, A=>nx170);
   ix8565 : inv01 port map ( Y=>nx8564, A=>nx152);
   ix8559 : inv01 port map ( Y=>nx8558, A=>nx134);
   ix8553 : inv01 port map ( Y=>nx8552, A=>nx116);
   ix8547 : inv01 port map ( Y=>nx8546, A=>nx98);
   ix8541 : inv01 port map ( Y=>nx8540, A=>nx68);
   ix8535 : inv01 port map ( Y=>nx8534, A=>nx32);
   ix8585 : inv02 port map ( Y=>nx8586, A=>nx8816);
   ix8587 : inv02 port map ( Y=>nx8588, A=>nx8816);
   ix8589 : inv02 port map ( Y=>nx8590, A=>nx8816);
   ix8591 : inv02 port map ( Y=>nx8592, A=>nx8816);
   ix8593 : inv02 port map ( Y=>nx8594, A=>nx8816);
   ix8595 : inv02 port map ( Y=>nx8596, A=>nx8816);
   ix8597 : inv02 port map ( Y=>nx8598, A=>nx8816);
   ix8599 : inv02 port map ( Y=>nx8600, A=>nx8818);
   ix8601 : inv02 port map ( Y=>nx8602, A=>nx8818);
   ix8603 : inv02 port map ( Y=>nx8604, A=>nx8818);
   ix8605 : inv02 port map ( Y=>nx8606, A=>nx8818);
   ix8607 : inv02 port map ( Y=>nx8608, A=>nx8818);
   ix8609 : inv02 port map ( Y=>nx8610, A=>nx8818);
   ix8611 : inv02 port map ( Y=>nx8612, A=>nx8818);
   ix8613 : inv02 port map ( Y=>nx8614, A=>nx8820);
   ix8615 : inv02 port map ( Y=>nx8616, A=>nx8820);
   ix8617 : inv02 port map ( Y=>nx8618, A=>nx8820);
   ix8619 : inv02 port map ( Y=>nx8620, A=>nx8820);
   ix8621 : inv02 port map ( Y=>nx8622, A=>nx8820);
   ix8623 : inv02 port map ( Y=>nx8624, A=>nx8820);
   ix8625 : inv02 port map ( Y=>nx8626, A=>nx8820);
   ix8627 : inv02 port map ( Y=>nx8628, A=>nx8822);
   ix8629 : inv02 port map ( Y=>nx8630, A=>nx8822);
   ix8631 : inv02 port map ( Y=>nx8632, A=>nx8822);
   ix8633 : inv02 port map ( Y=>nx8634, A=>nx8822);
   ix8635 : inv02 port map ( Y=>nx8636, A=>nx8822);
   ix8637 : inv02 port map ( Y=>nx8638, A=>nx8822);
   ix8639 : inv02 port map ( Y=>nx8640, A=>nx8822);
   ix8641 : inv02 port map ( Y=>nx8642, A=>nx8824);
   ix8643 : inv02 port map ( Y=>nx8644, A=>nx8824);
   ix8645 : inv02 port map ( Y=>nx8646, A=>nx8824);
   ix8647 : inv02 port map ( Y=>nx8648, A=>nx8824);
   ix8649 : inv02 port map ( Y=>nx8650, A=>nx8824);
   ix8651 : inv02 port map ( Y=>nx8652, A=>nx8824);
   ix8653 : inv02 port map ( Y=>nx8654, A=>nx8824);
   ix8655 : inv02 port map ( Y=>nx8656, A=>nx8826);
   ix8657 : inv02 port map ( Y=>nx8658, A=>nx8826);
   ix8659 : inv02 port map ( Y=>nx8660, A=>nx8826);
   ix8661 : inv02 port map ( Y=>nx8662, A=>nx8826);
   ix8663 : inv02 port map ( Y=>nx8664, A=>nx8826);
   ix8665 : inv02 port map ( Y=>nx8666, A=>nx8826);
   ix8667 : inv02 port map ( Y=>nx8668, A=>nx8826);
   ix8669 : inv02 port map ( Y=>nx8670, A=>nx8828);
   ix8671 : inv02 port map ( Y=>nx8672, A=>nx8828);
   ix8673 : inv02 port map ( Y=>nx8674, A=>nx8828);
   ix8675 : inv02 port map ( Y=>nx8676, A=>nx8828);
   ix8677 : inv02 port map ( Y=>nx8678, A=>nx8828);
   ix8679 : inv02 port map ( Y=>nx8680, A=>nx8828);
   ix8681 : inv02 port map ( Y=>nx8682, A=>nx8828);
   ix8683 : inv02 port map ( Y=>nx8684, A=>nx8830);
   ix8685 : inv02 port map ( Y=>nx8686, A=>nx8830);
   ix8687 : inv02 port map ( Y=>nx8688, A=>nx8830);
   ix8689 : inv02 port map ( Y=>nx8690, A=>nx8830);
   ix8691 : inv02 port map ( Y=>nx8692, A=>nx8830);
   ix8695 : inv02 port map ( Y=>nx8696, A=>nx8926);
   ix8697 : inv02 port map ( Y=>nx8698, A=>nx8926);
   ix8699 : inv02 port map ( Y=>nx8700, A=>nx8926);
   ix8701 : inv02 port map ( Y=>nx8702, A=>nx8926);
   ix8703 : inv02 port map ( Y=>nx8704, A=>nx8926);
   ix8705 : inv02 port map ( Y=>nx8706, A=>nx8926);
   ix8707 : inv02 port map ( Y=>nx8708, A=>nx8832);
   ix8709 : inv02 port map ( Y=>nx8710, A=>nx8834);
   ix8711 : inv02 port map ( Y=>nx8712, A=>nx8834);
   ix8713 : inv02 port map ( Y=>nx8714, A=>nx8834);
   ix8715 : inv02 port map ( Y=>nx8716, A=>nx8834);
   ix8717 : inv02 port map ( Y=>nx8718, A=>nx8834);
   ix8719 : inv02 port map ( Y=>nx8720, A=>nx8834);
   ix8721 : inv02 port map ( Y=>nx8722, A=>nx8834);
   ix8723 : inv02 port map ( Y=>nx8724, A=>nx8836);
   ix8725 : inv02 port map ( Y=>nx8726, A=>nx8836);
   ix8727 : inv02 port map ( Y=>nx8728, A=>nx8836);
   ix8729 : inv02 port map ( Y=>nx8730, A=>nx8836);
   ix8731 : inv02 port map ( Y=>nx8732, A=>nx8836);
   ix8733 : inv02 port map ( Y=>nx8734, A=>nx8836);
   ix8735 : inv02 port map ( Y=>nx8736, A=>nx8836);
   ix8737 : inv02 port map ( Y=>nx8738, A=>nx8838);
   ix8739 : inv02 port map ( Y=>nx8740, A=>nx8838);
   ix8741 : inv02 port map ( Y=>nx8742, A=>nx8838);
   ix8743 : inv02 port map ( Y=>nx8744, A=>nx8838);
   ix8745 : inv02 port map ( Y=>nx8746, A=>nx8838);
   ix8747 : inv02 port map ( Y=>nx8748, A=>nx8838);
   ix8749 : inv02 port map ( Y=>nx8750, A=>nx8838);
   ix8751 : inv02 port map ( Y=>nx8752, A=>nx8840);
   ix8753 : inv02 port map ( Y=>nx8754, A=>nx8840);
   ix8755 : inv02 port map ( Y=>nx8756, A=>nx8840);
   ix8757 : inv02 port map ( Y=>nx8758, A=>nx8840);
   ix8759 : inv02 port map ( Y=>nx8760, A=>nx8840);
   ix8761 : inv02 port map ( Y=>nx8762, A=>nx8840);
   ix8763 : inv02 port map ( Y=>nx8764, A=>nx8840);
   ix8765 : inv02 port map ( Y=>nx8766, A=>nx8842);
   ix8767 : inv02 port map ( Y=>nx8768, A=>nx8842);
   ix8769 : inv02 port map ( Y=>nx8770, A=>nx8842);
   ix8771 : inv02 port map ( Y=>nx8772, A=>nx8842);
   ix8773 : inv02 port map ( Y=>nx8774, A=>nx8842);
   ix8775 : inv02 port map ( Y=>nx8776, A=>nx8842);
   ix8777 : inv02 port map ( Y=>nx8778, A=>nx8842);
   ix8779 : inv02 port map ( Y=>nx8780, A=>nx8844);
   ix8781 : inv02 port map ( Y=>nx8782, A=>nx8844);
   ix8783 : inv02 port map ( Y=>nx8784, A=>nx8844);
   ix8785 : inv02 port map ( Y=>nx8786, A=>nx8844);
   ix8787 : inv02 port map ( Y=>nx8788, A=>nx8844);
   ix8789 : inv02 port map ( Y=>nx8790, A=>nx8844);
   ix8791 : inv02 port map ( Y=>nx8792, A=>nx8844);
   ix8793 : inv02 port map ( Y=>nx8794, A=>nx8846);
   ix8795 : inv02 port map ( Y=>nx8796, A=>nx8846);
   ix8797 : inv02 port map ( Y=>nx8798, A=>nx8846);
   ix8799 : inv02 port map ( Y=>nx8800, A=>nx8846);
   ix8801 : inv02 port map ( Y=>nx8802, A=>nx8846);
   ix8803 : inv02 port map ( Y=>nx8804, A=>LayerInfo(15));
   ix8805 : inv02 port map ( Y=>nx8806, A=>nx8856);
   ix8807 : inv02 port map ( Y=>nx8808, A=>nx8856);
   ix8809 : inv02 port map ( Y=>nx8810, A=>nx8856);
   ix8811 : inv02 port map ( Y=>nx8812, A=>nx12);
   ix8813 : inv02 port map ( Y=>nx8814, A=>nx8904);
   ix8815 : inv02 port map ( Y=>nx8816, A=>nx510);
   ix8817 : inv02 port map ( Y=>nx8818, A=>nx510);
   ix8819 : inv02 port map ( Y=>nx8820, A=>nx510);
   ix8821 : inv02 port map ( Y=>nx8822, A=>nx510);
   ix8823 : inv02 port map ( Y=>nx8824, A=>nx510);
   ix8825 : inv02 port map ( Y=>nx8826, A=>nx510);
   ix8827 : inv02 port map ( Y=>nx8828, A=>nx510);
   ix8829 : inv02 port map ( Y=>nx8830, A=>nx510);
   ix8831 : inv02 port map ( Y=>nx8832, A=>nx516);
   ix8833 : inv02 port map ( Y=>nx8834, A=>nx8912);
   ix8835 : inv02 port map ( Y=>nx8836, A=>nx8912);
   ix8837 : inv02 port map ( Y=>nx8838, A=>nx8912);
   ix8839 : inv02 port map ( Y=>nx8840, A=>nx8912);
   ix8841 : inv02 port map ( Y=>nx8842, A=>nx8912);
   ix8843 : inv02 port map ( Y=>nx8844, A=>nx8914);
   ix8845 : inv02 port map ( Y=>nx8846, A=>nx8914);
   ix517 : nor02ii port map ( Y=>nx516, A0=>nx8856, A1=>nx8902);
   ix35 : and02 port map ( Y=>nx34, A0=>nx8892, A1=>nx8856);
   ix21 : nor02ii port map ( Y=>nx20, A0=>nx8892, A1=>nx8906);
   ix49 : nor02ii port map ( Y=>nx48, A0=>nx8892, A1=>nx8856);
   ix255 : and02 port map ( Y=>ConvOuput_15_EXMPLR, A0=>nx8856, A1=>nx6);
   ix8851 : inv02 port map ( Y=>nx8852, A=>nx8804);
   ix8853 : inv02 port map ( Y=>nx8854, A=>nx8804);
   ix8855 : inv02 port map ( Y=>nx8856, A=>nx8804);
   ix8857 : inv02 port map ( Y=>nx8858, A=>nx8916);
   ix8859 : inv02 port map ( Y=>nx8860, A=>nx8916);
   ix8861 : inv02 port map ( Y=>nx8862, A=>nx8916);
   ix8863 : inv02 port map ( Y=>nx8864, A=>nx8918);
   ix8865 : inv02 port map ( Y=>nx8866, A=>nx8918);
   ix8867 : inv02 port map ( Y=>nx8868, A=>nx8918);
   ix8869 : inv02 port map ( Y=>nx8870, A=>nx8918);
   ix8871 : inv02 port map ( Y=>nx8872, A=>nx8918);
   ix8873 : inv02 port map ( Y=>nx8874, A=>nx8918);
   ix8875 : inv02 port map ( Y=>nx8876, A=>nx8918);
   ix8877 : inv02 port map ( Y=>nx8878, A=>nx8920);
   ix8879 : inv02 port map ( Y=>nx8880, A=>nx8920);
   ix8881 : inv02 port map ( Y=>nx8882, A=>nx8920);
   ix8883 : inv02 port map ( Y=>nx8884, A=>nx8920);
   ix8885 : inv02 port map ( Y=>nx8886, A=>nx8920);
   ix8887 : inv02 port map ( Y=>nx8888, A=>nx8920);
   ix8889 : inv02 port map ( Y=>nx8890, A=>nx8920);
   ix8891 : inv02 port map ( Y=>nx8892, A=>nx8922);
   ix8893 : inv01 port map ( Y=>nx8894, A=>QImgStat);
   ix8895 : inv02 port map ( Y=>nx8896, A=>nx8894);
   ix8897 : inv02 port map ( Y=>nx8898, A=>nx8894);
   ix8899 : inv02 port map ( Y=>nx8900, A=>nx8894);
   ix8901 : inv02 port map ( Y=>nx8902, A=>nx8894);
   ix8903 : inv02 port map ( Y=>nx8904, A=>nx8812);
   ix8905 : inv02 port map ( Y=>nx8906, A=>nx8812);
   ix8907 : buf02 port map ( Y=>nx8908, A=>nx48);
   ix8909 : buf02 port map ( Y=>nx8910, A=>nx48);
   ix8911 : inv01 port map ( Y=>nx8912, A=>nx8926);
   ix8913 : inv01 port map ( Y=>nx8914, A=>nx8832);
   ix8915 : inv02 port map ( Y=>nx8916, A=>LayerInfo(14));
   ix8917 : inv02 port map ( Y=>nx8918, A=>LayerInfo(14));
   ix8919 : inv02 port map ( Y=>nx8920, A=>LayerInfo(14));
   ix8921 : inv02 port map ( Y=>nx8922, A=>LayerInfo(14));
   ix8923 : inv02 port map ( Y=>nx8924, A=>LayerInfo(15));
   ix8925 : inv02 port map ( Y=>nx8926, A=>nx516);
end ConvArch ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Counter_5 is
   port (
      enable : IN std_logic ;
      reset : IN std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      output : OUT std_logic_vector (4 DOWNTO 0) ;
      input : IN std_logic_vector (4 DOWNTO 0)) ;
end Counter_5 ;

architecture CounterImplementation of Counter_5 is
   component my_nadder_5
      port (
         a : IN std_logic_vector (4 DOWNTO 0) ;
         b : IN std_logic_vector (4 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (4 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal output_4_EXMPLR, output_3_EXMPLR, output_2_EXMPLR, output_1_EXMPLR, 
      output_0_EXMPLR, addResult_4, addResult_3, addResult_2, addResult_1, 
      addResult_0, one_0, one_4, nx64, NOT_clk, nx8, nx12, nx58, nx20, nx24, 
      nx52, nx32, nx36, nx46, nx44, nx49, nx40, nx57, nx61, nx172, nx182, 
      nx192, nx202, nx212, nx221, nx262, nx268, nx270: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   output(4) <= output_4_EXMPLR ;
   output(3) <= output_3_EXMPLR ;
   output(2) <= output_2_EXMPLR ;
   output(1) <= output_1_EXMPLR ;
   output(0) <= output_0_EXMPLR ;
   A1 : my_nadder_5 port map ( a(4)=>output_4_EXMPLR, a(3)=>output_3_EXMPLR, 
      a(2)=>output_2_EXMPLR, a(1)=>output_1_EXMPLR, a(0)=>output_0_EXMPLR, 
      b(4)=>one_4, b(3)=>one_4, b(2)=>one_4, b(1)=>one_4, b(0)=>one_0, cin=>
      one_4, s(4)=>addResult_4, s(3)=>addResult_3, s(2)=>addResult_2, s(1)=>
      addResult_1, s(0)=>addResult_0, cout=>DANGLING(0));
   ix146 : fake_gnd port map ( Y=>one_4);
   ix144 : fake_vcc port map ( Y=>one_0);
   reg_toOutput_0_dup_1 : dffsr_ni port map ( Q=>output_0_EXMPLR, QB=>OPEN, 
      D=>nx172, CLK=>clk, S=>nx8, R=>nx12);
   ix173 : mux21_ni port map ( Y=>nx172, A0=>output_0_EXMPLR, A1=>
      addResult_0, S0=>nx268);
   ix9 : nor02ii port map ( Y=>nx8, A0=>nx262, A1=>nx64);
   ix222 : nor02_2x port map ( Y=>nx221, A0=>nx270, A1=>load);
   ix65 : dffr port map ( Q=>nx64, QB=>OPEN, D=>input(0), CLK=>NOT_clk, R=>
      nx270);
   ix225 : inv01 port map ( Y=>NOT_clk, A=>clk);
   ix13 : nor02_2x port map ( Y=>nx12, A0=>nx64, A1=>nx262);
   reg_toOutput_1_dup_1 : dffsr_ni port map ( Q=>output_1_EXMPLR, QB=>OPEN, 
      D=>nx182, CLK=>clk, S=>nx20, R=>nx24);
   ix183 : mux21_ni port map ( Y=>nx182, A0=>output_1_EXMPLR, A1=>
      addResult_1, S0=>nx268);
   ix21 : nor02ii port map ( Y=>nx20, A0=>nx262, A1=>nx58);
   ix59 : dffr port map ( Q=>nx58, QB=>OPEN, D=>input(1), CLK=>NOT_clk, R=>
      nx270);
   ix25 : nor02_2x port map ( Y=>nx24, A0=>nx58, A1=>nx262);
   reg_toOutput_2_dup_1 : dffsr_ni port map ( Q=>output_2_EXMPLR, QB=>OPEN, 
      D=>nx192, CLK=>clk, S=>nx32, R=>nx36);
   ix193 : mux21_ni port map ( Y=>nx192, A0=>output_2_EXMPLR, A1=>
      addResult_2, S0=>nx268);
   ix33 : nor02ii port map ( Y=>nx32, A0=>nx262, A1=>nx52);
   ix53 : dffr port map ( Q=>nx52, QB=>OPEN, D=>input(2), CLK=>NOT_clk, R=>
      nx270);
   ix37 : nor02_2x port map ( Y=>nx36, A0=>nx52, A1=>nx262);
   reg_toOutput_3_dup_1 : dffsr_ni port map ( Q=>output_3_EXMPLR, QB=>OPEN, 
      D=>nx202, CLK=>clk, S=>nx44, R=>nx49);
   ix203 : mux21_ni port map ( Y=>nx202, A0=>output_3_EXMPLR, A1=>
      addResult_3, S0=>nx268);
   ix45 : nor02ii port map ( Y=>nx44, A0=>nx262, A1=>nx46);
   ix47 : dffr port map ( Q=>nx46, QB=>OPEN, D=>input(3), CLK=>NOT_clk, R=>
      nx270);
   ix50 : nor02_2x port map ( Y=>nx49, A0=>nx46, A1=>nx221);
   reg_toOutput_4_dup_1 : dffsr_ni port map ( Q=>output_4_EXMPLR, QB=>OPEN, 
      D=>nx212, CLK=>clk, S=>nx57, R=>nx61);
   ix213 : mux21_ni port map ( Y=>nx212, A0=>output_4_EXMPLR, A1=>
      addResult_4, S0=>nx268);
   ix58 : nor02ii port map ( Y=>nx57, A0=>nx221, A1=>nx40);
   ix54 : dffr port map ( Q=>nx40, QB=>OPEN, D=>input(4), CLK=>NOT_clk, R=>
      nx270);
   ix62 : nor02_2x port map ( Y=>nx61, A0=>nx40, A1=>nx221);
   ix261 : nor02_2x port map ( Y=>nx262, A0=>nx270, A1=>load);
   ix267 : buf02 port map ( Y=>nx268, A=>enable);
   ix269 : buf02 port map ( Y=>nx270, A=>reset);
end CounterImplementation ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Counter_13 is
   port (
      enable : IN std_logic ;
      reset : IN std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      output : OUT std_logic_vector (12 DOWNTO 0) ;
      input : IN std_logic_vector (12 DOWNTO 0)) ;
end Counter_13 ;

architecture CounterImplementation of Counter_13 is
   component my_nadder_13
      port (
         a : IN std_logic_vector (12 DOWNTO 0) ;
         b : IN std_logic_vector (12 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (12 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal output_12_EXMPLR, output_11_EXMPLR, output_10_EXMPLR, 
      output_9_EXMPLR, output_8_EXMPLR, output_7_EXMPLR, output_6_EXMPLR, 
      output_5_EXMPLR, output_4_EXMPLR, output_3_EXMPLR, output_2_EXMPLR, 
      output_1_EXMPLR, output_0_EXMPLR, addResult_12, addResult_11, 
      addResult_10, addResult_9, addResult_8, addResult_7, addResult_6, 
      addResult_5, addResult_4, addResult_3, addResult_2, addResult_1, 
      addResult_0, one_0, one_12, nx160, nx8, nx12, nx154, nx20, nx24, nx148, 
      nx32, nx36, nx142, nx44, nx48, nx136, nx56, nx60, nx130, nx68, nx72, 
      nx124, nx80, nx84, nx118, nx92, nx96, nx112, nx104, nx108, nx106, 
      nx117, nx121, nx100, nx129, nx133, nx94, nx141, nx145, nx88, nx153, 
      nx157, nx404, nx414, nx424, nx434, nx444, nx454, nx464, nx474, nx484, 
      nx494, nx504, nx514, nx524, nx533, nx630, nx632, nx634, nx648, nx650, 
      nx652, nx654, nx656, nx658, nx660, nx662, nx664, nx666, nx668: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   output(12) <= output_12_EXMPLR ;
   output(11) <= output_11_EXMPLR ;
   output(10) <= output_10_EXMPLR ;
   output(9) <= output_9_EXMPLR ;
   output(8) <= output_8_EXMPLR ;
   output(7) <= output_7_EXMPLR ;
   output(6) <= output_6_EXMPLR ;
   output(5) <= output_5_EXMPLR ;
   output(4) <= output_4_EXMPLR ;
   output(3) <= output_3_EXMPLR ;
   output(2) <= output_2_EXMPLR ;
   output(1) <= output_1_EXMPLR ;
   output(0) <= output_0_EXMPLR ;
   A1 : my_nadder_13 port map ( a(12)=>output_12_EXMPLR, a(11)=>
      output_11_EXMPLR, a(10)=>output_10_EXMPLR, a(9)=>output_9_EXMPLR, a(8)
      =>output_8_EXMPLR, a(7)=>output_7_EXMPLR, a(6)=>output_6_EXMPLR, a(5)
      =>output_5_EXMPLR, a(4)=>output_4_EXMPLR, a(3)=>output_3_EXMPLR, a(2)
      =>output_2_EXMPLR, a(1)=>output_1_EXMPLR, a(0)=>output_0_EXMPLR, b(12)
      =>one_12, b(11)=>one_12, b(10)=>one_12, b(9)=>one_12, b(8)=>one_12, 
      b(7)=>one_12, b(6)=>one_12, b(5)=>one_12, b(4)=>one_12, b(3)=>one_12, 
      b(2)=>one_12, b(1)=>one_12, b(0)=>one_0, cin=>one_12, s(12)=>
      addResult_12, s(11)=>addResult_11, s(10)=>addResult_10, s(9)=>
      addResult_9, s(8)=>addResult_8, s(7)=>addResult_7, s(6)=>addResult_6, 
      s(5)=>addResult_5, s(4)=>addResult_4, s(3)=>addResult_3, s(2)=>
      addResult_2, s(1)=>addResult_1, s(0)=>addResult_0, cout=>DANGLING(0));
   ix354 : fake_gnd port map ( Y=>one_12);
   ix352 : fake_vcc port map ( Y=>one_0);
   reg_toOutput_0_dup_1 : dffsr_ni port map ( Q=>output_0_EXMPLR, QB=>OPEN, 
      D=>nx404, CLK=>nx648, S=>nx8, R=>nx12);
   ix405 : mux21_ni port map ( Y=>nx404, A0=>output_0_EXMPLR, A1=>
      addResult_0, S0=>nx658);
   ix534 : nor02_2x port map ( Y=>nx533, A0=>nx654, A1=>load);
   ix161 : dffr port map ( Q=>nx160, QB=>OPEN, D=>input(0), CLK=>nx662, R=>
      nx654);
   reg_toOutput_1_dup_1 : dffsr_ni port map ( Q=>output_1_EXMPLR, QB=>OPEN, 
      D=>nx414, CLK=>nx648, S=>nx20, R=>nx24);
   ix415 : mux21_ni port map ( Y=>nx414, A0=>output_1_EXMPLR, A1=>
      addResult_1, S0=>nx658);
   ix155 : dffr port map ( Q=>nx154, QB=>OPEN, D=>input(1), CLK=>nx662, R=>
      nx654);
   reg_toOutput_2_dup_1 : dffsr_ni port map ( Q=>output_2_EXMPLR, QB=>OPEN, 
      D=>nx424, CLK=>nx648, S=>nx32, R=>nx36);
   ix425 : mux21_ni port map ( Y=>nx424, A0=>output_2_EXMPLR, A1=>
      addResult_2, S0=>nx658);
   ix149 : dffr port map ( Q=>nx148, QB=>OPEN, D=>input(2), CLK=>nx662, R=>
      nx654);
   reg_toOutput_3_dup_1 : dffsr_ni port map ( Q=>output_3_EXMPLR, QB=>OPEN, 
      D=>nx434, CLK=>nx648, S=>nx44, R=>nx48);
   ix435 : mux21_ni port map ( Y=>nx434, A0=>output_3_EXMPLR, A1=>
      addResult_3, S0=>nx658);
   ix143 : dffr port map ( Q=>nx142, QB=>OPEN, D=>input(3), CLK=>nx662, R=>
      nx654);
   reg_toOutput_4_dup_1 : dffsr_ni port map ( Q=>output_4_EXMPLR, QB=>OPEN, 
      D=>nx444, CLK=>nx648, S=>nx56, R=>nx60);
   ix445 : mux21_ni port map ( Y=>nx444, A0=>output_4_EXMPLR, A1=>
      addResult_4, S0=>nx658);
   ix137 : dffr port map ( Q=>nx136, QB=>OPEN, D=>input(4), CLK=>nx662, R=>
      nx654);
   reg_toOutput_5_dup_1 : dffsr_ni port map ( Q=>output_5_EXMPLR, QB=>OPEN, 
      D=>nx454, CLK=>nx650, S=>nx68, R=>nx72);
   ix455 : mux21_ni port map ( Y=>nx454, A0=>output_5_EXMPLR, A1=>
      addResult_5, S0=>nx658);
   ix131 : dffr port map ( Q=>nx130, QB=>OPEN, D=>input(5), CLK=>nx662, R=>
      nx654);
   reg_toOutput_6_dup_1 : dffsr_ni port map ( Q=>output_6_EXMPLR, QB=>OPEN, 
      D=>nx464, CLK=>nx650, S=>nx80, R=>nx84);
   ix465 : mux21_ni port map ( Y=>nx464, A0=>output_6_EXMPLR, A1=>
      addResult_6, S0=>nx658);
   ix125 : dffr port map ( Q=>nx124, QB=>OPEN, D=>input(6), CLK=>nx662, R=>
      nx656);
   reg_toOutput_7_dup_1 : dffsr_ni port map ( Q=>output_7_EXMPLR, QB=>OPEN, 
      D=>nx474, CLK=>nx650, S=>nx92, R=>nx96);
   ix475 : mux21_ni port map ( Y=>nx474, A0=>output_7_EXMPLR, A1=>
      addResult_7, S0=>nx660);
   ix119 : dffr port map ( Q=>nx118, QB=>OPEN, D=>input(7), CLK=>nx632, R=>
      nx656);
   reg_toOutput_8_dup_1 : dffsr_ni port map ( Q=>output_8_EXMPLR, QB=>OPEN, 
      D=>nx484, CLK=>nx650, S=>nx104, R=>nx108);
   ix485 : mux21_ni port map ( Y=>nx484, A0=>output_8_EXMPLR, A1=>
      addResult_8, S0=>nx660);
   ix113 : dffr port map ( Q=>nx112, QB=>OPEN, D=>input(8), CLK=>nx632, R=>
      nx656);
   reg_toOutput_9_dup_1 : dffsr_ni port map ( Q=>output_9_EXMPLR, QB=>OPEN, 
      D=>nx494, CLK=>nx650, S=>nx117, R=>nx121);
   ix495 : mux21_ni port map ( Y=>nx494, A0=>output_9_EXMPLR, A1=>
      addResult_9, S0=>nx660);
   ix114 : dffr port map ( Q=>nx106, QB=>OPEN, D=>input(9), CLK=>nx632, R=>
      nx656);
   reg_toOutput_10_dup_1 : dffsr_ni port map ( Q=>output_10_EXMPLR, QB=>OPEN, 
      D=>nx504, CLK=>nx652, S=>nx129, R=>nx133);
   ix505 : mux21_ni port map ( Y=>nx504, A0=>output_10_EXMPLR, A1=>
      addResult_10, S0=>nx660);
   ix126 : dffr port map ( Q=>nx100, QB=>OPEN, D=>input(10), CLK=>nx632, R=>
      nx656);
   reg_toOutput_11_dup_1 : dffsr_ni port map ( Q=>output_11_EXMPLR, QB=>OPEN, 
      D=>nx514, CLK=>nx652, S=>nx141, R=>nx145);
   ix515 : mux21_ni port map ( Y=>nx514, A0=>output_11_EXMPLR, A1=>
      addResult_11, S0=>nx660);
   ix138 : dffr port map ( Q=>nx94, QB=>OPEN, D=>input(11), CLK=>nx632, R=>
      nx656);
   reg_toOutput_12_dup_1 : dffsr_ni port map ( Q=>output_12_EXMPLR, QB=>OPEN, 
      D=>nx524, CLK=>nx652, S=>nx153, R=>nx157);
   ix525 : mux21_ni port map ( Y=>nx524, A0=>output_12_EXMPLR, A1=>
      addResult_12, S0=>nx660);
   ix150 : dffr port map ( Q=>nx88, QB=>OPEN, D=>input(12), CLK=>nx632, R=>
      nx656);
   ix629 : inv02 port map ( Y=>nx630, A=>clk);
   ix631 : inv02 port map ( Y=>nx632, A=>nx652);
   ix633 : inv01 port map ( Y=>nx634, A=>nx533);
   ix9 : and02 port map ( Y=>nx8, A0=>nx664, A1=>nx160);
   ix13 : nor02ii port map ( Y=>nx12, A0=>nx160, A1=>nx664);
   ix21 : and02 port map ( Y=>nx20, A0=>nx664, A1=>nx154);
   ix25 : nor02ii port map ( Y=>nx24, A0=>nx154, A1=>nx664);
   ix33 : and02 port map ( Y=>nx32, A0=>nx664, A1=>nx148);
   ix37 : nor02ii port map ( Y=>nx36, A0=>nx148, A1=>nx664);
   ix45 : and02 port map ( Y=>nx44, A0=>nx664, A1=>nx142);
   ix49 : nor02ii port map ( Y=>nx48, A0=>nx142, A1=>nx666);
   ix57 : and02 port map ( Y=>nx56, A0=>nx666, A1=>nx136);
   ix61 : nor02ii port map ( Y=>nx60, A0=>nx136, A1=>nx666);
   ix69 : and02 port map ( Y=>nx68, A0=>nx666, A1=>nx130);
   ix73 : nor02ii port map ( Y=>nx72, A0=>nx130, A1=>nx666);
   ix81 : and02 port map ( Y=>nx80, A0=>nx666, A1=>nx124);
   ix85 : nor02ii port map ( Y=>nx84, A0=>nx124, A1=>nx666);
   ix93 : and02 port map ( Y=>nx92, A0=>nx668, A1=>nx118);
   ix97 : nor02ii port map ( Y=>nx96, A0=>nx118, A1=>nx668);
   ix105 : and02 port map ( Y=>nx104, A0=>nx668, A1=>nx112);
   ix109 : nor02ii port map ( Y=>nx108, A0=>nx112, A1=>nx668);
   ix118 : and02 port map ( Y=>nx117, A0=>nx668, A1=>nx106);
   ix122 : nor02ii port map ( Y=>nx121, A0=>nx106, A1=>nx668);
   ix130 : and02 port map ( Y=>nx129, A0=>nx668, A1=>nx100);
   ix134 : nor02ii port map ( Y=>nx133, A0=>nx100, A1=>nx634);
   ix142 : and02 port map ( Y=>nx141, A0=>nx634, A1=>nx94);
   ix146 : nor02ii port map ( Y=>nx145, A0=>nx94, A1=>nx634);
   ix154 : and02 port map ( Y=>nx153, A0=>nx634, A1=>nx88);
   ix158 : nor02ii port map ( Y=>nx157, A0=>nx88, A1=>nx634);
   ix647 : inv01 port map ( Y=>nx648, A=>nx630);
   ix649 : inv01 port map ( Y=>nx650, A=>nx630);
   ix651 : inv01 port map ( Y=>nx652, A=>nx630);
   ix653 : buf02 port map ( Y=>nx654, A=>reset);
   ix655 : buf02 port map ( Y=>nx656, A=>reset);
   ix657 : buf02 port map ( Y=>nx658, A=>enable);
   ix659 : buf02 port map ( Y=>nx660, A=>enable);
   ix661 : inv02 port map ( Y=>nx662, A=>clk);
   ix663 : inv01 port map ( Y=>nx664, A=>nx533);
   ix665 : inv01 port map ( Y=>nx666, A=>nx533);
   ix667 : inv01 port map ( Y=>nx668, A=>nx533);
end CounterImplementation ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity addressCounter is
   port (
      reset : IN std_logic ;
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      outputAddress : OUT std_logic_vector (12 DOWNTO 0) ;
      RealOutputCounter : OUT std_logic_vector (12 DOWNTO 0) ;
      AddresCounterLoad : IN std_logic_vector (12 DOWNTO 0) ;
      X : IN std_logic ;
      Y : IN std_logic ;
      clk : IN std_logic) ;
end addressCounter ;

architecture addressCounterArch of addressCounter is
   component Counter_13
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (12 DOWNTO 0) ;
         input : IN std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   signal RealOutputCounter_12_EXMPLR, RealOutputCounter_11_EXMPLR, 
      RealOutputCounter_10_EXMPLR, RealOutputCounter_9_EXMPLR, 
      RealOutputCounter_8_EXMPLR, RealOutputCounter_7_EXMPLR, 
      RealOutputCounter_6_EXMPLR, RealOutputCounter_5_EXMPLR, 
      RealOutputCounter_4_EXMPLR, RealOutputCounter_3_EXMPLR, 
      RealOutputCounter_2_EXMPLR, RealOutputCounter_1_EXMPLR, 
      RealOutputCounter_0_EXMPLR, CounterClk, CounterRest, Load, nx110: 
   std_logic ;

begin
   RealOutputCounter(12) <= RealOutputCounter_12_EXMPLR ;
   RealOutputCounter(11) <= RealOutputCounter_11_EXMPLR ;
   RealOutputCounter(10) <= RealOutputCounter_10_EXMPLR ;
   RealOutputCounter(9) <= RealOutputCounter_9_EXMPLR ;
   RealOutputCounter(8) <= RealOutputCounter_8_EXMPLR ;
   RealOutputCounter(7) <= RealOutputCounter_7_EXMPLR ;
   RealOutputCounter(6) <= RealOutputCounter_6_EXMPLR ;
   RealOutputCounter(5) <= RealOutputCounter_5_EXMPLR ;
   RealOutputCounter(4) <= RealOutputCounter_4_EXMPLR ;
   RealOutputCounter(3) <= RealOutputCounter_3_EXMPLR ;
   RealOutputCounter(2) <= RealOutputCounter_2_EXMPLR ;
   RealOutputCounter(1) <= RealOutputCounter_1_EXMPLR ;
   RealOutputCounter(0) <= RealOutputCounter_0_EXMPLR ;
   myCounter : Counter_13 port map ( enable=>current_state(8), reset=>
      CounterRest, clk=>CounterClk, load=>Load, output(12)=>
      RealOutputCounter_12_EXMPLR, output(11)=>RealOutputCounter_11_EXMPLR, 
      output(10)=>RealOutputCounter_10_EXMPLR, output(9)=>
      RealOutputCounter_9_EXMPLR, output(8)=>RealOutputCounter_8_EXMPLR, 
      output(7)=>RealOutputCounter_7_EXMPLR, output(6)=>
      RealOutputCounter_6_EXMPLR, output(5)=>RealOutputCounter_5_EXMPLR, 
      output(4)=>RealOutputCounter_4_EXMPLR, output(3)=>
      RealOutputCounter_3_EXMPLR, output(2)=>RealOutputCounter_2_EXMPLR, 
      output(1)=>RealOutputCounter_1_EXMPLR, output(0)=>
      RealOutputCounter_0_EXMPLR, input(12)=>AddresCounterLoad(12), 
      input(11)=>AddresCounterLoad(11), input(10)=>AddresCounterLoad(10), 
      input(9)=>AddresCounterLoad(9), input(8)=>AddresCounterLoad(8), 
      input(7)=>AddresCounterLoad(7), input(6)=>AddresCounterLoad(6), 
      input(5)=>AddresCounterLoad(5), input(4)=>AddresCounterLoad(4), 
      input(3)=>AddresCounterLoad(3), input(2)=>AddresCounterLoad(2), 
      input(1)=>AddresCounterLoad(1), input(0)=>AddresCounterLoad(0));
   outOfAddressCounter : triStateBuffer_13 port map ( D(12)=>
      RealOutputCounter_12_EXMPLR, D(11)=>RealOutputCounter_11_EXMPLR, D(10)
      =>RealOutputCounter_10_EXMPLR, D(9)=>RealOutputCounter_9_EXMPLR, D(8)
      =>RealOutputCounter_8_EXMPLR, D(7)=>RealOutputCounter_7_EXMPLR, D(6)=>
      RealOutputCounter_6_EXMPLR, D(5)=>RealOutputCounter_5_EXMPLR, D(4)=>
      RealOutputCounter_4_EXMPLR, D(3)=>RealOutputCounter_3_EXMPLR, D(2)=>
      RealOutputCounter_2_EXMPLR, D(1)=>RealOutputCounter_1_EXMPLR, D(0)=>
      RealOutputCounter_0_EXMPLR, EN=>current_state(8), F(12)=>
      outputAddress(12), F(11)=>outputAddress(11), F(10)=>outputAddress(10), 
      F(9)=>outputAddress(9), F(8)=>outputAddress(8), F(7)=>outputAddress(7), 
      F(6)=>outputAddress(6), F(5)=>outputAddress(5), F(4)=>outputAddress(4), 
      F(3)=>outputAddress(3), F(2)=>outputAddress(2), F(1)=>outputAddress(1), 
      F(0)=>outputAddress(0));
   ix11 : aoi21 port map ( Y=>Load, A0=>X, A1=>Y, B0=>nx110);
   ix111 : inv01 port map ( Y=>nx110, A=>current_state(9));
   ix13 : or02 port map ( Y=>CounterRest, A0=>reset, A1=>current_state(12));
   ix3 : ao21 port map ( Y=>CounterClk, A0=>clk, A1=>current_state(9), B0=>
      current_state(8));
end addressCounterArch ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity depthNotZero is
   port (
      fromOutDMA : IN std_logic_vector (15 DOWNTO 0) ;
      fromOutReg : IN std_logic_vector (15 DOWNTO 0) ;
      Depth : IN std_logic_vector (3 DOWNTO 0) ;
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      output : OUT std_logic_vector (15 DOWNTO 0)) ;
end depthNotZero ;

architecture DepthNotZeroArch of depthNotZero is
   component my_nadder_16
      port (
         a : IN std_logic_vector (15 DOWNTO 0) ;
         b : IN std_logic_vector (15 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (15 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component triStateBuffer_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal outputAdder_15, outputAdder_14, outputAdder_13, outputAdder_12, 
      outputAdder_11, outputAdder_10, outputAdder_9, outputAdder_8, 
      outputAdder_7, outputAdder_6, outputAdder_5, outputAdder_4, 
      outputAdder_3, outputAdder_2, outputAdder_1, outputAdder_0, Enable, 
      GND, nx117: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   myNadder : my_nadder_16 port map ( a(15)=>fromOutReg(15), a(14)=>
      fromOutReg(14), a(13)=>fromOutReg(13), a(12)=>fromOutReg(12), a(11)=>
      fromOutReg(11), a(10)=>fromOutReg(10), a(9)=>fromOutReg(9), a(8)=>
      fromOutReg(8), a(7)=>fromOutReg(7), a(6)=>fromOutReg(6), a(5)=>
      fromOutReg(5), a(4)=>fromOutReg(4), a(3)=>fromOutReg(3), a(2)=>
      fromOutReg(2), a(1)=>fromOutReg(1), a(0)=>fromOutReg(0), b(15)=>
      fromOutDMA(15), b(14)=>fromOutDMA(14), b(13)=>fromOutDMA(13), b(12)=>
      fromOutDMA(12), b(11)=>fromOutDMA(11), b(10)=>fromOutDMA(10), b(9)=>
      fromOutDMA(9), b(8)=>fromOutDMA(8), b(7)=>fromOutDMA(7), b(6)=>
      fromOutDMA(6), b(5)=>fromOutDMA(5), b(4)=>fromOutDMA(4), b(3)=>
      fromOutDMA(3), b(2)=>fromOutDMA(2), b(1)=>fromOutDMA(1), b(0)=>
      fromOutDMA(0), cin=>GND, s(15)=>outputAdder_15, s(14)=>outputAdder_14, 
      s(13)=>outputAdder_13, s(12)=>outputAdder_12, s(11)=>outputAdder_11, 
      s(10)=>outputAdder_10, s(9)=>outputAdder_9, s(8)=>outputAdder_8, s(7)
      =>outputAdder_7, s(6)=>outputAdder_6, s(5)=>outputAdder_5, s(4)=>
      outputAdder_4, s(3)=>outputAdder_3, s(2)=>outputAdder_2, s(1)=>
      outputAdder_1, s(0)=>outputAdder_0, cout=>DANGLING(0));
   depth0 : triStateBuffer_16 port map ( D(15)=>outputAdder_15, D(14)=>
      outputAdder_14, D(13)=>outputAdder_13, D(12)=>outputAdder_12, D(11)=>
      outputAdder_11, D(10)=>outputAdder_10, D(9)=>outputAdder_9, D(8)=>
      outputAdder_8, D(7)=>outputAdder_7, D(6)=>outputAdder_6, D(5)=>
      outputAdder_5, D(4)=>outputAdder_4, D(3)=>outputAdder_3, D(2)=>
      outputAdder_2, D(1)=>outputAdder_1, D(0)=>outputAdder_0, EN=>Enable, 
      F(15)=>output(15), F(14)=>output(14), F(13)=>output(13), F(12)=>
      output(12), F(11)=>output(11), F(10)=>output(10), F(9)=>output(9), 
      F(8)=>output(8), F(7)=>output(7), F(6)=>output(6), F(5)=>output(5), 
      F(4)=>output(4), F(3)=>output(3), F(2)=>output(2), F(1)=>output(1), 
      F(0)=>output(0));
   ix104 : fake_gnd port map ( Y=>GND);
   ix7 : nor02ii port map ( Y=>Enable, A0=>nx117, A1=>current_state(8));
   ix118 : nor04 port map ( Y=>nx117, A0=>Depth(0), A1=>Depth(1), A2=>
      Depth(2), A3=>Depth(3));
end DepthNotZeroArch ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity mux7 is
   port (
      a1 : IN std_logic_vector (15 DOWNTO 0) ;
      a2 : IN std_logic_vector (15 DOWNTO 0) ;
      a3 : IN std_logic_vector (15 DOWNTO 0) ;
      a4 : IN std_logic_vector (15 DOWNTO 0) ;
      a5 : IN std_logic_vector (15 DOWNTO 0) ;
      a6 : IN std_logic_vector (15 DOWNTO 0) ;
      a7 : IN std_logic_vector (15 DOWNTO 0) ;
      a8 : IN std_logic_vector (15 DOWNTO 0) ;
      sel : IN std_logic_vector (3 DOWNTO 0) ;
      output : OUT std_logic_vector (15 DOWNTO 0)) ;
end mux7 ;

architecture mux7Arch of mux7 is
   signal nx12, nx18, nx80, nx217, nx221, nx223, nx227, nx231, nx233, nx239, 
      nx241, nx247, nx255, nx257, nx259, nx261, nx265, nx267, nx269, nx271, 
      nx275, nx277, nx279, nx281, nx285, nx287, nx289, nx291, nx295, nx297, 
      nx299, nx301, nx305, nx307, nx309, nx311, nx315, nx317, nx319, nx321, 
      nx325, nx327, nx329, nx331, nx335, nx337, nx339, nx341, nx345, nx347, 
      nx349, nx351, nx355, nx357, nx359, nx361, nx365, nx367, nx369, nx371, 
      nx375, nx377, nx379, nx381, nx385, nx387, nx389, nx391, nx395, nx397, 
      nx399, nx401, nx408, nx410, nx412, nx414, nx416, nx418, nx421, nx423, 
      nx425, nx427, nx429, nx431, nx433, nx435, nx437, nx439, nx441, nx443, 
      nx445, nx447, nx449, nx451, nx453, nx455, nx457, nx459, nx461, nx463, 
      nx465, nx467: std_logic ;

begin
   ix89 : nand04 port map ( Y=>output(0), A0=>nx217, A1=>nx233, A2=>nx241, 
      A3=>nx247);
   ix218 : aoi22 port map ( Y=>nx217, A0=>a7(0), A1=>nx459, B0=>a8(0), B1=>
      nx465);
   ix222 : inv01 port map ( Y=>nx221, A=>sel(2));
   ix224 : inv01 port map ( Y=>nx223, A=>sel(1));
   ix81 : nand02 port map ( Y=>nx80, A0=>nx227, A1=>nx231);
   ix228 : nand03 port map ( Y=>nx227, A0=>nx18, A1=>sel(2), A2=>sel(1));
   ix19 : nor02ii port map ( Y=>nx18, A0=>sel(3), A1=>sel(0));
   ix232 : inv01 port map ( Y=>nx231, A=>sel(3));
   ix234 : aoi22 port map ( Y=>nx233, A0=>a3(0), A1=>nx451, B0=>a2(0), B1=>
      nx443);
   ix242 : aoi22 port map ( Y=>nx241, A0=>a5(0), A1=>nx435, B0=>a6(0), B1=>
      nx427);
   ix248 : aoi22 port map ( Y=>nx247, A0=>a1(0), A1=>nx410, B0=>a4(0), B1=>
      nx418);
   ix13 : nor04 port map ( Y=>nx12, A0=>sel(3), A1=>sel(0), A2=>sel(2), A3=>
      sel(1));
   ix119 : nand04 port map ( Y=>output(1), A0=>nx255, A1=>nx257, A2=>nx259, 
      A3=>nx261);
   ix256 : aoi22 port map ( Y=>nx255, A0=>a7(1), A1=>nx459, B0=>a8(1), B1=>
      nx465);
   ix258 : aoi22 port map ( Y=>nx257, A0=>a3(1), A1=>nx451, B0=>a2(1), B1=>
      nx443);
   ix260 : aoi22 port map ( Y=>nx259, A0=>a5(1), A1=>nx435, B0=>a6(1), B1=>
      nx427);
   ix262 : aoi22 port map ( Y=>nx261, A0=>a1(1), A1=>nx410, B0=>a4(1), B1=>
      nx418);
   ix149 : nand04 port map ( Y=>output(2), A0=>nx265, A1=>nx267, A2=>nx269, 
      A3=>nx271);
   ix266 : aoi22 port map ( Y=>nx265, A0=>a7(2), A1=>nx459, B0=>a8(2), B1=>
      nx465);
   ix268 : aoi22 port map ( Y=>nx267, A0=>a3(2), A1=>nx451, B0=>a2(2), B1=>
      nx443);
   ix270 : aoi22 port map ( Y=>nx269, A0=>a5(2), A1=>nx435, B0=>a6(2), B1=>
      nx427);
   ix272 : aoi22 port map ( Y=>nx271, A0=>a1(2), A1=>nx410, B0=>a4(2), B1=>
      nx418);
   ix179 : nand04 port map ( Y=>output(3), A0=>nx275, A1=>nx277, A2=>nx279, 
      A3=>nx281);
   ix276 : aoi22 port map ( Y=>nx275, A0=>a7(3), A1=>nx459, B0=>a8(3), B1=>
      nx465);
   ix278 : aoi22 port map ( Y=>nx277, A0=>a3(3), A1=>nx451, B0=>a2(3), B1=>
      nx443);
   ix280 : aoi22 port map ( Y=>nx279, A0=>a5(3), A1=>nx435, B0=>a6(3), B1=>
      nx427);
   ix282 : aoi22 port map ( Y=>nx281, A0=>a1(3), A1=>nx410, B0=>a4(3), B1=>
      nx418);
   ix209 : nand04 port map ( Y=>output(4), A0=>nx285, A1=>nx287, A2=>nx289, 
      A3=>nx291);
   ix286 : aoi22 port map ( Y=>nx285, A0=>a7(4), A1=>nx459, B0=>a8(4), B1=>
      nx465);
   ix288 : aoi22 port map ( Y=>nx287, A0=>a3(4), A1=>nx451, B0=>a2(4), B1=>
      nx443);
   ix290 : aoi22 port map ( Y=>nx289, A0=>a5(4), A1=>nx435, B0=>a6(4), B1=>
      nx427);
   ix292 : aoi22 port map ( Y=>nx291, A0=>a1(4), A1=>nx410, B0=>a4(4), B1=>
      nx418);
   ix239 : nand04 port map ( Y=>output(5), A0=>nx295, A1=>nx297, A2=>nx299, 
      A3=>nx301);
   ix296 : aoi22 port map ( Y=>nx295, A0=>a7(5), A1=>nx459, B0=>a8(5), B1=>
      nx465);
   ix298 : aoi22 port map ( Y=>nx297, A0=>a3(5), A1=>nx451, B0=>a2(5), B1=>
      nx443);
   ix300 : aoi22 port map ( Y=>nx299, A0=>a5(5), A1=>nx435, B0=>a6(5), B1=>
      nx427);
   ix302 : aoi22 port map ( Y=>nx301, A0=>a1(5), A1=>nx410, B0=>a4(5), B1=>
      nx418);
   ix269 : nand04 port map ( Y=>output(6), A0=>nx305, A1=>nx307, A2=>nx309, 
      A3=>nx311);
   ix306 : aoi22 port map ( Y=>nx305, A0=>a7(6), A1=>nx459, B0=>a8(6), B1=>
      nx465);
   ix308 : aoi22 port map ( Y=>nx307, A0=>a3(6), A1=>nx451, B0=>a2(6), B1=>
      nx443);
   ix310 : aoi22 port map ( Y=>nx309, A0=>a5(6), A1=>nx435, B0=>a6(6), B1=>
      nx427);
   ix312 : aoi22 port map ( Y=>nx311, A0=>a1(6), A1=>nx410, B0=>a4(6), B1=>
      nx418);
   ix299 : nand04 port map ( Y=>output(7), A0=>nx315, A1=>nx317, A2=>nx319, 
      A3=>nx321);
   ix316 : aoi22 port map ( Y=>nx315, A0=>a7(7), A1=>nx461, B0=>a8(7), B1=>
      nx467);
   ix318 : aoi22 port map ( Y=>nx317, A0=>a3(7), A1=>nx453, B0=>a2(7), B1=>
      nx445);
   ix320 : aoi22 port map ( Y=>nx319, A0=>a5(7), A1=>nx437, B0=>a6(7), B1=>
      nx429);
   ix322 : aoi22 port map ( Y=>nx321, A0=>a1(7), A1=>nx412, B0=>a4(7), B1=>
      nx421);
   ix329 : nand04 port map ( Y=>output(8), A0=>nx325, A1=>nx327, A2=>nx329, 
      A3=>nx331);
   ix326 : aoi22 port map ( Y=>nx325, A0=>a7(8), A1=>nx461, B0=>a8(8), B1=>
      nx467);
   ix328 : aoi22 port map ( Y=>nx327, A0=>a3(8), A1=>nx453, B0=>a2(8), B1=>
      nx445);
   ix330 : aoi22 port map ( Y=>nx329, A0=>a5(8), A1=>nx437, B0=>a6(8), B1=>
      nx429);
   ix332 : aoi22 port map ( Y=>nx331, A0=>a1(8), A1=>nx412, B0=>a4(8), B1=>
      nx421);
   ix359 : nand04 port map ( Y=>output(9), A0=>nx335, A1=>nx337, A2=>nx339, 
      A3=>nx341);
   ix336 : aoi22 port map ( Y=>nx335, A0=>a7(9), A1=>nx461, B0=>a8(9), B1=>
      nx467);
   ix338 : aoi22 port map ( Y=>nx337, A0=>a3(9), A1=>nx453, B0=>a2(9), B1=>
      nx445);
   ix340 : aoi22 port map ( Y=>nx339, A0=>a5(9), A1=>nx437, B0=>a6(9), B1=>
      nx429);
   ix342 : aoi22 port map ( Y=>nx341, A0=>a1(9), A1=>nx412, B0=>a4(9), B1=>
      nx421);
   ix389 : nand04 port map ( Y=>output(10), A0=>nx345, A1=>nx347, A2=>nx349, 
      A3=>nx351);
   ix346 : aoi22 port map ( Y=>nx345, A0=>a7(10), A1=>nx461, B0=>a8(10), B1
      =>nx467);
   ix348 : aoi22 port map ( Y=>nx347, A0=>a3(10), A1=>nx453, B0=>a2(10), B1
      =>nx445);
   ix350 : aoi22 port map ( Y=>nx349, A0=>a5(10), A1=>nx437, B0=>a6(10), B1
      =>nx429);
   ix352 : aoi22 port map ( Y=>nx351, A0=>a1(10), A1=>nx412, B0=>a4(10), B1
      =>nx421);
   ix419 : nand04 port map ( Y=>output(11), A0=>nx355, A1=>nx357, A2=>nx359, 
      A3=>nx361);
   ix356 : aoi22 port map ( Y=>nx355, A0=>a7(11), A1=>nx461, B0=>a8(11), B1
      =>nx467);
   ix358 : aoi22 port map ( Y=>nx357, A0=>a3(11), A1=>nx453, B0=>a2(11), B1
      =>nx445);
   ix360 : aoi22 port map ( Y=>nx359, A0=>a5(11), A1=>nx437, B0=>a6(11), B1
      =>nx429);
   ix362 : aoi22 port map ( Y=>nx361, A0=>a1(11), A1=>nx412, B0=>a4(11), B1
      =>nx421);
   ix449 : nand04 port map ( Y=>output(12), A0=>nx365, A1=>nx367, A2=>nx369, 
      A3=>nx371);
   ix366 : aoi22 port map ( Y=>nx365, A0=>a7(12), A1=>nx461, B0=>a8(12), B1
      =>nx467);
   ix368 : aoi22 port map ( Y=>nx367, A0=>a3(12), A1=>nx453, B0=>a2(12), B1
      =>nx445);
   ix370 : aoi22 port map ( Y=>nx369, A0=>a5(12), A1=>nx437, B0=>a6(12), B1
      =>nx429);
   ix372 : aoi22 port map ( Y=>nx371, A0=>a1(12), A1=>nx412, B0=>a4(12), B1
      =>nx421);
   ix479 : nand04 port map ( Y=>output(13), A0=>nx375, A1=>nx377, A2=>nx379, 
      A3=>nx381);
   ix376 : aoi22 port map ( Y=>nx375, A0=>a7(13), A1=>nx461, B0=>a8(13), B1
      =>nx467);
   ix378 : aoi22 port map ( Y=>nx377, A0=>a3(13), A1=>nx453, B0=>a2(13), B1
      =>nx445);
   ix380 : aoi22 port map ( Y=>nx379, A0=>a5(13), A1=>nx437, B0=>a6(13), B1
      =>nx429);
   ix382 : aoi22 port map ( Y=>nx381, A0=>a1(13), A1=>nx412, B0=>a4(13), B1
      =>nx421);
   ix509 : nand04 port map ( Y=>output(14), A0=>nx385, A1=>nx387, A2=>nx389, 
      A3=>nx391);
   ix386 : aoi22 port map ( Y=>nx385, A0=>a7(14), A1=>nx463, B0=>a8(14), B1
      =>nx80);
   ix388 : aoi22 port map ( Y=>nx387, A0=>a3(14), A1=>nx455, B0=>a2(14), B1
      =>nx447);
   ix390 : aoi22 port map ( Y=>nx389, A0=>a5(14), A1=>nx439, B0=>a6(14), B1
      =>nx431);
   ix392 : aoi22 port map ( Y=>nx391, A0=>a1(14), A1=>nx414, B0=>a4(14), B1
      =>nx423);
   ix539 : nand04 port map ( Y=>output(15), A0=>nx395, A1=>nx397, A2=>nx399, 
      A3=>nx401);
   ix396 : aoi22 port map ( Y=>nx395, A0=>a7(15), A1=>nx463, B0=>a8(15), B1
      =>nx80);
   ix398 : aoi22 port map ( Y=>nx397, A0=>a3(15), A1=>nx455, B0=>a2(15), B1
      =>nx447);
   ix400 : aoi22 port map ( Y=>nx399, A0=>a5(15), A1=>nx439, B0=>a6(15), B1
      =>nx431);
   ix402 : aoi22 port map ( Y=>nx401, A0=>a1(15), A1=>nx414, B0=>a4(15), B1
      =>nx423);
   ix240 : inv01 port map ( Y=>nx239, A=>nx18);
   ix407 : inv01 port map ( Y=>nx408, A=>nx12);
   ix409 : inv02 port map ( Y=>nx410, A=>nx408);
   ix411 : inv02 port map ( Y=>nx412, A=>nx408);
   ix413 : inv02 port map ( Y=>nx414, A=>nx408);
   ix417 : inv02 port map ( Y=>nx418, A=>nx416);
   ix420 : inv02 port map ( Y=>nx421, A=>nx416);
   ix422 : inv02 port map ( Y=>nx423, A=>nx416);
   ix426 : inv02 port map ( Y=>nx427, A=>nx425);
   ix428 : inv02 port map ( Y=>nx429, A=>nx425);
   ix430 : inv02 port map ( Y=>nx431, A=>nx425);
   ix434 : inv02 port map ( Y=>nx435, A=>nx433);
   ix436 : inv02 port map ( Y=>nx437, A=>nx433);
   ix438 : inv02 port map ( Y=>nx439, A=>nx433);
   ix442 : inv02 port map ( Y=>nx443, A=>nx441);
   ix444 : inv02 port map ( Y=>nx445, A=>nx441);
   ix446 : inv02 port map ( Y=>nx447, A=>nx441);
   ix450 : inv02 port map ( Y=>nx451, A=>nx449);
   ix452 : inv02 port map ( Y=>nx453, A=>nx449);
   ix454 : inv02 port map ( Y=>nx455, A=>nx449);
   ix458 : inv02 port map ( Y=>nx459, A=>nx457);
   ix460 : inv02 port map ( Y=>nx461, A=>nx457);
   ix462 : inv02 port map ( Y=>nx463, A=>nx457);
   ix464 : nand02 port map ( Y=>nx465, A0=>nx227, A1=>nx231);
   ix466 : nand02 port map ( Y=>nx467, A0=>nx227, A1=>nx231);
   ix73 : or04 port map ( Y=>nx457, A0=>sel(3), A1=>sel(0), A2=>nx221, A3=>
      nx223);
   ix68 : or04 port map ( Y=>nx449, A0=>sel(3), A1=>sel(0), A2=>sel(2), A3=>
      nx223);
   ix57 : or03 port map ( Y=>nx441, A0=>nx239, A1=>sel(2), A2=>sel(1));
   ix43 : or04 port map ( Y=>nx433, A0=>sel(3), A1=>sel(0), A2=>nx221, A3=>
      sel(1));
   ix35 : nand03 port map ( Y=>nx425, A0=>nx18, A1=>sel(2), A2=>nx223);
   ix25 : nand03 port map ( Y=>nx416, A0=>nx18, A1=>nx221, A2=>sel(1));
end mux7Arch ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity depthZero is
   port (
      fromOutReg : IN std_logic_vector (15 DOWNTO 0) ;
      bias1 : IN std_logic_vector (15 DOWNTO 0) ;
      bias2 : IN std_logic_vector (15 DOWNTO 0) ;
      bias3 : IN std_logic_vector (15 DOWNTO 0) ;
      bias4 : IN std_logic_vector (15 DOWNTO 0) ;
      bias5 : IN std_logic_vector (15 DOWNTO 0) ;
      bias6 : IN std_logic_vector (15 DOWNTO 0) ;
      bias7 : IN std_logic_vector (15 DOWNTO 0) ;
      bias8 : IN std_logic_vector (15 DOWNTO 0) ;
      counterNumber : IN std_logic_vector (3 DOWNTO 0) ;
      Depth : IN std_logic_vector (3 DOWNTO 0) ;
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      output : OUT std_logic_vector (15 DOWNTO 0)) ;
end depthZero ;

architecture DepthZeroArch of depthZero is
   component mux7
      port (
         a1 : IN std_logic_vector (15 DOWNTO 0) ;
         a2 : IN std_logic_vector (15 DOWNTO 0) ;
         a3 : IN std_logic_vector (15 DOWNTO 0) ;
         a4 : IN std_logic_vector (15 DOWNTO 0) ;
         a5 : IN std_logic_vector (15 DOWNTO 0) ;
         a6 : IN std_logic_vector (15 DOWNTO 0) ;
         a7 : IN std_logic_vector (15 DOWNTO 0) ;
         a8 : IN std_logic_vector (15 DOWNTO 0) ;
         sel : IN std_logic_vector (3 DOWNTO 0) ;
         output : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component my_nadder_16
      port (
         a : IN std_logic_vector (15 DOWNTO 0) ;
         b : IN std_logic_vector (15 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (15 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component triStateBuffer_16
      port (
         D : IN std_logic_vector (15 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal outputMux_15, outputMux_14, outputMux_13, outputMux_12, 
      outputMux_11, outputMux_10, outputMux_9, outputMux_8, outputMux_7, 
      outputMux_6, outputMux_5, outputMux_4, outputMux_3, outputMux_2, 
      outputMux_1, outputMux_0, outputAdder_15, outputAdder_14, 
      outputAdder_13, outputAdder_12, outputAdder_11, outputAdder_10, 
      outputAdder_9, outputAdder_8, outputAdder_7, outputAdder_6, 
      outputAdder_5, outputAdder_4, outputAdder_3, outputAdder_2, 
      outputAdder_1, outputAdder_0, Enable, GND, nx163, nx165: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   myMux : mux7 port map ( a1(15)=>bias1(15), a1(14)=>bias1(14), a1(13)=>
      bias1(13), a1(12)=>bias1(12), a1(11)=>bias1(11), a1(10)=>bias1(10), 
      a1(9)=>bias1(9), a1(8)=>bias1(8), a1(7)=>bias1(7), a1(6)=>bias1(6), 
      a1(5)=>bias1(5), a1(4)=>bias1(4), a1(3)=>bias1(3), a1(2)=>bias1(2), 
      a1(1)=>bias1(1), a1(0)=>bias1(0), a2(15)=>bias2(15), a2(14)=>bias2(14), 
      a2(13)=>bias2(13), a2(12)=>bias2(12), a2(11)=>bias2(11), a2(10)=>
      bias2(10), a2(9)=>bias2(9), a2(8)=>bias2(8), a2(7)=>bias2(7), a2(6)=>
      bias2(6), a2(5)=>bias2(5), a2(4)=>bias2(4), a2(3)=>bias2(3), a2(2)=>
      bias2(2), a2(1)=>bias2(1), a2(0)=>bias2(0), a3(15)=>bias3(15), a3(14)
      =>bias3(14), a3(13)=>bias3(13), a3(12)=>bias3(12), a3(11)=>bias3(11), 
      a3(10)=>bias3(10), a3(9)=>bias3(9), a3(8)=>bias3(8), a3(7)=>bias3(7), 
      a3(6)=>bias3(6), a3(5)=>bias3(5), a3(4)=>bias3(4), a3(3)=>bias3(3), 
      a3(2)=>bias3(2), a3(1)=>bias3(1), a3(0)=>bias3(0), a4(15)=>bias4(15), 
      a4(14)=>bias4(14), a4(13)=>bias4(13), a4(12)=>bias4(12), a4(11)=>
      bias4(11), a4(10)=>bias4(10), a4(9)=>bias4(9), a4(8)=>bias4(8), a4(7)
      =>bias4(7), a4(6)=>bias4(6), a4(5)=>bias4(5), a4(4)=>bias4(4), a4(3)=>
      bias4(3), a4(2)=>bias4(2), a4(1)=>bias4(1), a4(0)=>bias4(0), a5(15)=>
      bias5(15), a5(14)=>bias5(14), a5(13)=>bias5(13), a5(12)=>bias5(12), 
      a5(11)=>bias5(11), a5(10)=>bias5(10), a5(9)=>bias5(9), a5(8)=>bias5(8), 
      a5(7)=>bias5(7), a5(6)=>bias5(6), a5(5)=>bias5(5), a5(4)=>bias5(4), 
      a5(3)=>bias5(3), a5(2)=>bias5(2), a5(1)=>bias5(1), a5(0)=>bias5(0), 
      a6(15)=>bias6(15), a6(14)=>bias6(14), a6(13)=>bias6(13), a6(12)=>
      bias6(12), a6(11)=>bias6(11), a6(10)=>bias6(10), a6(9)=>bias6(9), 
      a6(8)=>bias6(8), a6(7)=>bias6(7), a6(6)=>bias6(6), a6(5)=>bias6(5), 
      a6(4)=>bias6(4), a6(3)=>bias6(3), a6(2)=>bias6(2), a6(1)=>bias6(1), 
      a6(0)=>bias6(0), a7(15)=>bias7(15), a7(14)=>bias7(14), a7(13)=>
      bias7(13), a7(12)=>bias7(12), a7(11)=>bias7(11), a7(10)=>bias7(10), 
      a7(9)=>bias7(9), a7(8)=>bias7(8), a7(7)=>bias7(7), a7(6)=>bias7(6), 
      a7(5)=>bias7(5), a7(4)=>bias7(4), a7(3)=>bias7(3), a7(2)=>bias7(2), 
      a7(1)=>bias7(1), a7(0)=>bias7(0), a8(15)=>bias8(15), a8(14)=>bias8(14), 
      a8(13)=>bias8(13), a8(12)=>bias8(12), a8(11)=>bias8(11), a8(10)=>
      bias8(10), a8(9)=>bias8(9), a8(8)=>bias8(8), a8(7)=>bias8(7), a8(6)=>
      bias8(6), a8(5)=>bias8(5), a8(4)=>bias8(4), a8(3)=>bias8(3), a8(2)=>
      bias8(2), a8(1)=>bias8(1), a8(0)=>bias8(0), sel(3)=>counterNumber(3), 
      sel(2)=>counterNumber(2), sel(1)=>counterNumber(1), sel(0)=>
      counterNumber(0), output(15)=>outputMux_15, output(14)=>outputMux_14, 
      output(13)=>outputMux_13, output(12)=>outputMux_12, output(11)=>
      outputMux_11, output(10)=>outputMux_10, output(9)=>outputMux_9, 
      output(8)=>outputMux_8, output(7)=>outputMux_7, output(6)=>outputMux_6, 
      output(5)=>outputMux_5, output(4)=>outputMux_4, output(3)=>outputMux_3, 
      output(2)=>outputMux_2, output(1)=>outputMux_1, output(0)=>outputMux_0
   );
   myNadder : my_nadder_16 port map ( a(15)=>fromOutReg(15), a(14)=>
      fromOutReg(14), a(13)=>fromOutReg(13), a(12)=>fromOutReg(12), a(11)=>
      fromOutReg(11), a(10)=>fromOutReg(10), a(9)=>fromOutReg(9), a(8)=>
      fromOutReg(8), a(7)=>fromOutReg(7), a(6)=>fromOutReg(6), a(5)=>
      fromOutReg(5), a(4)=>fromOutReg(4), a(3)=>fromOutReg(3), a(2)=>
      fromOutReg(2), a(1)=>fromOutReg(1), a(0)=>fromOutReg(0), b(15)=>
      outputMux_15, b(14)=>outputMux_14, b(13)=>outputMux_13, b(12)=>
      outputMux_12, b(11)=>outputMux_11, b(10)=>outputMux_10, b(9)=>
      outputMux_9, b(8)=>outputMux_8, b(7)=>outputMux_7, b(6)=>outputMux_6, 
      b(5)=>outputMux_5, b(4)=>outputMux_4, b(3)=>outputMux_3, b(2)=>
      outputMux_2, b(1)=>outputMux_1, b(0)=>outputMux_0, cin=>GND, s(15)=>
      outputAdder_15, s(14)=>outputAdder_14, s(13)=>outputAdder_13, s(12)=>
      outputAdder_12, s(11)=>outputAdder_11, s(10)=>outputAdder_10, s(9)=>
      outputAdder_9, s(8)=>outputAdder_8, s(7)=>outputAdder_7, s(6)=>
      outputAdder_6, s(5)=>outputAdder_5, s(4)=>outputAdder_4, s(3)=>
      outputAdder_3, s(2)=>outputAdder_2, s(1)=>outputAdder_1, s(0)=>
      outputAdder_0, cout=>DANGLING(0));
   depth0 : triStateBuffer_16 port map ( D(15)=>outputAdder_15, D(14)=>
      outputAdder_14, D(13)=>outputAdder_13, D(12)=>outputAdder_12, D(11)=>
      outputAdder_11, D(10)=>outputAdder_10, D(9)=>outputAdder_9, D(8)=>
      outputAdder_8, D(7)=>outputAdder_7, D(6)=>outputAdder_6, D(5)=>
      outputAdder_5, D(4)=>outputAdder_4, D(3)=>outputAdder_3, D(2)=>
      outputAdder_2, D(1)=>outputAdder_1, D(0)=>outputAdder_0, EN=>Enable, 
      F(15)=>output(15), F(14)=>output(14), F(13)=>output(13), F(12)=>
      output(12), F(11)=>output(11), F(10)=>output(10), F(9)=>output(9), 
      F(8)=>output(8), F(7)=>output(7), F(6)=>output(6), F(5)=>output(5), 
      F(4)=>output(4), F(3)=>output(3), F(2)=>output(2), F(1)=>output(1), 
      F(0)=>output(0));
   ix150 : fake_gnd port map ( Y=>GND);
   ix15 : nor04 port map ( Y=>Enable, A0=>Depth(1), A1=>Depth(3), A2=>
      Depth(2), A3=>nx163);
   ix164 : nand02 port map ( Y=>nx163, A0=>nx165, A1=>current_state(8));
   ix166 : inv01 port map ( Y=>nx165, A=>Depth(0));
end DepthZeroArch ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity saveState is
   port (
      DMAOutput : IN std_logic_vector (15 DOWNTO 0) ;
      RegisterOutput : IN std_logic_vector (15 DOWNTO 0) ;
      bias1 : IN std_logic_vector (15 DOWNTO 0) ;
      bias2 : IN std_logic_vector (15 DOWNTO 0) ;
      bias3 : IN std_logic_vector (15 DOWNTO 0) ;
      bias4 : IN std_logic_vector (15 DOWNTO 0) ;
      bias5 : IN std_logic_vector (15 DOWNTO 0) ;
      bias6 : IN std_logic_vector (15 DOWNTO 0) ;
      bias7 : IN std_logic_vector (15 DOWNTO 0) ;
      bias8 : IN std_logic_vector (15 DOWNTO 0) ;
      Depth : IN std_logic_vector (3 DOWNTO 0) ;
      NumberOfFiltersCounter : IN std_logic_vector (3 DOWNTO 0) ;
      rst : IN std_logic ;
      stateinput : IN std_logic_vector (14 DOWNTO 0) ;
      clk : IN std_logic ;
      outputCounterToDma : OUT std_logic_vector (12 DOWNTO 0) ;
      RealOutputCounter : OUT std_logic_vector (12 DOWNTO 0) ;
      output : OUT std_logic_vector (15 DOWNTO 0) ;
      ShiftLeftCounterOutput : OUT std_logic_vector (4 DOWNTO 0) ;
      ShiftCounterRst : IN std_logic ;
      AddresCounterLoad : IN std_logic_vector (12 DOWNTO 0) ;
      X : IN std_logic ;
      Y : IN std_logic) ;
end saveState ;

architecture saveStateArch of saveState is
   component Counter_5
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (4 DOWNTO 0) ;
         input : IN std_logic_vector (4 DOWNTO 0)) ;
   end component ;
   component addressCounter
      port (
         reset : IN std_logic ;
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         outputAddress : OUT std_logic_vector (12 DOWNTO 0) ;
         RealOutputCounter : OUT std_logic_vector (12 DOWNTO 0) ;
         AddresCounterLoad : IN std_logic_vector (12 DOWNTO 0) ;
         X : IN std_logic ;
         Y : IN std_logic ;
         clk : IN std_logic) ;
   end component ;
   component depthNotZero
      port (
         fromOutDMA : IN std_logic_vector (15 DOWNTO 0) ;
         fromOutReg : IN std_logic_vector (15 DOWNTO 0) ;
         Depth : IN std_logic_vector (3 DOWNTO 0) ;
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         output : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component depthZero
      port (
         fromOutReg : IN std_logic_vector (15 DOWNTO 0) ;
         bias1 : IN std_logic_vector (15 DOWNTO 0) ;
         bias2 : IN std_logic_vector (15 DOWNTO 0) ;
         bias3 : IN std_logic_vector (15 DOWNTO 0) ;
         bias4 : IN std_logic_vector (15 DOWNTO 0) ;
         bias5 : IN std_logic_vector (15 DOWNTO 0) ;
         bias6 : IN std_logic_vector (15 DOWNTO 0) ;
         bias7 : IN std_logic_vector (15 DOWNTO 0) ;
         bias8 : IN std_logic_vector (15 DOWNTO 0) ;
         counterNumber : IN std_logic_vector (3 DOWNTO 0) ;
         Depth : IN std_logic_vector (3 DOWNTO 0) ;
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         output : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal output_15_EXMPLR, output_14_EXMPLR, output_13_EXMPLR, 
      output_12_EXMPLR, output_11_EXMPLR, output_10_EXMPLR, output_9_EXMPLR, 
      output_8_EXMPLR, output_7_EXMPLR, output_6_EXMPLR, output_5_EXMPLR, 
      output_4_EXMPLR, output_3_EXMPLR, output_2_EXMPLR, output_1_EXMPLR, 
      output_0_EXMPLR, ShiftRegClk, resetCounter, Enable, GND0, nx238, nx240
   : std_logic ;

begin
   output(15) <= output_15_EXMPLR ;
   output(14) <= output_14_EXMPLR ;
   output(13) <= output_13_EXMPLR ;
   output(12) <= output_12_EXMPLR ;
   output(11) <= output_11_EXMPLR ;
   output(10) <= output_10_EXMPLR ;
   output(9) <= output_9_EXMPLR ;
   output(8) <= output_8_EXMPLR ;
   output(7) <= output_7_EXMPLR ;
   output(6) <= output_6_EXMPLR ;
   output(5) <= output_5_EXMPLR ;
   output(4) <= output_4_EXMPLR ;
   output(3) <= output_3_EXMPLR ;
   output(2) <= output_2_EXMPLR ;
   output(1) <= output_1_EXMPLR ;
   output(0) <= output_0_EXMPLR ;
   Scounter : Counter_5 port map ( enable=>Enable, reset=>ShiftCounterRst, 
      clk=>ShiftRegClk, load=>GND0, output(4)=>ShiftLeftCounterOutput(4), 
      output(3)=>ShiftLeftCounterOutput(3), output(2)=>
      ShiftLeftCounterOutput(2), output(1)=>ShiftLeftCounterOutput(1), 
      output(0)=>ShiftLeftCounterOutput(0), input(4)=>GND0, input(3)=>GND0, 
      input(2)=>GND0, input(1)=>GND0, input(0)=>GND0);
   first : addressCounter port map ( reset=>resetCounter, current_state(14)
      =>GND0, current_state(13)=>GND0, current_state(12)=>stateinput(12), 
      current_state(11)=>GND0, current_state(10)=>GND0, current_state(9)=>
      stateinput(9), current_state(8)=>nx238, current_state(7)=>GND0, 
      current_state(6)=>GND0, current_state(5)=>GND0, current_state(4)=>GND0, 
      current_state(3)=>GND0, current_state(2)=>GND0, current_state(1)=>GND0, 
      current_state(0)=>GND0, outputAddress(12)=>outputCounterToDma(12), 
      outputAddress(11)=>outputCounterToDma(11), outputAddress(10)=>
      outputCounterToDma(10), outputAddress(9)=>outputCounterToDma(9), 
      outputAddress(8)=>outputCounterToDma(8), outputAddress(7)=>
      outputCounterToDma(7), outputAddress(6)=>outputCounterToDma(6), 
      outputAddress(5)=>outputCounterToDma(5), outputAddress(4)=>
      outputCounterToDma(4), outputAddress(3)=>outputCounterToDma(3), 
      outputAddress(2)=>outputCounterToDma(2), outputAddress(1)=>
      outputCounterToDma(1), outputAddress(0)=>outputCounterToDma(0), 
      RealOutputCounter(12)=>RealOutputCounter(12), RealOutputCounter(11)=>
      RealOutputCounter(11), RealOutputCounter(10)=>RealOutputCounter(10), 
      RealOutputCounter(9)=>RealOutputCounter(9), RealOutputCounter(8)=>
      RealOutputCounter(8), RealOutputCounter(7)=>RealOutputCounter(7), 
      RealOutputCounter(6)=>RealOutputCounter(6), RealOutputCounter(5)=>
      RealOutputCounter(5), RealOutputCounter(4)=>RealOutputCounter(4), 
      RealOutputCounter(3)=>RealOutputCounter(3), RealOutputCounter(2)=>
      RealOutputCounter(2), RealOutputCounter(1)=>RealOutputCounter(1), 
      RealOutputCounter(0)=>RealOutputCounter(0), AddresCounterLoad(12)=>
      AddresCounterLoad(12), AddresCounterLoad(11)=>AddresCounterLoad(11), 
      AddresCounterLoad(10)=>AddresCounterLoad(10), AddresCounterLoad(9)=>
      AddresCounterLoad(9), AddresCounterLoad(8)=>AddresCounterLoad(8), 
      AddresCounterLoad(7)=>AddresCounterLoad(7), AddresCounterLoad(6)=>
      AddresCounterLoad(6), AddresCounterLoad(5)=>AddresCounterLoad(5), 
      AddresCounterLoad(4)=>AddresCounterLoad(4), AddresCounterLoad(3)=>
      AddresCounterLoad(3), AddresCounterLoad(2)=>AddresCounterLoad(2), 
      AddresCounterLoad(1)=>AddresCounterLoad(1), AddresCounterLoad(0)=>
      AddresCounterLoad(0), X=>X, Y=>Y, clk=>clk);
   second : depthNotZero port map ( fromOutDMA(15)=>DMAOutput(15), 
      fromOutDMA(14)=>DMAOutput(14), fromOutDMA(13)=>DMAOutput(13), 
      fromOutDMA(12)=>DMAOutput(12), fromOutDMA(11)=>DMAOutput(11), 
      fromOutDMA(10)=>DMAOutput(10), fromOutDMA(9)=>DMAOutput(9), 
      fromOutDMA(8)=>DMAOutput(8), fromOutDMA(7)=>DMAOutput(7), 
      fromOutDMA(6)=>DMAOutput(6), fromOutDMA(5)=>DMAOutput(5), 
      fromOutDMA(4)=>DMAOutput(4), fromOutDMA(3)=>DMAOutput(3), 
      fromOutDMA(2)=>DMAOutput(2), fromOutDMA(1)=>DMAOutput(1), 
      fromOutDMA(0)=>DMAOutput(0), fromOutReg(15)=>RegisterOutput(15), 
      fromOutReg(14)=>RegisterOutput(14), fromOutReg(13)=>RegisterOutput(13), 
      fromOutReg(12)=>RegisterOutput(12), fromOutReg(11)=>RegisterOutput(11), 
      fromOutReg(10)=>RegisterOutput(10), fromOutReg(9)=>RegisterOutput(9), 
      fromOutReg(8)=>RegisterOutput(8), fromOutReg(7)=>RegisterOutput(7), 
      fromOutReg(6)=>RegisterOutput(6), fromOutReg(5)=>RegisterOutput(5), 
      fromOutReg(4)=>RegisterOutput(4), fromOutReg(3)=>RegisterOutput(3), 
      fromOutReg(2)=>RegisterOutput(2), fromOutReg(1)=>RegisterOutput(1), 
      fromOutReg(0)=>RegisterOutput(0), Depth(3)=>Depth(3), Depth(2)=>
      Depth(2), Depth(1)=>Depth(1), Depth(0)=>Depth(0), current_state(14)=>
      GND0, current_state(13)=>GND0, current_state(12)=>GND0, 
      current_state(11)=>GND0, current_state(10)=>GND0, current_state(9)=>
      GND0, current_state(8)=>nx238, current_state(7)=>GND0, 
      current_state(6)=>GND0, current_state(5)=>GND0, current_state(4)=>GND0, 
      current_state(3)=>GND0, current_state(2)=>GND0, current_state(1)=>GND0, 
      current_state(0)=>GND0, output(15)=>output_15_EXMPLR, output(14)=>
      output_14_EXMPLR, output(13)=>output_13_EXMPLR, output(12)=>
      output_12_EXMPLR, output(11)=>output_11_EXMPLR, output(10)=>
      output_10_EXMPLR, output(9)=>output_9_EXMPLR, output(8)=>
      output_8_EXMPLR, output(7)=>output_7_EXMPLR, output(6)=>
      output_6_EXMPLR, output(5)=>output_5_EXMPLR, output(4)=>
      output_4_EXMPLR, output(3)=>output_3_EXMPLR, output(2)=>
      output_2_EXMPLR, output(1)=>output_1_EXMPLR, output(0)=>
      output_0_EXMPLR);
   third : depthZero port map ( fromOutReg(15)=>RegisterOutput(15), 
      fromOutReg(14)=>RegisterOutput(14), fromOutReg(13)=>RegisterOutput(13), 
      fromOutReg(12)=>RegisterOutput(12), fromOutReg(11)=>RegisterOutput(11), 
      fromOutReg(10)=>RegisterOutput(10), fromOutReg(9)=>RegisterOutput(9), 
      fromOutReg(8)=>RegisterOutput(8), fromOutReg(7)=>RegisterOutput(7), 
      fromOutReg(6)=>RegisterOutput(6), fromOutReg(5)=>RegisterOutput(5), 
      fromOutReg(4)=>RegisterOutput(4), fromOutReg(3)=>RegisterOutput(3), 
      fromOutReg(2)=>RegisterOutput(2), fromOutReg(1)=>RegisterOutput(1), 
      fromOutReg(0)=>RegisterOutput(0), bias1(15)=>bias1(15), bias1(14)=>
      bias1(14), bias1(13)=>bias1(13), bias1(12)=>bias1(12), bias1(11)=>
      bias1(11), bias1(10)=>bias1(10), bias1(9)=>bias1(9), bias1(8)=>
      bias1(8), bias1(7)=>bias1(7), bias1(6)=>bias1(6), bias1(5)=>bias1(5), 
      bias1(4)=>bias1(4), bias1(3)=>bias1(3), bias1(2)=>bias1(2), bias1(1)=>
      bias1(1), bias1(0)=>bias1(0), bias2(15)=>bias2(15), bias2(14)=>
      bias2(14), bias2(13)=>bias2(13), bias2(12)=>bias2(12), bias2(11)=>
      bias2(11), bias2(10)=>bias2(10), bias2(9)=>bias2(9), bias2(8)=>
      bias2(8), bias2(7)=>bias2(7), bias2(6)=>bias2(6), bias2(5)=>bias2(5), 
      bias2(4)=>bias2(4), bias2(3)=>bias2(3), bias2(2)=>bias2(2), bias2(1)=>
      bias2(1), bias2(0)=>bias2(0), bias3(15)=>bias3(15), bias3(14)=>
      bias3(14), bias3(13)=>bias3(13), bias3(12)=>bias3(12), bias3(11)=>
      bias3(11), bias3(10)=>bias3(10), bias3(9)=>bias3(9), bias3(8)=>
      bias3(8), bias3(7)=>bias3(7), bias3(6)=>bias3(6), bias3(5)=>bias3(5), 
      bias3(4)=>bias3(4), bias3(3)=>bias3(3), bias3(2)=>bias3(2), bias3(1)=>
      bias3(1), bias3(0)=>bias3(0), bias4(15)=>bias4(15), bias4(14)=>
      bias4(14), bias4(13)=>bias4(13), bias4(12)=>bias4(12), bias4(11)=>
      bias4(11), bias4(10)=>bias4(10), bias4(9)=>bias4(9), bias4(8)=>
      bias4(8), bias4(7)=>bias4(7), bias4(6)=>bias4(6), bias4(5)=>bias4(5), 
      bias4(4)=>bias4(4), bias4(3)=>bias4(3), bias4(2)=>bias4(2), bias4(1)=>
      bias4(1), bias4(0)=>bias4(0), bias5(15)=>bias5(15), bias5(14)=>
      bias5(14), bias5(13)=>bias5(13), bias5(12)=>bias5(12), bias5(11)=>
      bias5(11), bias5(10)=>bias5(10), bias5(9)=>bias5(9), bias5(8)=>
      bias5(8), bias5(7)=>bias5(7), bias5(6)=>bias5(6), bias5(5)=>bias5(5), 
      bias5(4)=>bias5(4), bias5(3)=>bias5(3), bias5(2)=>bias5(2), bias5(1)=>
      bias5(1), bias5(0)=>bias5(0), bias6(15)=>bias6(15), bias6(14)=>
      bias6(14), bias6(13)=>bias6(13), bias6(12)=>bias6(12), bias6(11)=>
      bias6(11), bias6(10)=>bias6(10), bias6(9)=>bias6(9), bias6(8)=>
      bias6(8), bias6(7)=>bias6(7), bias6(6)=>bias6(6), bias6(5)=>bias6(5), 
      bias6(4)=>bias6(4), bias6(3)=>bias6(3), bias6(2)=>bias6(2), bias6(1)=>
      bias6(1), bias6(0)=>bias6(0), bias7(15)=>bias7(15), bias7(14)=>
      bias7(14), bias7(13)=>bias7(13), bias7(12)=>bias7(12), bias7(11)=>
      bias7(11), bias7(10)=>bias7(10), bias7(9)=>bias7(9), bias7(8)=>
      bias7(8), bias7(7)=>bias7(7), bias7(6)=>bias7(6), bias7(5)=>bias7(5), 
      bias7(4)=>bias7(4), bias7(3)=>bias7(3), bias7(2)=>bias7(2), bias7(1)=>
      bias7(1), bias7(0)=>bias7(0), bias8(15)=>bias8(15), bias8(14)=>
      bias8(14), bias8(13)=>bias8(13), bias8(12)=>bias8(12), bias8(11)=>
      bias8(11), bias8(10)=>bias8(10), bias8(9)=>bias8(9), bias8(8)=>
      bias8(8), bias8(7)=>bias8(7), bias8(6)=>bias8(6), bias8(5)=>bias8(5), 
      bias8(4)=>bias8(4), bias8(3)=>bias8(3), bias8(2)=>bias8(2), bias8(1)=>
      bias8(1), bias8(0)=>bias8(0), counterNumber(3)=>
      NumberOfFiltersCounter(3), counterNumber(2)=>NumberOfFiltersCounter(2), 
      counterNumber(1)=>NumberOfFiltersCounter(1), counterNumber(0)=>
      NumberOfFiltersCounter(0), Depth(3)=>Depth(3), Depth(2)=>Depth(2), 
      Depth(1)=>Depth(1), Depth(0)=>Depth(0), current_state(14)=>GND0, 
      current_state(13)=>GND0, current_state(12)=>GND0, current_state(11)=>
      GND0, current_state(10)=>GND0, current_state(9)=>GND0, 
      current_state(8)=>nx238, current_state(7)=>GND0, current_state(6)=>
      GND0, current_state(5)=>GND0, current_state(4)=>GND0, current_state(3)
      =>GND0, current_state(2)=>GND0, current_state(1)=>GND0, 
      current_state(0)=>GND0, output(15)=>output_15_EXMPLR, output(14)=>
      output_14_EXMPLR, output(13)=>output_13_EXMPLR, output(12)=>
      output_12_EXMPLR, output(11)=>output_11_EXMPLR, output(10)=>
      output_10_EXMPLR, output(9)=>output_9_EXMPLR, output(8)=>
      output_8_EXMPLR, output(7)=>output_7_EXMPLR, output(6)=>
      output_6_EXMPLR, output(5)=>output_5_EXMPLR, output(4)=>
      output_4_EXMPLR, output(3)=>output_3_EXMPLR, output(2)=>
      output_2_EXMPLR, output(1)=>output_1_EXMPLR, output(0)=>
      output_0_EXMPLR);
   ix214 : fake_gnd port map ( Y=>GND0);
   ix5 : or02 port map ( Y=>Enable, A0=>nx240, A1=>stateinput(10));
   ix7 : or02 port map ( Y=>resetCounter, A0=>rst, A1=>stateinput(13));
   ix3 : ao21 port map ( Y=>ShiftRegClk, A0=>clk, A1=>stateinput(10), B0=>
      nx240);
   ix237 : buf02 port map ( Y=>nx238, A=>stateinput(8));
   ix239 : buf02 port map ( Y=>nx240, A=>stateinput(8));
end saveStateArch ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Counter_4 is
   port (
      enable : IN std_logic ;
      reset : IN std_logic ;
      clk : IN std_logic ;
      load : IN std_logic ;
      output : OUT std_logic_vector (3 DOWNTO 0) ;
      input : IN std_logic_vector (3 DOWNTO 0)) ;
end Counter_4 ;

architecture CounterImplementation of Counter_4 is
   component my_nadder_4
      port (
         a : IN std_logic_vector (3 DOWNTO 0) ;
         b : IN std_logic_vector (3 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (3 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal output_3_EXMPLR, output_2_EXMPLR, output_1_EXMPLR, output_0_EXMPLR, 
      addResult_3, addResult_2, addResult_1, addResult_0, one_0, one_3, nx52, 
      NOT_clk, nx8, nx12, nx46, nx20, nx24, nx40, nx32, nx36, nx34, nx45, 
      nx49, nx143, nx153, nx163, nx173, nx182, nx216: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   output(3) <= output_3_EXMPLR ;
   output(2) <= output_2_EXMPLR ;
   output(1) <= output_1_EXMPLR ;
   output(0) <= output_0_EXMPLR ;
   A1 : my_nadder_4 port map ( a(3)=>output_3_EXMPLR, a(2)=>output_2_EXMPLR, 
      a(1)=>output_1_EXMPLR, a(0)=>output_0_EXMPLR, b(3)=>one_3, b(2)=>one_3, 
      b(1)=>one_3, b(0)=>one_0, cin=>one_3, s(3)=>addResult_3, s(2)=>
      addResult_2, s(1)=>addResult_1, s(0)=>addResult_0, cout=>DANGLING(0));
   ix120 : fake_gnd port map ( Y=>one_3);
   ix118 : fake_vcc port map ( Y=>one_0);
   reg_toOutput_0_dup_1 : dffsr_ni port map ( Q=>output_0_EXMPLR, QB=>OPEN, 
      D=>nx143, CLK=>clk, S=>nx8, R=>nx12);
   ix144 : mux21_ni port map ( Y=>nx143, A0=>output_0_EXMPLR, A1=>
      addResult_0, S0=>enable);
   ix9 : nor02ii port map ( Y=>nx8, A0=>nx182, A1=>nx52);
   ix183 : nor02_2x port map ( Y=>nx182, A0=>nx216, A1=>load);
   ix53 : dffr port map ( Q=>nx52, QB=>OPEN, D=>input(0), CLK=>NOT_clk, R=>
      nx216);
   ix186 : inv01 port map ( Y=>NOT_clk, A=>clk);
   ix13 : nor02_2x port map ( Y=>nx12, A0=>nx52, A1=>nx182);
   reg_toOutput_1_dup_1 : dffsr_ni port map ( Q=>output_1_EXMPLR, QB=>OPEN, 
      D=>nx153, CLK=>clk, S=>nx20, R=>nx24);
   ix154 : mux21_ni port map ( Y=>nx153, A0=>output_1_EXMPLR, A1=>
      addResult_1, S0=>enable);
   ix21 : nor02ii port map ( Y=>nx20, A0=>nx182, A1=>nx46);
   ix47 : dffr port map ( Q=>nx46, QB=>OPEN, D=>input(1), CLK=>NOT_clk, R=>
      nx216);
   ix25 : nor02_2x port map ( Y=>nx24, A0=>nx46, A1=>nx182);
   reg_toOutput_2_dup_1 : dffsr_ni port map ( Q=>output_2_EXMPLR, QB=>OPEN, 
      D=>nx163, CLK=>clk, S=>nx32, R=>nx36);
   ix164 : mux21_ni port map ( Y=>nx163, A0=>output_2_EXMPLR, A1=>
      addResult_2, S0=>enable);
   ix33 : nor02ii port map ( Y=>nx32, A0=>nx182, A1=>nx40);
   ix41 : dffr port map ( Q=>nx40, QB=>OPEN, D=>input(2), CLK=>NOT_clk, R=>
      nx216);
   ix37 : nor02_2x port map ( Y=>nx36, A0=>nx40, A1=>nx182);
   reg_toOutput_3_dup_1 : dffsr_ni port map ( Q=>output_3_EXMPLR, QB=>OPEN, 
      D=>nx173, CLK=>clk, S=>nx45, R=>nx49);
   ix174 : mux21_ni port map ( Y=>nx173, A0=>output_3_EXMPLR, A1=>
      addResult_3, S0=>enable);
   ix46 : nor02ii port map ( Y=>nx45, A0=>nx182, A1=>nx34);
   ix42 : dffr port map ( Q=>nx34, QB=>OPEN, D=>input(3), CLK=>NOT_clk, R=>
      nx216);
   ix50 : nor02_2x port map ( Y=>nx49, A0=>nx34, A1=>nx182);
   ix215 : buf02 port map ( Y=>nx216, A=>reset);
end CounterImplementation ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity ImageState is
   port (
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      WSquared : IN std_logic_vector (9 DOWNTO 0) ;
      AddresCounterIN : IN std_logic_vector (12 DOWNTO 0) ;
      AddresCounterLoad : OUT std_logic_vector (12 DOWNTO 0) ;
      NoOfShiftsCounter : IN std_logic_vector (4 DOWNTO 0) ;
      LayerInfoIn : IN std_logic_vector (15 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      Q : OUT std_logic ;
      NumOfFilters : OUT std_logic_vector (3 DOWNTO 0) ;
      NumOfHeight : OUT std_logic_vector (4 DOWNTO 0) ;
      X1 : OUT std_logic ;
      Y1 : OUT std_logic ;
      K1 : OUT std_logic) ;
end ImageState ;

architecture archImgState of ImageState is
   component nBitRegister_1
      port (
         D : IN std_logic_vector (0 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (0 DOWNTO 0)) ;
   end component ;
   component Counter_5
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (4 DOWNTO 0) ;
         input : IN std_logic_vector (4 DOWNTO 0)) ;
   end component ;
   component Counter_4
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (3 DOWNTO 0) ;
         input : IN std_logic_vector (3 DOWNTO 0)) ;
   end component ;
   component nBitRegister_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component my_nadder_13
      port (
         a : IN std_logic_vector (12 DOWNTO 0) ;
         b : IN std_logic_vector (12 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (12 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   signal AddresCounterLoad_12_EXMPLR, AddresCounterLoad_11_EXMPLR, 
      AddresCounterLoad_10_EXMPLR, AddresCounterLoad_9_EXMPLR, 
      AddresCounterLoad_8_EXMPLR, AddresCounterLoad_7_EXMPLR, 
      AddresCounterLoad_6_EXMPLR, AddresCounterLoad_5_EXMPLR, 
      AddresCounterLoad_4_EXMPLR, AddresCounterLoad_3_EXMPLR, 
      AddresCounterLoad_2_EXMPLR, AddresCounterLoad_1_EXMPLR, 
      AddresCounterLoad_0_EXMPLR, Q_EXMPLR, NumOfFilters_3_EXMPLR, 
      NumOfFilters_2_EXMPLR, NumOfFilters_1_EXMPLR, NumOfFilters_0_EXMPLR, 
      NumOfHeight_4_EXMPLR, NumOfHeight_3_EXMPLR, NumOfHeight_2_EXMPLR, 
      NumOfHeight_1_EXMPLR, NumOfHeight_0_EXMPLR, Qbar_0, newSliceRegOUT_12, 
      newSliceRegOUT_11, newSliceRegOUT_10, newSliceRegOUT_9, 
      newSliceRegOUT_8, newSliceRegOUT_7, newSliceRegOUT_6, newSliceRegOUT_5, 
      newSliceRegOUT_4, newSliceRegOUT_3, newSliceRegOUT_2, newSliceRegOUT_1, 
      newSliceRegOUT_0, adder0Out_12, adder0Out_11, adder0Out_10, 
      adder0Out_9, adder0Out_8, adder0Out_7, adder0Out_6, adder0Out_5, 
      adder0Out_4, adder0Out_3, adder0Out_2, adder0Out_1, adder0Out_0, 
      adder1Out_12, adder1Out_11, adder1Out_10, adder1Out_9, adder1Out_8, 
      adder1Out_7, adder1Out_6, adder1Out_5, adder1Out_4, adder1Out_3, 
      adder1Out_2, adder1Out_1, adder1Out_0, QRST, cnhRST, cnfCLK, 
      FilterCounterRst, newSliceRegRST, newSliceRegEn, triStateBuffer1EN, 
      X1_EXMPLR, Y1_EXMPLR, K1_EXMPLR, PWR, adder0b_12, YBar, nx253, nx255, 
      nx257, nx259, nx264, nx266, nx268, nx270, nx272, nx274, nx278, nx280, 
      nx282, nx284, nx286, nx288, nx295, nx297, nx300, nx310, nx316, nx318, 
      nx320, nx322, nx324: std_logic ;
   
   signal DANGLING : std_logic_vector (1 downto 0 );

begin
   AddresCounterLoad(12) <= AddresCounterLoad_12_EXMPLR ;
   AddresCounterLoad(11) <= AddresCounterLoad_11_EXMPLR ;
   AddresCounterLoad(10) <= AddresCounterLoad_10_EXMPLR ;
   AddresCounterLoad(9) <= AddresCounterLoad_9_EXMPLR ;
   AddresCounterLoad(8) <= AddresCounterLoad_8_EXMPLR ;
   AddresCounterLoad(7) <= AddresCounterLoad_7_EXMPLR ;
   AddresCounterLoad(6) <= AddresCounterLoad_6_EXMPLR ;
   AddresCounterLoad(5) <= AddresCounterLoad_5_EXMPLR ;
   AddresCounterLoad(4) <= AddresCounterLoad_4_EXMPLR ;
   AddresCounterLoad(3) <= AddresCounterLoad_3_EXMPLR ;
   AddresCounterLoad(2) <= AddresCounterLoad_2_EXMPLR ;
   AddresCounterLoad(1) <= AddresCounterLoad_1_EXMPLR ;
   AddresCounterLoad(0) <= AddresCounterLoad_0_EXMPLR ;
   Q <= Q_EXMPLR ;
   NumOfFilters(3) <= NumOfFilters_3_EXMPLR ;
   NumOfFilters(2) <= NumOfFilters_2_EXMPLR ;
   NumOfFilters(1) <= NumOfFilters_1_EXMPLR ;
   NumOfFilters(0) <= NumOfFilters_0_EXMPLR ;
   NumOfHeight(4) <= NumOfHeight_4_EXMPLR ;
   NumOfHeight(3) <= NumOfHeight_3_EXMPLR ;
   NumOfHeight(2) <= NumOfHeight_2_EXMPLR ;
   NumOfHeight(1) <= NumOfHeight_1_EXMPLR ;
   NumOfHeight(0) <= NumOfHeight_0_EXMPLR ;
   X1 <= X1_EXMPLR ;
   Y1 <= Y1_EXMPLR ;
   K1 <= K1_EXMPLR ;
   DDF0 : nBitRegister_1 port map ( D(0)=>Qbar_0, CLK=>nx310, RST=>QRST, EN
      =>PWR, Q(0)=>Q_EXMPLR);
   counterNoHeight0 : Counter_5 port map ( enable=>PWR, reset=>cnhRST, clk=>
      YBar, load=>adder0b_12, output(4)=>NumOfHeight_4_EXMPLR, output(3)=>
      NumOfHeight_3_EXMPLR, output(2)=>NumOfHeight_2_EXMPLR, output(1)=>
      NumOfHeight_1_EXMPLR, output(0)=>NumOfHeight_0_EXMPLR, input(4)=>
      adder0b_12, input(3)=>adder0b_12, input(2)=>adder0b_12, input(1)=>
      adder0b_12, input(0)=>PWR);
   counterNoFilters0 : Counter_4 port map ( enable=>PWR, reset=>
      FilterCounterRst, clk=>nx310, load=>adder0b_12, output(3)=>
      NumOfFilters_3_EXMPLR, output(2)=>NumOfFilters_2_EXMPLR, output(1)=>
      NumOfFilters_1_EXMPLR, output(0)=>NumOfFilters_0_EXMPLR, input(3)=>
      adder0b_12, input(2)=>adder0b_12, input(1)=>adder0b_12, input(0)=>PWR
   );
   newSliceReg0 : nBitRegister_13 port map ( D(12)=>adder0Out_12, D(11)=>
      adder0Out_11, D(10)=>adder0Out_10, D(9)=>adder0Out_9, D(8)=>
      adder0Out_8, D(7)=>adder0Out_7, D(6)=>adder0Out_6, D(5)=>adder0Out_5, 
      D(4)=>adder0Out_4, D(3)=>adder0Out_3, D(2)=>adder0Out_2, D(1)=>
      adder0Out_1, D(0)=>adder0Out_0, CLK=>CLK, RST=>newSliceRegRST, EN=>
      newSliceRegEn, Q(12)=>newSliceRegOUT_12, Q(11)=>newSliceRegOUT_11, 
      Q(10)=>newSliceRegOUT_10, Q(9)=>newSliceRegOUT_9, Q(8)=>
      newSliceRegOUT_8, Q(7)=>newSliceRegOUT_7, Q(6)=>newSliceRegOUT_6, Q(5)
      =>newSliceRegOUT_5, Q(4)=>newSliceRegOUT_4, Q(3)=>newSliceRegOUT_3, 
      Q(2)=>newSliceRegOUT_2, Q(1)=>newSliceRegOUT_1, Q(0)=>newSliceRegOUT_0
   );
   adder0 : my_nadder_13 port map ( a(12)=>newSliceRegOUT_12, a(11)=>
      newSliceRegOUT_11, a(10)=>newSliceRegOUT_10, a(9)=>newSliceRegOUT_9, 
      a(8)=>newSliceRegOUT_8, a(7)=>newSliceRegOUT_7, a(6)=>newSliceRegOUT_6, 
      a(5)=>newSliceRegOUT_5, a(4)=>newSliceRegOUT_4, a(3)=>newSliceRegOUT_3, 
      a(2)=>newSliceRegOUT_2, a(1)=>newSliceRegOUT_1, a(0)=>newSliceRegOUT_0, 
      b(12)=>adder0b_12, b(11)=>adder0b_12, b(10)=>adder0b_12, b(9)=>
      adder0b_12, b(8)=>adder0b_12, b(7)=>adder0b_12, b(6)=>adder0b_12, b(5)
      =>adder0b_12, b(4)=>nx316, b(3)=>nx318, b(2)=>nx320, b(1)=>nx322, b(0)
      =>nx324, cin=>adder0b_12, s(12)=>adder0Out_12, s(11)=>adder0Out_11, 
      s(10)=>adder0Out_10, s(9)=>adder0Out_9, s(8)=>adder0Out_8, s(7)=>
      adder0Out_7, s(6)=>adder0Out_6, s(5)=>adder0Out_5, s(4)=>adder0Out_4, 
      s(3)=>adder0Out_3, s(2)=>adder0Out_2, s(1)=>adder0Out_1, s(0)=>
      adder0Out_0, cout=>DANGLING(0));
   triStateBuffer0 : triStateBuffer_13 port map ( D(12)=>adder0Out_12, D(11)
      =>adder0Out_11, D(10)=>adder0Out_10, D(9)=>adder0Out_9, D(8)=>
      adder0Out_8, D(7)=>adder0Out_7, D(6)=>adder0Out_6, D(5)=>adder0Out_5, 
      D(4)=>adder0Out_4, D(3)=>adder0Out_3, D(2)=>adder0Out_2, D(1)=>
      adder0Out_1, D(0)=>adder0Out_0, EN=>newSliceRegEn, F(12)=>
      AddresCounterLoad_12_EXMPLR, F(11)=>AddresCounterLoad_11_EXMPLR, F(10)
      =>AddresCounterLoad_10_EXMPLR, F(9)=>AddresCounterLoad_9_EXMPLR, F(8)
      =>AddresCounterLoad_8_EXMPLR, F(7)=>AddresCounterLoad_7_EXMPLR, F(6)=>
      AddresCounterLoad_6_EXMPLR, F(5)=>AddresCounterLoad_5_EXMPLR, F(4)=>
      AddresCounterLoad_4_EXMPLR, F(3)=>AddresCounterLoad_3_EXMPLR, F(2)=>
      AddresCounterLoad_2_EXMPLR, F(1)=>AddresCounterLoad_1_EXMPLR, F(0)=>
      AddresCounterLoad_0_EXMPLR);
   adder1 : my_nadder_13 port map ( a(12)=>AddresCounterIN(12), a(11)=>
      AddresCounterIN(11), a(10)=>AddresCounterIN(10), a(9)=>
      AddresCounterIN(9), a(8)=>AddresCounterIN(8), a(7)=>AddresCounterIN(7), 
      a(6)=>AddresCounterIN(6), a(5)=>AddresCounterIN(5), a(4)=>
      AddresCounterIN(4), a(3)=>AddresCounterIN(3), a(2)=>AddresCounterIN(2), 
      a(1)=>AddresCounterIN(1), a(0)=>AddresCounterIN(0), b(12)=>adder0b_12, 
      b(11)=>adder0b_12, b(10)=>adder0b_12, b(9)=>WSquared(9), b(8)=>
      WSquared(8), b(7)=>WSquared(7), b(6)=>WSquared(6), b(5)=>WSquared(5), 
      b(4)=>WSquared(4), b(3)=>WSquared(3), b(2)=>WSquared(2), b(1)=>
      WSquared(1), b(0)=>WSquared(0), cin=>adder0b_12, s(12)=>adder1Out_12, 
      s(11)=>adder1Out_11, s(10)=>adder1Out_10, s(9)=>adder1Out_9, s(8)=>
      adder1Out_8, s(7)=>adder1Out_7, s(6)=>adder1Out_6, s(5)=>adder1Out_5, 
      s(4)=>adder1Out_4, s(3)=>adder1Out_3, s(2)=>adder1Out_2, s(1)=>
      adder1Out_1, s(0)=>adder1Out_0, cout=>DANGLING(1));
   triStateBuffer1 : triStateBuffer_13 port map ( D(12)=>adder1Out_12, D(11)
      =>adder1Out_11, D(10)=>adder1Out_10, D(9)=>adder1Out_9, D(8)=>
      adder1Out_8, D(7)=>adder1Out_7, D(6)=>adder1Out_6, D(5)=>adder1Out_5, 
      D(4)=>adder1Out_4, D(3)=>adder1Out_3, D(2)=>adder1Out_2, D(1)=>
      adder1Out_1, D(0)=>adder1Out_0, EN=>triStateBuffer1EN, F(12)=>
      AddresCounterLoad_12_EXMPLR, F(11)=>AddresCounterLoad_11_EXMPLR, F(10)
      =>AddresCounterLoad_10_EXMPLR, F(9)=>AddresCounterLoad_9_EXMPLR, F(8)
      =>AddresCounterLoad_8_EXMPLR, F(7)=>AddresCounterLoad_7_EXMPLR, F(6)=>
      AddresCounterLoad_6_EXMPLR, F(5)=>AddresCounterLoad_5_EXMPLR, F(4)=>
      AddresCounterLoad_4_EXMPLR, F(3)=>AddresCounterLoad_3_EXMPLR, F(2)=>
      AddresCounterLoad_2_EXMPLR, F(1)=>AddresCounterLoad_1_EXMPLR, F(0)=>
      AddresCounterLoad_0_EXMPLR);
   ix254 : xnor2 port map ( Y=>nx253, A0=>LayerInfoIn(3), A1=>
      NumOfFilters_3_EXMPLR);
   ix256 : xnor2 port map ( Y=>nx255, A0=>LayerInfoIn(2), A1=>
      NumOfFilters_2_EXMPLR);
   ix258 : xnor2 port map ( Y=>nx257, A0=>LayerInfoIn(1), A1=>
      NumOfFilters_1_EXMPLR);
   ix260 : xnor2 port map ( Y=>nx259, A0=>LayerInfoIn(0), A1=>
      NumOfFilters_0_EXMPLR);
   ix221 : fake_gnd port map ( Y=>adder0b_12);
   ix219 : fake_vcc port map ( Y=>PWR);
   ix17 : nand04 port map ( Y=>K1_EXMPLR, A0=>nx264, A1=>nx270, A2=>nx272, 
      A3=>nx274);
   ix265 : and02 port map ( Y=>nx264, A0=>nx266, A1=>nx268);
   ix267 : xnor2 port map ( Y=>nx266, A0=>nx318, A1=>NumOfHeight_3_EXMPLR);
   ix269 : xnor2 port map ( Y=>nx268, A0=>nx320, A1=>NumOfHeight_2_EXMPLR);
   ix271 : xnor2 port map ( Y=>nx270, A0=>nx324, A1=>NumOfHeight_0_EXMPLR);
   ix273 : xnor2 port map ( Y=>nx272, A0=>nx316, A1=>NumOfHeight_4_EXMPLR);
   ix275 : xnor2 port map ( Y=>nx274, A0=>nx322, A1=>NumOfHeight_1_EXMPLR);
   ix49 : nand04 port map ( Y=>Y1_EXMPLR, A0=>nx253, A1=>nx255, A2=>nx257, 
      A3=>nx259);
   ix35 : nand04 port map ( Y=>X1_EXMPLR, A0=>nx278, A1=>nx284, A2=>nx286, 
      A3=>nx288);
   ix279 : and02 port map ( Y=>nx278, A0=>nx280, A1=>nx282);
   ix281 : xnor2 port map ( Y=>nx280, A0=>nx318, A1=>NoOfShiftsCounter(3));
   ix283 : xnor2 port map ( Y=>nx282, A0=>nx320, A1=>NoOfShiftsCounter(2));
   ix285 : xnor2 port map ( Y=>nx284, A0=>nx324, A1=>NoOfShiftsCounter(0));
   ix287 : xnor2 port map ( Y=>nx286, A0=>nx316, A1=>NoOfShiftsCounter(4));
   ix289 : xnor2 port map ( Y=>nx288, A0=>nx322, A1=>NoOfShiftsCounter(1));
   ix61 : nor02ii port map ( Y=>triStateBuffer1EN, A0=>newSliceRegEn, A1=>
      nx310);
   ix53 : nor02ii port map ( Y=>newSliceRegEn, A0=>Y1_EXMPLR, A1=>
      current_state(9));
   ix57 : nor02ii port map ( Y=>cnfCLK, A0=>X1_EXMPLR, A1=>current_state(9)
   );
   ix63 : or02 port map ( Y=>newSliceRegRST, A0=>RST, A1=>current_state(12)
   );
   ix69 : oai21 port map ( Y=>FilterCounterRst, A0=>nx295, A1=>Y1_EXMPLR, B0
      =>nx297);
   ix296 : inv01 port map ( Y=>nx295, A=>current_state(11));
   ix298 : inv01 port map ( Y=>nx297, A=>RST);
   ix77 : oai21 port map ( Y=>cnhRST, A0=>nx300, A1=>K1_EXMPLR, B0=>nx297);
   ix301 : inv01 port map ( Y=>nx300, A=>current_state(12));
   ix79 : or02 port map ( Y=>QRST, A0=>RST, A1=>current_state(13));
   ix304 : inv01 port map ( Y=>Qbar_0, A=>Q_EXMPLR);
   ix252 : inv01 port map ( Y=>YBar, A=>Y1_EXMPLR);
   ix309 : buf02 port map ( Y=>nx310, A=>cnfCLK);
   ix315 : buf02 port map ( Y=>nx316, A=>LayerInfoIn(8));
   ix317 : buf02 port map ( Y=>nx318, A=>LayerInfoIn(7));
   ix319 : buf02 port map ( Y=>nx320, A=>LayerInfoIn(6));
   ix321 : buf02 port map ( Y=>nx322, A=>LayerInfoIn(5));
   ix323 : buf02 port map ( Y=>nx324, A=>LayerInfoIn(4));
end archImgState ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity StateChecks is
   port (
      current_state : IN std_logic_vector (14 DOWNTO 0) ;
      noOfLayers : IN std_logic_vector (15 DOWNTO 0) ;
      LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
      CLK : IN std_logic ;
      RST : IN std_logic ;
      L : OUT std_logic ;
      D : OUT std_logic ;
      CNDoutput : OUT std_logic_vector (3 DOWNTO 0) ;
      CNLoutput : OUT std_logic_vector (1 DOWNTO 0)) ;
end StateChecks ;

architecture archCHECKS of StateChecks is
   component Counter_4
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (3 DOWNTO 0) ;
         input : IN std_logic_vector (3 DOWNTO 0)) ;
   end component ;
   component Counter_2
      port (
         enable : IN std_logic ;
         reset : IN std_logic ;
         clk : IN std_logic ;
         load : IN std_logic ;
         output : OUT std_logic_vector (1 DOWNTO 0) ;
         input : IN std_logic_vector (1 DOWNTO 0)) ;
   end component ;
   signal CNDoutput_3_EXMPLR, CNDoutput_2_EXMPLR, CNDoutput_1_EXMPLR, 
      CNDoutput_0_EXMPLR, CNLoutput_1_EXMPLR, CNLoutput_0_EXMPLR, 
      DepthCounterRst, SDbar, D_EXMPLR, GND0, PWR, nx62, nx64, nx67, nx69, 
      nx71, nx73: std_logic ;

begin
   D <= D_EXMPLR ;
   CNDoutput(3) <= CNDoutput_3_EXMPLR ;
   CNDoutput(2) <= CNDoutput_2_EXMPLR ;
   CNDoutput(1) <= CNDoutput_1_EXMPLR ;
   CNDoutput(0) <= CNDoutput_0_EXMPLR ;
   CNLoutput(1) <= CNLoutput_1_EXMPLR ;
   CNLoutput(0) <= CNLoutput_0_EXMPLR ;
   counterNoDepth0 : Counter_4 port map ( enable=>PWR, reset=>
      DepthCounterRst, clk=>current_state(12), load=>GND0, output(3)=>
      CNDoutput_3_EXMPLR, output(2)=>CNDoutput_2_EXMPLR, output(1)=>
      CNDoutput_1_EXMPLR, output(0)=>CNDoutput_0_EXMPLR, input(3)=>GND0, 
      input(2)=>GND0, input(1)=>GND0, input(0)=>PWR);
   counterNoLayer0 : Counter_2 port map ( enable=>PWR, reset=>RST, clk=>
      SDbar, load=>GND0, output(1)=>CNLoutput_1_EXMPLR, output(0)=>
      CNLoutput_0_EXMPLR, input(1)=>GND0, input(0)=>PWR);
   ix44 : fake_vcc port map ( Y=>PWR);
   ix42 : fake_gnd port map ( Y=>GND0);
   ix5 : nand02 port map ( Y=>L, A0=>nx62, A1=>nx64);
   ix63 : xnor2 port map ( Y=>nx62, A0=>CNLoutput_1_EXMPLR, A1=>
      noOfLayers(1));
   ix65 : xnor2 port map ( Y=>nx64, A0=>CNLoutput_0_EXMPLR, A1=>
      noOfLayers(0));
   ix19 : nand04 port map ( Y=>D_EXMPLR, A0=>nx67, A1=>nx69, A2=>nx71, A3=>
      nx73);
   ix68 : xnor2 port map ( Y=>nx67, A0=>CNDoutput_3_EXMPLR, A1=>
      LayerInfo(12));
   ix70 : xnor2 port map ( Y=>nx69, A0=>CNDoutput_2_EXMPLR, A1=>
      LayerInfo(11));
   ix72 : xnor2 port map ( Y=>nx71, A0=>CNDoutput_1_EXMPLR, A1=>
      LayerInfo(10));
   ix74 : xnor2 port map ( Y=>nx73, A0=>CNDoutput_0_EXMPLR, A1=>LayerInfo(9)
   );
   ix23 : or02 port map ( Y=>DepthCounterRst, A0=>RST, A1=>current_state(13)
   );
   ix76 : inv01 port map ( Y=>SDbar, A=>D_EXMPLR);
end archCHECKS ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity outWidthState is
   port (
      currentState : IN std_logic_vector (14 DOWNTO 0) ;
      infoReg : IN std_logic_vector (15 DOWNTO 0) ;
      address : OUT std_logic_vector (12 DOWNTO 0) ;
      outWidth : OUT std_logic_vector (15 DOWNTO 0)) ;
end outWidthState ;

architecture archOutWidthState of outWidthState is
   signal nx263, nx268, nx271, nx274, nx277, nx280, nx311, nx313, nx315, 
      nx317, nx319, nx321: std_logic ;

begin
   ix264 : fake_vcc port map ( Y=>nx263);
   tri_outwidthbefore_0 : tri01 port map ( Y=>outWidth(0), A=>nx268, E=>
      nx313);
   ix269 : inv01 port map ( Y=>nx268, A=>infoReg(4));
   tri_outwidthbefore_1 : tri01 port map ( Y=>outWidth(1), A=>nx271, E=>
      nx313);
   ix272 : inv01 port map ( Y=>nx271, A=>infoReg(5));
   tri_outwidthbefore_2 : tri01 port map ( Y=>outWidth(2), A=>nx274, E=>
      nx313);
   ix275 : inv01 port map ( Y=>nx274, A=>infoReg(6));
   tri_outwidthbefore_3 : tri01 port map ( Y=>outWidth(3), A=>nx277, E=>
      nx313);
   ix278 : inv01 port map ( Y=>nx277, A=>infoReg(7));
   tri_outwidthbefore_4 : tri01 port map ( Y=>outWidth(4), A=>nx280, E=>
      nx313);
   ix281 : inv01 port map ( Y=>nx280, A=>infoReg(8));
   tri_outwidthbefore_5 : tri01 port map ( Y=>outWidth(5), A=>nx263, E=>
      nx313);
   tri_outwidthbefore_6 : tri01 port map ( Y=>outWidth(6), A=>nx263, E=>
      nx313);
   tri_outwidthbefore_7 : tri01 port map ( Y=>outWidth(7), A=>nx263, E=>
      nx315);
   tri_outwidthbefore_8 : tri01 port map ( Y=>outWidth(8), A=>nx263, E=>
      nx315);
   tri_outwidthbefore_9 : tri01 port map ( Y=>outWidth(9), A=>nx263, E=>
      nx315);
   tri_outwidthbefore_10 : tri01 port map ( Y=>outWidth(10), A=>nx263, E=>
      nx315);
   tri_outwidthbefore_11 : tri01 port map ( Y=>outWidth(11), A=>nx263, E=>
      nx315);
   tri_outwidthbefore_12 : tri01 port map ( Y=>outWidth(12), A=>nx263, E=>
      nx315);
   tri_outwidthbefore_13 : tri01 port map ( Y=>outWidth(13), A=>nx263, E=>
      nx315);
   tri_outwidthbefore_14 : tri01 port map ( Y=>outWidth(14), A=>nx263, E=>
      nx317);
   tri_outwidthbefore_15 : tri01 port map ( Y=>outWidth(15), A=>nx263, E=>
      nx317);
   tri_address_0 : tri01 port map ( Y=>address(0), A=>nx263, E=>nx317);
   tri_address_1 : tri01 port map ( Y=>address(1), A=>nx263, E=>nx317);
   tri_address_2 : tri01 port map ( Y=>address(2), A=>nx263, E=>nx317);
   tri_address_3 : tri01 port map ( Y=>address(3), A=>nx263, E=>nx317);
   tri_address_4 : tri01 port map ( Y=>address(4), A=>nx263, E=>nx317);
   tri_address_5 : tri01 port map ( Y=>address(5), A=>nx263, E=>nx319);
   tri_address_6 : tri01 port map ( Y=>address(6), A=>nx263, E=>nx319);
   tri_address_7 : tri01 port map ( Y=>address(7), A=>nx263, E=>nx319);
   tri_address_8 : tri01 port map ( Y=>address(8), A=>nx263, E=>nx319);
   tri_address_9 : tri01 port map ( Y=>address(9), A=>nx263, E=>nx319);
   tri_address_10 : tri01 port map ( Y=>address(10), A=>nx263, E=>nx319);
   tri_address_11 : tri01 port map ( Y=>address(11), A=>nx263, E=>nx319);
   tri_address_12 : tri01 port map ( Y=>address(12), A=>nx263, E=>nx321);
   ix310 : inv01 port map ( Y=>nx311, A=>currentState(13));
   ix312 : inv01 port map ( Y=>nx313, A=>nx311);
   ix314 : inv01 port map ( Y=>nx315, A=>nx311);
   ix316 : inv01 port map ( Y=>nx317, A=>nx311);
   ix318 : inv01 port map ( Y=>nx319, A=>nx311);
   ix320 : inv01 port map ( Y=>nx321, A=>nx311);
end archOutWidthState ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity Main is
   port (
      rst : IN std_logic ;
      cl : IN std_logic ;
      start : IN std_logic ;
      dmaStartSignal : INOUT std_logic ;
      done : OUT std_logic) ;
end Main ;

architecture vlsi of Main is
   component nBitRegister_1
      port (
         D : IN std_logic_vector (0 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (0 DOWNTO 0)) ;
   end component ;
   component triStateBuffer_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         EN : IN std_logic ;
         F : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component nBitRegister_13
      port (
         D : IN std_logic_vector (12 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         EN : IN std_logic ;
         Q : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component RAM_25
      port (
         reset : IN std_logic ;
         CLK : IN std_logic ;
         W : IN std_logic ;
         R : IN std_logic ;
         address : IN std_logic_vector (12 DOWNTO 0) ;
         dataIn : IN std_logic_vector (15 DOWNTO 0) ;
         dataOut : OUT std_logic_vector (399 DOWNTO 0) ;
         MFC : OUT std_logic ;
         counterOut : OUT std_logic_vector (3 DOWNTO 0)) ;
   end component ;
   component memoryDMA
      port (
         resetEN : IN std_logic ;
         AddressIn : IN std_logic_vector (12 DOWNTO 0) ;
         dataIn : IN std_logic_vector (15 DOWNTO 0) ;
         switcherEN : IN std_logic ;
         ramSelector : IN std_logic ;
         readEn : IN std_logic ;
         writeEn : IN std_logic ;
         CLK : IN std_logic ;
         Normal : IN std_logic ;
         MFC : OUT std_logic ;
         counterOut : OUT std_logic_vector (3 DOWNTO 0) ;
         dataOut : OUT std_logic_vector (447 DOWNTO 0)) ;
   end component ;
   component ReadInfoState
      port (
         CLK : IN std_logic ;
         S : IN std_logic_vector (14 DOWNTO 0) ;
         reset : IN std_logic ;
         MFC : IN std_logic ;
         filterAddressReg_out : IN std_logic_vector (12 DOWNTO 0) ;
         filterRamData : IN std_logic_vector (15 DOWNTO 0) ;
         noOfLayersReg_out : OUT std_logic_vector (15 DOWNTO 0) ;
         filterRamAddress : OUT std_logic_vector (12 DOWNTO 0)) ;
   
   end component ;
   component my_nadder_13
      port (
         a : IN std_logic_vector (12 DOWNTO 0) ;
         b : IN std_logic_vector (12 DOWNTO 0) ;
         cin : IN std_logic ;
         s : OUT std_logic_vector (12 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   component ReadLayerInfo
      port (
         LayerInfoIn : IN std_logic_vector (15 DOWNTO 0) ;
         ImgWidthIn : IN std_logic_vector (15 DOWNTO 0) ;
         FilterAdd : IN std_logic_vector (12 DOWNTO 0) ;
         ImgAdd : IN std_logic_vector (12 DOWNTO 0) ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         ACKF : IN std_logic ;
         ACKI : IN std_logic ;
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         LayerInfoOut : OUT std_logic_vector (15 DOWNTO 0) ;
         ImgWidthOut : OUT std_logic_vector (15 DOWNTO 0) ;
         FilterAddToDMA : OUT std_logic_vector (12 DOWNTO 0) ;
         ImgAddToDMA : OUT std_logic_vector (12 DOWNTO 0)) ;
   end component ;
   component CalculateInfo
      port (
         WSquareOut : OUT std_logic_vector (9 DOWNTO 0) ;
         CounOut : OUT std_logic_vector (1 DOWNTO 0) ;
         LayerInfoIn : IN std_logic_vector (15 DOWNTO 0) ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         ACK : OUT std_logic ;
         ACKI : IN std_logic ;
         Wmin1 : OUT std_logic_vector (4 DOWNTO 0)) ;
   end component ;
   component ReadBias
      port (
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         BIAS : IN std_logic_vector (399 DOWNTO 0) ;
         FilterAddress : IN std_logic_vector (12 DOWNTO 0) ;
         DMAAddressToFilter : OUT std_logic_vector (12 DOWNTO 0) ;
         UpdatedAddress : OUT std_logic_vector (12 DOWNTO 0) ;
         changerAdd : OUT std_logic_vector (12 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
         outBias0 : OUT std_logic_vector (15 DOWNTO 0) ;
         outBias1 : OUT std_logic_vector (15 DOWNTO 0) ;
         outBias2 : OUT std_logic_vector (15 DOWNTO 0) ;
         outBias3 : OUT std_logic_vector (15 DOWNTO 0) ;
         outBias4 : OUT std_logic_vector (15 DOWNTO 0) ;
         outBias5 : OUT std_logic_vector (15 DOWNTO 0) ;
         outBias6 : OUT std_logic_vector (15 DOWNTO 0) ;
         outBias7 : OUT std_logic_vector (15 DOWNTO 0) ;
         ACKF : IN std_logic) ;
   end component ;
   component ReadFilter
      port (
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
         depthcounter : IN std_logic_vector (3 DOWNTO 0) ;
         FilterCounter : IN std_logic_vector (3 DOWNTO 0) ;
         Heightcounter : IN std_logic_vector (4 DOWNTO 0) ;
         FILTER : IN std_logic_vector (399 DOWNTO 0) ;
         FilterAddress : IN std_logic_vector (12 DOWNTO 0) ;
         msbNoOfFilters : IN std_logic ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         QImgStat : IN std_logic ;
         ACKF : IN std_logic ;
         IndicatorFilter : OUT std_logic_vector (0 DOWNTO 0) ;
         DMAAddress : OUT std_logic_vector (12 DOWNTO 0) ;
         UpdatedAddress : OUT std_logic_vector (12 DOWNTO 0) ;
         outFilter0 : OUT std_logic_vector (399 DOWNTO 0) ;
         outFilter1 : OUT std_logic_vector (399 DOWNTO 0) ;
         donttrust : OUT std_logic ;
         LastFilterIND : OUT std_logic ;
         LastHeightOut : OUT std_logic ;
         lastDepthOut : OUT std_logic) ;
   end component ;
   component ReadImage
      port (
         WI : IN std_logic ;
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         ACK : IN std_logic ;
         ImgAddress : IN std_logic_vector (12 DOWNTO 0) ;
         ImgWidth : IN std_logic_vector (15 DOWNTO 0) ;
         DATA : IN std_logic_vector (447 DOWNTO 0) ;
         OutputImg0 : OUT std_logic_vector (447 DOWNTO 0) ;
         OutputImg1 : OUT std_logic_vector (447 DOWNTO 0) ;
         OutputImg2 : OUT std_logic_vector (447 DOWNTO 0) ;
         OutputImg3 : OUT std_logic_vector (447 DOWNTO 0) ;
         OutputImg4 : OUT std_logic_vector (447 DOWNTO 0) ;
         OutputImg5 : OUT std_logic_vector (447 DOWNTO 0) ;
         ImgCounterOuput : OUT std_logic_vector (2 DOWNTO 0) ;
         ImgAddToDma : OUT std_logic_vector (12 DOWNTO 0) ;
         UpdatedAddress : OUT std_logic_vector (12 DOWNTO 0) ;
         ImgIndic : OUT std_logic_vector (0 DOWNTO 0) ;
         ImgEn : OUT std_logic_vector (5 DOWNTO 0) ;
         dontTrust : IN std_logic) ;
   end component ;
   component Convolution
      port (
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         QImgStat : IN std_logic ;
         ACK : OUT std_logic ;
         LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
         ImgAddress : IN std_logic_vector (12 DOWNTO 0) ;
         OutputImg0 : IN std_logic_vector (79 DOWNTO 0) ;
         OutputImg1 : IN std_logic_vector (79 DOWNTO 0) ;
         OutputImg2 : IN std_logic_vector (79 DOWNTO 0) ;
         OutputImg3 : IN std_logic_vector (79 DOWNTO 0) ;
         OutputImg4 : IN std_logic_vector (79 DOWNTO 0) ;
         outFilter0 : IN std_logic_vector (399 DOWNTO 0) ;
         outFilter1 : IN std_logic_vector (399 DOWNTO 0) ;
         ConvOuput : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   component saveState
      port (
         DMAOutput : IN std_logic_vector (15 DOWNTO 0) ;
         RegisterOutput : IN std_logic_vector (15 DOWNTO 0) ;
         bias1 : IN std_logic_vector (15 DOWNTO 0) ;
         bias2 : IN std_logic_vector (15 DOWNTO 0) ;
         bias3 : IN std_logic_vector (15 DOWNTO 0) ;
         bias4 : IN std_logic_vector (15 DOWNTO 0) ;
         bias5 : IN std_logic_vector (15 DOWNTO 0) ;
         bias6 : IN std_logic_vector (15 DOWNTO 0) ;
         bias7 : IN std_logic_vector (15 DOWNTO 0) ;
         bias8 : IN std_logic_vector (15 DOWNTO 0) ;
         Depth : IN std_logic_vector (3 DOWNTO 0) ;
         NumberOfFiltersCounter : IN std_logic_vector (3 DOWNTO 0) ;
         rst : IN std_logic ;
         stateinput : IN std_logic_vector (14 DOWNTO 0) ;
         clk : IN std_logic ;
         outputCounterToDma : OUT std_logic_vector (12 DOWNTO 0) ;
         RealOutputCounter : OUT std_logic_vector (12 DOWNTO 0) ;
         output : OUT std_logic_vector (15 DOWNTO 0) ;
         ShiftLeftCounterOutput : OUT std_logic_vector (4 DOWNTO 0) ;
         ShiftCounterRst : IN std_logic ;
         AddresCounterLoad : IN std_logic_vector (12 DOWNTO 0) ;
         X : IN std_logic ;
         Y : IN std_logic) ;
   end component ;
   component ImageState
      port (
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         WSquared : IN std_logic_vector (9 DOWNTO 0) ;
         AddresCounterIN : IN std_logic_vector (12 DOWNTO 0) ;
         AddresCounterLoad : OUT std_logic_vector (12 DOWNTO 0) ;
         NoOfShiftsCounter : IN std_logic_vector (4 DOWNTO 0) ;
         LayerInfoIn : IN std_logic_vector (15 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         Q : OUT std_logic ;
         NumOfFilters : OUT std_logic_vector (3 DOWNTO 0) ;
         NumOfHeight : OUT std_logic_vector (4 DOWNTO 0) ;
         X1 : OUT std_logic ;
         Y1 : OUT std_logic ;
         K1 : OUT std_logic) ;
   end component ;
   component StateChecks
      port (
         current_state : IN std_logic_vector (14 DOWNTO 0) ;
         noOfLayers : IN std_logic_vector (15 DOWNTO 0) ;
         LayerInfo : IN std_logic_vector (15 DOWNTO 0) ;
         CLK : IN std_logic ;
         RST : IN std_logic ;
         L : OUT std_logic ;
         D : OUT std_logic ;
         CNDoutput : OUT std_logic_vector (3 DOWNTO 0) ;
         CNLoutput : OUT std_logic_vector (1 DOWNTO 0)) ;
   end component ;
   component outWidthState
      port (
         currentState : IN std_logic_vector (14 DOWNTO 0) ;
         infoReg : IN std_logic_vector (15 DOWNTO 0) ;
         address : OUT std_logic_vector (12 DOWNTO 0) ;
         outWidth : OUT std_logic_vector (15 DOWNTO 0)) ;
   end component ;
   signal done_EXMPLR, current_state_11, current_state_10, current_state_9, 
      current_state_8, current_state_6, current_state_5, current_state_4, 
      current_state_3, current_state_2, current_state_0, FilterAddressIN_12, 
      FilterAddressIN_11, FilterAddressIN_10, FilterAddressIN_9, 
      FilterAddressIN_8, FilterAddressIN_7, FilterAddressIN_6, 
      FilterAddressIN_5, FilterAddressIN_4, FilterAddressIN_3, 
      FilterAddressIN_2, FilterAddressIN_1, FilterAddressIN_0, 
      FilterAddressOut_12, FilterAddressOut_11, FilterAddressOut_10, 
      FilterAddressOut_9, FilterAddressOut_8, FilterAddressOut_7, 
      FilterAddressOut_6, FilterAddressOut_5, FilterAddressOut_4, 
      FilterAddressOut_3, FilterAddressOut_2, FilterAddressOut_1, 
      FilterAddressOut_0, AddressChangerIN_12, AddressChangerIN_11, 
      AddressChangerIN_10, AddressChangerIN_9, AddressChangerIN_8, 
      AddressChangerIN_7, AddressChangerIN_6, AddressChangerIN_5, 
      AddressChangerIN_4, AddressChangerIN_3, AddressChangerIN_2, 
      AddressChangerIN_1, AddressChangerIN_0, AddressChangerOut_12, 
      AddressChangerOut_11, AddressChangerOut_10, AddressChangerOut_9, 
      AddressChangerOut_8, AddressChangerOut_7, AddressChangerOut_6, 
      AddressChangerOut_5, AddressChangerOut_4, AddressChangerOut_3, 
      AddressChangerOut_2, AddressChangerOut_1, AddressChangerOut_0, 
      ImgAddRegIN_12, ImgAddRegIN_11, ImgAddRegIN_10, ImgAddRegIN_9, 
      ImgAddRegIN_8, ImgAddRegIN_7, ImgAddRegIN_6, ImgAddRegIN_5, 
      ImgAddRegIN_4, ImgAddRegIN_3, ImgAddRegIN_2, ImgAddRegIN_1, 
      ImgAddRegIN_0, ImgAddRegOut_12, ImgAddRegOut_11, ImgAddRegOut_10, 
      ImgAddRegOut_9, ImgAddRegOut_8, ImgAddRegOut_7, ImgAddRegOut_6, 
      ImgAddRegOut_5, ImgAddRegOut_4, ImgAddRegOut_3, ImgAddRegOut_2, 
      ImgAddRegOut_1, ImgAddRegOut_0, TriStateCounterOUT_12, 
      TriStateCounterOUT_11, TriStateCounterOUT_10, TriStateCounterOUT_9, 
      TriStateCounterOUT_8, TriStateCounterOUT_7, TriStateCounterOUT_6, 
      TriStateCounterOUT_5, TriStateCounterOUT_4, TriStateCounterOUT_3, 
      TriStateCounterOUT_2, TriStateCounterOUT_1, TriStateCounterOUT_0, 
      ImgAddACKTriIN_0, ReadF, AddressF_12, AddressF_11, AddressF_10, 
      AddressF_9, AddressF_8, AddressF_7, AddressF_6, AddressF_5, AddressF_4, 
      AddressF_3, AddressF_2, AddressF_1, AddressF_0, DataFOut_399, ACKF, 
      WriteI, ReadI, AddressI_12, AddressI_11, AddressI_10, AddressI_9, 
      AddressI_8, AddressI_7, AddressI_6, AddressI_5, AddressI_4, AddressI_3, 
      AddressI_2, AddressI_1, AddressI_0, DataIIn_15, DataIIn_14, DataIIn_13, 
      DataIIn_12, DataIIn_11, DataIIn_10, DataIIn_9, DataIIn_8, DataIIn_7, 
      DataIIn_6, DataIIn_5, DataIIn_4, DataIIn_3, DataIIn_2, DataIIn_1, 
      DataIIn_0, DataIOut_447, DataIOut_446, DataIOut_445, DataIOut_444, 
      DataIOut_443, DataIOut_442, DataIOut_441, DataIOut_440, DataIOut_439, 
      DataIOut_438, DataIOut_437, DataIOut_436, DataIOut_435, DataIOut_434, 
      DataIOut_433, DataIOut_432, DataIOut_431, DataIOut_430, DataIOut_429, 
      DataIOut_428, DataIOut_427, DataIOut_426, DataIOut_425, DataIOut_424, 
      DataIOut_423, DataIOut_422, DataIOut_421, DataIOut_420, DataIOut_419, 
      DataIOut_418, DataIOut_417, DataIOut_416, DataIOut_415, DataIOut_414, 
      DataIOut_413, DataIOut_412, DataIOut_411, DataIOut_410, DataIOut_409, 
      DataIOut_408, DataIOut_407, DataIOut_406, DataIOut_405, DataIOut_404, 
      DataIOut_403, DataIOut_402, DataIOut_401, DataIOut_400, DataIOut_399, 
      DataIOut_398, DataIOut_397, DataIOut_396, DataIOut_395, DataIOut_394, 
      DataIOut_393, DataIOut_392, DataIOut_391, DataIOut_390, DataIOut_389, 
      DataIOut_388, DataIOut_387, DataIOut_386, DataIOut_385, DataIOut_384, 
      DataIOut_383, DataIOut_382, DataIOut_381, DataIOut_380, DataIOut_379, 
      DataIOut_378, DataIOut_377, DataIOut_376, DataIOut_375, DataIOut_374, 
      DataIOut_373, DataIOut_372, DataIOut_371, DataIOut_370, DataIOut_369, 
      DataIOut_368, DataIOut_367, DataIOut_366, DataIOut_365, DataIOut_364, 
      DataIOut_363, DataIOut_362, DataIOut_361, DataIOut_360, DataIOut_359, 
      DataIOut_358, DataIOut_357, DataIOut_356, DataIOut_355, DataIOut_354, 
      DataIOut_353, DataIOut_352, DataIOut_351, DataIOut_350, DataIOut_349, 
      DataIOut_348, DataIOut_347, DataIOut_346, DataIOut_345, DataIOut_344, 
      DataIOut_343, DataIOut_342, DataIOut_341, DataIOut_340, DataIOut_339, 
      DataIOut_338, DataIOut_337, DataIOut_336, DataIOut_335, DataIOut_334, 
      DataIOut_333, DataIOut_332, DataIOut_331, DataIOut_330, DataIOut_329, 
      DataIOut_328, DataIOut_327, DataIOut_326, DataIOut_325, DataIOut_324, 
      DataIOut_323, DataIOut_322, DataIOut_321, DataIOut_320, DataIOut_319, 
      DataIOut_318, DataIOut_317, DataIOut_316, DataIOut_315, DataIOut_314, 
      DataIOut_313, DataIOut_312, DataIOut_311, DataIOut_310, DataIOut_309, 
      DataIOut_308, DataIOut_307, DataIOut_306, DataIOut_305, DataIOut_304, 
      DataIOut_303, DataIOut_302, DataIOut_301, DataIOut_300, DataIOut_299, 
      DataIOut_298, DataIOut_297, DataIOut_296, DataIOut_295, DataIOut_294, 
      DataIOut_293, DataIOut_292, DataIOut_291, DataIOut_290, DataIOut_289, 
      DataIOut_288, DataIOut_287, DataIOut_286, DataIOut_285, DataIOut_284, 
      DataIOut_283, DataIOut_282, DataIOut_281, DataIOut_280, DataIOut_279, 
      DataIOut_278, DataIOut_277, DataIOut_276, DataIOut_275, DataIOut_274, 
      DataIOut_273, DataIOut_272, DataIOut_271, DataIOut_270, DataIOut_269, 
      DataIOut_268, DataIOut_267, DataIOut_266, DataIOut_265, DataIOut_264, 
      DataIOut_263, DataIOut_262, DataIOut_261, DataIOut_260, DataIOut_259, 
      DataIOut_258, DataIOut_257, DataIOut_256, DataIOut_255, DataIOut_254, 
      DataIOut_253, DataIOut_252, DataIOut_251, DataIOut_250, DataIOut_249, 
      DataIOut_248, DataIOut_247, DataIOut_246, DataIOut_245, DataIOut_244, 
      DataIOut_243, DataIOut_242, DataIOut_241, DataIOut_240, DataIOut_239, 
      DataIOut_238, DataIOut_237, DataIOut_236, DataIOut_235, DataIOut_234, 
      DataIOut_233, DataIOut_232, DataIOut_231, DataIOut_230, DataIOut_229, 
      DataIOut_228, DataIOut_227, DataIOut_226, DataIOut_225, DataIOut_224, 
      DataIOut_223, DataIOut_222, DataIOut_221, DataIOut_220, DataIOut_219, 
      DataIOut_218, DataIOut_217, DataIOut_216, DataIOut_215, DataIOut_214, 
      DataIOut_213, DataIOut_212, DataIOut_211, DataIOut_210, DataIOut_209, 
      DataIOut_208, DataIOut_207, DataIOut_206, DataIOut_205, DataIOut_204, 
      DataIOut_203, DataIOut_202, DataIOut_201, DataIOut_200, DataIOut_199, 
      DataIOut_198, DataIOut_197, DataIOut_196, DataIOut_195, DataIOut_194, 
      DataIOut_193, DataIOut_192, DataIOut_191, DataIOut_190, DataIOut_189, 
      DataIOut_188, DataIOut_187, DataIOut_186, DataIOut_185, DataIOut_184, 
      DataIOut_183, DataIOut_182, DataIOut_181, DataIOut_180, DataIOut_179, 
      DataIOut_178, DataIOut_177, DataIOut_176, DataIOut_175, DataIOut_174, 
      DataIOut_173, DataIOut_172, DataIOut_171, DataIOut_170, DataIOut_169, 
      DataIOut_168, DataIOut_167, DataIOut_166, DataIOut_165, DataIOut_164, 
      DataIOut_163, DataIOut_162, DataIOut_161, DataIOut_160, DataIOut_159, 
      DataIOut_158, DataIOut_157, DataIOut_156, DataIOut_155, DataIOut_154, 
      DataIOut_153, DataIOut_152, DataIOut_151, DataIOut_150, DataIOut_149, 
      DataIOut_148, DataIOut_147, DataIOut_146, DataIOut_145, DataIOut_144, 
      DataIOut_143, DataIOut_142, DataIOut_141, DataIOut_140, DataIOut_139, 
      DataIOut_138, DataIOut_137, DataIOut_136, DataIOut_135, DataIOut_134, 
      DataIOut_133, DataIOut_132, DataIOut_131, DataIOut_130, DataIOut_129, 
      DataIOut_128, DataIOut_127, DataIOut_126, DataIOut_125, DataIOut_124, 
      DataIOut_123, DataIOut_122, DataIOut_121, DataIOut_120, DataIOut_119, 
      DataIOut_118, DataIOut_117, DataIOut_116, DataIOut_115, DataIOut_114, 
      DataIOut_113, DataIOut_112, DataIOut_111, DataIOut_110, DataIOut_109, 
      DataIOut_108, DataIOut_107, DataIOut_106, DataIOut_105, DataIOut_104, 
      DataIOut_103, DataIOut_102, DataIOut_101, DataIOut_100, DataIOut_99, 
      DataIOut_98, DataIOut_97, DataIOut_96, DataIOut_95, DataIOut_94, 
      DataIOut_93, DataIOut_92, DataIOut_91, DataIOut_90, DataIOut_89, 
      DataIOut_88, DataIOut_87, DataIOut_86, DataIOut_85, DataIOut_84, 
      DataIOut_83, DataIOut_82, DataIOut_81, DataIOut_80, DataIOut_79, 
      DataIOut_78, DataIOut_77, DataIOut_76, DataIOut_75, DataIOut_74, 
      DataIOut_73, DataIOut_72, DataIOut_71, DataIOut_70, DataIOut_69, 
      DataIOut_68, DataIOut_67, DataIOut_66, DataIOut_65, DataIOut_64, 
      DataIOut_63, DataIOut_62, DataIOut_61, DataIOut_60, DataIOut_59, 
      DataIOut_58, DataIOut_57, DataIOut_56, DataIOut_55, DataIOut_54, 
      DataIOut_53, DataIOut_52, DataIOut_51, DataIOut_50, DataIOut_49, 
      DataIOut_48, DataIOut_47, DataIOut_46, DataIOut_45, DataIOut_44, 
      DataIOut_43, DataIOut_42, DataIOut_41, DataIOut_40, DataIOut_39, 
      DataIOut_38, DataIOut_37, DataIOut_36, DataIOut_35, DataIOut_34, 
      DataIOut_33, DataIOut_32, DataIOut_31, DataIOut_30, DataIOut_29, 
      DataIOut_28, DataIOut_27, DataIOut_26, DataIOut_25, DataIOut_24, 
      DataIOut_23, DataIOut_22, DataIOut_21, DataIOut_20, DataIOut_19, 
      DataIOut_18, DataIOut_17, DataIOut_16, DataIOut_15, DataIOut_14, 
      DataIOut_13, DataIOut_12, DataIOut_11, DataIOut_10, DataIOut_9, 
      DataIOut_8, DataIOut_7, DataIOut_6, DataIOut_5, DataIOut_4, DataIOut_3, 
      DataIOut_2, DataIOut_1, DataIOut_0, NoOfLayers_1, NoOfLayers_0, 
      LayerInfoOut_15, LayerInfoOut_14, LayerInfoOut_12, LayerInfoOut_11, 
      LayerInfoOut_10, LayerInfoOut_9, LayerInfoOut_8, LayerInfoOut_7, 
      LayerInfoOut_6, LayerInfoOut_5, LayerInfoOut_4, LayerInfoOut_3, 
      LayerInfoOut_2, LayerInfoOut_1, LayerInfoOut_0, ImgWidthOut_15, 
      ImgWidthOut_14, ImgWidthOut_13, ImgWidthOut_12, ImgWidthOut_11, 
      ImgWidthOut_10, ImgWidthOut_9, ImgWidthOut_8, ImgWidthOut_7, 
      ImgWidthOut_6, ImgWidthOut_5, ImgWidthOut_4, ImgWidthOut_3, 
      ImgWidthOut_2, ImgWidthOut_1, ImgWidthOut_0, WidthSquareOut_9, 
      WidthSquareOut_8, WidthSquareOut_7, WidthSquareOut_6, WidthSquareOut_5, 
      WidthSquareOut_4, WidthSquareOut_3, WidthSquareOut_2, WidthSquareOut_1, 
      WidthSquareOut_0, Bias0_15, Bias0_14, Bias0_13, Bias0_12, Bias0_11, 
      Bias0_10, Bias0_9, Bias0_8, Bias0_7, Bias0_6, Bias0_5, Bias0_4, 
      Bias0_3, Bias0_2, Bias0_1, Bias0_0, Bias1_15, Bias1_14, Bias1_13, 
      Bias1_12, Bias1_11, Bias1_10, Bias1_9, Bias1_8, Bias1_7, Bias1_6, 
      Bias1_5, Bias1_4, Bias1_3, Bias1_2, Bias1_1, Bias1_0, Bias2_15, 
      Bias2_14, Bias2_13, Bias2_12, Bias2_11, Bias2_10, Bias2_9, Bias2_8, 
      Bias2_7, Bias2_6, Bias2_5, Bias2_4, Bias2_3, Bias2_2, Bias2_1, Bias2_0, 
      Bias3_15, Bias3_14, Bias3_13, Bias3_12, Bias3_11, Bias3_10, Bias3_9, 
      Bias3_8, Bias3_7, Bias3_6, Bias3_5, Bias3_4, Bias3_3, Bias3_2, Bias3_1, 
      Bias3_0, Bias4_15, Bias4_14, Bias4_13, Bias4_12, Bias4_11, Bias4_10, 
      Bias4_9, Bias4_8, Bias4_7, Bias4_6, Bias4_5, Bias4_4, Bias4_3, Bias4_2, 
      Bias4_1, Bias4_0, Bias5_15, Bias5_14, Bias5_13, Bias5_12, Bias5_11, 
      Bias5_10, Bias5_9, Bias5_8, Bias5_7, Bias5_6, Bias5_5, Bias5_4, 
      Bias5_3, Bias5_2, Bias5_1, Bias5_0, Bias6_15, Bias6_14, Bias6_13, 
      Bias6_12, Bias6_11, Bias6_10, Bias6_9, Bias6_8, Bias6_7, Bias6_6, 
      Bias6_5, Bias6_4, Bias6_3, Bias6_2, Bias6_1, Bias6_0, Bias7_15, 
      Bias7_14, Bias7_13, Bias7_12, Bias7_11, Bias7_10, Bias7_9, Bias7_8, 
      Bias7_7, Bias7_6, Bias7_5, Bias7_4, Bias7_3, Bias7_2, Bias7_1, Bias7_0, 
      IndicatorF_0, Filter2_399, Filter2_398, Filter2_397, Filter2_396, 
      Filter2_395, Filter2_394, Filter2_393, Filter2_392, Filter2_391, 
      Filter2_390, Filter2_389, Filter2_388, Filter2_387, Filter2_386, 
      Filter2_385, Filter2_384, Filter2_383, Filter2_382, Filter2_381, 
      Filter2_380, Filter2_379, Filter2_378, Filter2_377, Filter2_376, 
      Filter2_375, Filter2_374, Filter2_373, Filter2_372, Filter2_371, 
      Filter2_370, Filter2_369, Filter2_368, Filter2_367, Filter2_366, 
      Filter2_365, Filter2_364, Filter2_363, Filter2_362, Filter2_361, 
      Filter2_360, Filter2_359, Filter2_358, Filter2_357, Filter2_356, 
      Filter2_355, Filter2_354, Filter2_353, Filter2_352, Filter2_351, 
      Filter2_350, Filter2_349, Filter2_348, Filter2_347, Filter2_346, 
      Filter2_345, Filter2_344, Filter2_343, Filter2_342, Filter2_341, 
      Filter2_340, Filter2_339, Filter2_338, Filter2_337, Filter2_336, 
      Filter2_335, Filter2_334, Filter2_333, Filter2_332, Filter2_331, 
      Filter2_330, Filter2_329, Filter2_328, Filter2_327, Filter2_326, 
      Filter2_325, Filter2_324, Filter2_323, Filter2_322, Filter2_321, 
      Filter2_320, Filter2_319, Filter2_318, Filter2_317, Filter2_316, 
      Filter2_315, Filter2_314, Filter2_313, Filter2_312, Filter2_311, 
      Filter2_310, Filter2_309, Filter2_308, Filter2_307, Filter2_306, 
      Filter2_305, Filter2_304, Filter2_303, Filter2_302, Filter2_301, 
      Filter2_300, Filter2_299, Filter2_298, Filter2_297, Filter2_296, 
      Filter2_295, Filter2_294, Filter2_293, Filter2_292, Filter2_291, 
      Filter2_290, Filter2_289, Filter2_288, Filter2_287, Filter2_286, 
      Filter2_285, Filter2_284, Filter2_283, Filter2_282, Filter2_281, 
      Filter2_280, Filter2_279, Filter2_278, Filter2_277, Filter2_276, 
      Filter2_275, Filter2_274, Filter2_273, Filter2_272, Filter2_271, 
      Filter2_270, Filter2_269, Filter2_268, Filter2_267, Filter2_266, 
      Filter2_265, Filter2_264, Filter2_263, Filter2_262, Filter2_261, 
      Filter2_260, Filter2_259, Filter2_258, Filter2_257, Filter2_256, 
      Filter2_255, Filter2_254, Filter2_253, Filter2_252, Filter2_251, 
      Filter2_250, Filter2_249, Filter2_248, Filter2_247, Filter2_246, 
      Filter2_245, Filter2_244, Filter2_243, Filter2_242, Filter2_241, 
      Filter2_240, Filter2_239, Filter2_238, Filter2_237, Filter2_236, 
      Filter2_235, Filter2_234, Filter2_233, Filter2_232, Filter2_231, 
      Filter2_230, Filter2_229, Filter2_228, Filter2_227, Filter2_226, 
      Filter2_225, Filter2_224, Filter2_223, Filter2_222, Filter2_221, 
      Filter2_220, Filter2_219, Filter2_218, Filter2_217, Filter2_216, 
      Filter2_215, Filter2_214, Filter2_213, Filter2_212, Filter2_211, 
      Filter2_210, Filter2_209, Filter2_208, Filter2_207, Filter2_206, 
      Filter2_205, Filter2_204, Filter2_203, Filter2_202, Filter2_201, 
      Filter2_200, Filter2_199, Filter2_198, Filter2_197, Filter2_196, 
      Filter2_195, Filter2_194, Filter2_193, Filter2_192, Filter2_191, 
      Filter2_190, Filter2_189, Filter2_188, Filter2_187, Filter2_186, 
      Filter2_185, Filter2_184, Filter2_183, Filter2_182, Filter2_181, 
      Filter2_180, Filter2_179, Filter2_178, Filter2_177, Filter2_176, 
      Filter2_175, Filter2_174, Filter2_173, Filter2_172, Filter2_171, 
      Filter2_170, Filter2_169, Filter2_168, Filter2_167, Filter2_166, 
      Filter2_165, Filter2_164, Filter2_163, Filter2_162, Filter2_161, 
      Filter2_160, Filter2_159, Filter2_158, Filter2_157, Filter2_156, 
      Filter2_155, Filter2_154, Filter2_153, Filter2_152, Filter2_151, 
      Filter2_150, Filter2_149, Filter2_148, Filter2_147, Filter2_146, 
      Filter2_145, Filter2_144, Filter2_143, Filter2_142, Filter2_141, 
      Filter2_140, Filter2_139, Filter2_138, Filter2_137, Filter2_136, 
      Filter2_135, Filter2_134, Filter2_133, Filter2_132, Filter2_131, 
      Filter2_130, Filter2_129, Filter2_128, Filter2_127, Filter2_126, 
      Filter2_125, Filter2_124, Filter2_123, Filter2_122, Filter2_121, 
      Filter2_120, Filter2_119, Filter2_118, Filter2_117, Filter2_116, 
      Filter2_115, Filter2_114, Filter2_113, Filter2_112, Filter2_111, 
      Filter2_110, Filter2_109, Filter2_108, Filter2_107, Filter2_106, 
      Filter2_105, Filter2_104, Filter2_103, Filter2_102, Filter2_101, 
      Filter2_100, Filter2_99, Filter2_98, Filter2_97, Filter2_96, 
      Filter2_95, Filter2_94, Filter2_93, Filter2_92, Filter2_91, Filter2_90, 
      Filter2_89, Filter2_88, Filter2_87, Filter2_86, Filter2_85, Filter2_84, 
      Filter2_83, Filter2_82, Filter2_81, Filter2_80, Filter2_79, Filter2_78, 
      Filter2_77, Filter2_76, Filter2_75, Filter2_74, Filter2_73, Filter2_72, 
      Filter2_71, Filter2_70, Filter2_69, Filter2_68, Filter2_67, Filter2_66, 
      Filter2_65, Filter2_64, Filter2_63, Filter2_62, Filter2_61, Filter2_60, 
      Filter2_59, Filter2_58, Filter2_57, Filter2_56, Filter2_55, Filter2_54, 
      Filter2_53, Filter2_52, Filter2_51, Filter2_50, Filter2_49, Filter2_48, 
      Filter2_47, Filter2_46, Filter2_45, Filter2_44, Filter2_43, Filter2_42, 
      Filter2_41, Filter2_40, Filter2_39, Filter2_38, Filter2_37, Filter2_36, 
      Filter2_35, Filter2_34, Filter2_33, Filter2_32, Filter2_31, Filter2_30, 
      Filter2_29, Filter2_28, Filter2_27, Filter2_26, Filter2_25, Filter2_24, 
      Filter2_23, Filter2_22, Filter2_21, Filter2_20, Filter2_19, Filter2_18, 
      Filter2_17, Filter2_16, Filter2_15, Filter2_14, Filter2_13, Filter2_12, 
      Filter2_11, Filter2_10, Filter2_9, Filter2_8, Filter2_7, Filter2_6, 
      Filter2_5, Filter2_4, Filter2_3, Filter2_2, Filter2_1, Filter2_0, 
      Filter1_399, Filter1_398, Filter1_397, Filter1_396, Filter1_395, 
      Filter1_394, Filter1_393, Filter1_392, Filter1_391, Filter1_390, 
      Filter1_389, Filter1_388, Filter1_387, Filter1_386, Filter1_385, 
      Filter1_384, Filter1_383, Filter1_382, Filter1_381, Filter1_380, 
      Filter1_379, Filter1_378, Filter1_377, Filter1_376, Filter1_375, 
      Filter1_374, Filter1_373, Filter1_372, Filter1_371, Filter1_370, 
      Filter1_369, Filter1_368, Filter1_367, Filter1_366, Filter1_365, 
      Filter1_364, Filter1_363, Filter1_362, Filter1_361, Filter1_360, 
      Filter1_359, Filter1_358, Filter1_357, Filter1_356, Filter1_355, 
      Filter1_354, Filter1_353, Filter1_352, Filter1_351, Filter1_350, 
      Filter1_349, Filter1_348, Filter1_347, Filter1_346, Filter1_345, 
      Filter1_344, Filter1_343, Filter1_342, Filter1_341, Filter1_340, 
      Filter1_339, Filter1_338, Filter1_337, Filter1_336, Filter1_335, 
      Filter1_334, Filter1_333, Filter1_332, Filter1_331, Filter1_330, 
      Filter1_329, Filter1_328, Filter1_327, Filter1_326, Filter1_325, 
      Filter1_324, Filter1_323, Filter1_322, Filter1_321, Filter1_320, 
      Filter1_319, Filter1_318, Filter1_317, Filter1_316, Filter1_315, 
      Filter1_314, Filter1_313, Filter1_312, Filter1_311, Filter1_310, 
      Filter1_309, Filter1_308, Filter1_307, Filter1_306, Filter1_305, 
      Filter1_304, Filter1_303, Filter1_302, Filter1_301, Filter1_300, 
      Filter1_299, Filter1_298, Filter1_297, Filter1_296, Filter1_295, 
      Filter1_294, Filter1_293, Filter1_292, Filter1_291, Filter1_290, 
      Filter1_289, Filter1_288, Filter1_287, Filter1_286, Filter1_285, 
      Filter1_284, Filter1_283, Filter1_282, Filter1_281, Filter1_280, 
      Filter1_279, Filter1_278, Filter1_277, Filter1_276, Filter1_275, 
      Filter1_274, Filter1_273, Filter1_272, Filter1_271, Filter1_270, 
      Filter1_269, Filter1_268, Filter1_267, Filter1_266, Filter1_265, 
      Filter1_264, Filter1_263, Filter1_262, Filter1_261, Filter1_260, 
      Filter1_259, Filter1_258, Filter1_257, Filter1_256, Filter1_255, 
      Filter1_254, Filter1_253, Filter1_252, Filter1_251, Filter1_250, 
      Filter1_249, Filter1_248, Filter1_247, Filter1_246, Filter1_245, 
      Filter1_244, Filter1_243, Filter1_242, Filter1_241, Filter1_240, 
      Filter1_239, Filter1_238, Filter1_237, Filter1_236, Filter1_235, 
      Filter1_234, Filter1_233, Filter1_232, Filter1_231, Filter1_230, 
      Filter1_229, Filter1_228, Filter1_227, Filter1_226, Filter1_225, 
      Filter1_224, Filter1_223, Filter1_222, Filter1_221, Filter1_220, 
      Filter1_219, Filter1_218, Filter1_217, Filter1_216, Filter1_215, 
      Filter1_214, Filter1_213, Filter1_212, Filter1_211, Filter1_210, 
      Filter1_209, Filter1_208, Filter1_207, Filter1_206, Filter1_205, 
      Filter1_204, Filter1_203, Filter1_202, Filter1_201, Filter1_200, 
      Filter1_199, Filter1_198, Filter1_197, Filter1_196, Filter1_195, 
      Filter1_194, Filter1_193, Filter1_192, Filter1_191, Filter1_190, 
      Filter1_189, Filter1_188, Filter1_187, Filter1_186, Filter1_185, 
      Filter1_184, Filter1_183, Filter1_182, Filter1_181, Filter1_180, 
      Filter1_179, Filter1_178, Filter1_177, Filter1_176, Filter1_175, 
      Filter1_174, Filter1_173, Filter1_172, Filter1_171, Filter1_170, 
      Filter1_169, Filter1_168, Filter1_167, Filter1_166, Filter1_165, 
      Filter1_164, Filter1_163, Filter1_162, Filter1_161, Filter1_160, 
      Filter1_159, Filter1_158, Filter1_157, Filter1_156, Filter1_155, 
      Filter1_154, Filter1_153, Filter1_152, Filter1_151, Filter1_150, 
      Filter1_149, Filter1_148, Filter1_147, Filter1_146, Filter1_145, 
      Filter1_144, Filter1_143, Filter1_142, Filter1_141, Filter1_140, 
      Filter1_139, Filter1_138, Filter1_137, Filter1_136, Filter1_135, 
      Filter1_134, Filter1_133, Filter1_132, Filter1_131, Filter1_130, 
      Filter1_129, Filter1_128, Filter1_127, Filter1_126, Filter1_125, 
      Filter1_124, Filter1_123, Filter1_122, Filter1_121, Filter1_120, 
      Filter1_119, Filter1_118, Filter1_117, Filter1_116, Filter1_115, 
      Filter1_114, Filter1_113, Filter1_112, Filter1_111, Filter1_110, 
      Filter1_109, Filter1_108, Filter1_107, Filter1_106, Filter1_105, 
      Filter1_104, Filter1_103, Filter1_102, Filter1_101, Filter1_100, 
      Filter1_99, Filter1_98, Filter1_97, Filter1_96, Filter1_95, Filter1_94, 
      Filter1_93, Filter1_92, Filter1_91, Filter1_90, Filter1_89, Filter1_88, 
      Filter1_87, Filter1_86, Filter1_85, Filter1_84, Filter1_83, Filter1_82, 
      Filter1_81, Filter1_80, Filter1_79, Filter1_78, Filter1_77, Filter1_76, 
      Filter1_75, Filter1_74, Filter1_73, Filter1_72, Filter1_71, Filter1_70, 
      Filter1_69, Filter1_68, Filter1_67, Filter1_66, Filter1_65, Filter1_64, 
      Filter1_63, Filter1_62, Filter1_61, Filter1_60, Filter1_59, Filter1_58, 
      Filter1_57, Filter1_56, Filter1_55, Filter1_54, Filter1_53, Filter1_52, 
      Filter1_51, Filter1_50, Filter1_49, Filter1_48, Filter1_47, Filter1_46, 
      Filter1_45, Filter1_44, Filter1_43, Filter1_42, Filter1_41, Filter1_40, 
      Filter1_39, Filter1_38, Filter1_37, Filter1_36, Filter1_35, Filter1_34, 
      Filter1_33, Filter1_32, Filter1_31, Filter1_30, Filter1_29, Filter1_28, 
      Filter1_27, Filter1_26, Filter1_25, Filter1_24, Filter1_23, Filter1_22, 
      Filter1_21, Filter1_20, Filter1_19, Filter1_18, Filter1_17, Filter1_16, 
      Filter1_15, Filter1_14, Filter1_13, Filter1_12, Filter1_11, Filter1_10, 
      Filter1_9, Filter1_8, Filter1_7, Filter1_6, Filter1_5, Filter1_4, 
      Filter1_3, Filter1_2, Filter1_1, Filter1_0, IndicatorI_0, 
      ImgCounterOuput_2, ImgCounterOuput_1, ImgCounterOuput_0, OutputImg0_79, 
      OutputImg0_78, OutputImg0_77, OutputImg0_76, OutputImg0_75, 
      OutputImg0_74, OutputImg0_73, OutputImg0_72, OutputImg0_71, 
      OutputImg0_70, OutputImg0_69, OutputImg0_68, OutputImg0_67, 
      OutputImg0_66, OutputImg0_65, OutputImg0_64, OutputImg0_63, 
      OutputImg0_62, OutputImg0_61, OutputImg0_60, OutputImg0_59, 
      OutputImg0_58, OutputImg0_57, OutputImg0_56, OutputImg0_55, 
      OutputImg0_54, OutputImg0_53, OutputImg0_52, OutputImg0_51, 
      OutputImg0_50, OutputImg0_49, OutputImg0_48, OutputImg0_47, 
      OutputImg0_46, OutputImg0_45, OutputImg0_44, OutputImg0_43, 
      OutputImg0_42, OutputImg0_41, OutputImg0_40, OutputImg0_39, 
      OutputImg0_38, OutputImg0_37, OutputImg0_36, OutputImg0_35, 
      OutputImg0_34, OutputImg0_33, OutputImg0_32, OutputImg0_31, 
      OutputImg0_30, OutputImg0_29, OutputImg0_28, OutputImg0_27, 
      OutputImg0_26, OutputImg0_25, OutputImg0_24, OutputImg0_23, 
      OutputImg0_22, OutputImg0_21, OutputImg0_20, OutputImg0_19, 
      OutputImg0_18, OutputImg0_17, OutputImg0_16, OutputImg0_15, 
      OutputImg0_14, OutputImg0_13, OutputImg0_12, OutputImg0_11, 
      OutputImg0_10, OutputImg0_9, OutputImg0_8, OutputImg0_7, OutputImg0_6, 
      OutputImg0_5, OutputImg0_4, OutputImg0_3, OutputImg0_2, OutputImg0_1, 
      OutputImg0_0, OutputImg1_79, OutputImg1_78, OutputImg1_77, 
      OutputImg1_76, OutputImg1_75, OutputImg1_74, OutputImg1_73, 
      OutputImg1_72, OutputImg1_71, OutputImg1_70, OutputImg1_69, 
      OutputImg1_68, OutputImg1_67, OutputImg1_66, OutputImg1_65, 
      OutputImg1_64, OutputImg1_63, OutputImg1_62, OutputImg1_61, 
      OutputImg1_60, OutputImg1_59, OutputImg1_58, OutputImg1_57, 
      OutputImg1_56, OutputImg1_55, OutputImg1_54, OutputImg1_53, 
      OutputImg1_52, OutputImg1_51, OutputImg1_50, OutputImg1_49, 
      OutputImg1_48, OutputImg1_47, OutputImg1_46, OutputImg1_45, 
      OutputImg1_44, OutputImg1_43, OutputImg1_42, OutputImg1_41, 
      OutputImg1_40, OutputImg1_39, OutputImg1_38, OutputImg1_37, 
      OutputImg1_36, OutputImg1_35, OutputImg1_34, OutputImg1_33, 
      OutputImg1_32, OutputImg1_31, OutputImg1_30, OutputImg1_29, 
      OutputImg1_28, OutputImg1_27, OutputImg1_26, OutputImg1_25, 
      OutputImg1_24, OutputImg1_23, OutputImg1_22, OutputImg1_21, 
      OutputImg1_20, OutputImg1_19, OutputImg1_18, OutputImg1_17, 
      OutputImg1_16, OutputImg1_15, OutputImg1_14, OutputImg1_13, 
      OutputImg1_12, OutputImg1_11, OutputImg1_10, OutputImg1_9, 
      OutputImg1_8, OutputImg1_7, OutputImg1_6, OutputImg1_5, OutputImg1_4, 
      OutputImg1_3, OutputImg1_2, OutputImg1_1, OutputImg1_0, OutputImg2_79, 
      OutputImg2_78, OutputImg2_77, OutputImg2_76, OutputImg2_75, 
      OutputImg2_74, OutputImg2_73, OutputImg2_72, OutputImg2_71, 
      OutputImg2_70, OutputImg2_69, OutputImg2_68, OutputImg2_67, 
      OutputImg2_66, OutputImg2_65, OutputImg2_64, OutputImg2_63, 
      OutputImg2_62, OutputImg2_61, OutputImg2_60, OutputImg2_59, 
      OutputImg2_58, OutputImg2_57, OutputImg2_56, OutputImg2_55, 
      OutputImg2_54, OutputImg2_53, OutputImg2_52, OutputImg2_51, 
      OutputImg2_50, OutputImg2_49, OutputImg2_48, OutputImg2_47, 
      OutputImg2_46, OutputImg2_45, OutputImg2_44, OutputImg2_43, 
      OutputImg2_42, OutputImg2_41, OutputImg2_40, OutputImg2_39, 
      OutputImg2_38, OutputImg2_37, OutputImg2_36, OutputImg2_35, 
      OutputImg2_34, OutputImg2_33, OutputImg2_32, OutputImg2_31, 
      OutputImg2_30, OutputImg2_29, OutputImg2_28, OutputImg2_27, 
      OutputImg2_26, OutputImg2_25, OutputImg2_24, OutputImg2_23, 
      OutputImg2_22, OutputImg2_21, OutputImg2_20, OutputImg2_19, 
      OutputImg2_18, OutputImg2_17, OutputImg2_16, OutputImg2_15, 
      OutputImg2_14, OutputImg2_13, OutputImg2_12, OutputImg2_11, 
      OutputImg2_10, OutputImg2_9, OutputImg2_8, OutputImg2_7, OutputImg2_6, 
      OutputImg2_5, OutputImg2_4, OutputImg2_3, OutputImg2_2, OutputImg2_1, 
      OutputImg2_0, OutputImg3_79, OutputImg3_78, OutputImg3_77, 
      OutputImg3_76, OutputImg3_75, OutputImg3_74, OutputImg3_73, 
      OutputImg3_72, OutputImg3_71, OutputImg3_70, OutputImg3_69, 
      OutputImg3_68, OutputImg3_67, OutputImg3_66, OutputImg3_65, 
      OutputImg3_64, OutputImg3_63, OutputImg3_62, OutputImg3_61, 
      OutputImg3_60, OutputImg3_59, OutputImg3_58, OutputImg3_57, 
      OutputImg3_56, OutputImg3_55, OutputImg3_54, OutputImg3_53, 
      OutputImg3_52, OutputImg3_51, OutputImg3_50, OutputImg3_49, 
      OutputImg3_48, OutputImg3_47, OutputImg3_46, OutputImg3_45, 
      OutputImg3_44, OutputImg3_43, OutputImg3_42, OutputImg3_41, 
      OutputImg3_40, OutputImg3_39, OutputImg3_38, OutputImg3_37, 
      OutputImg3_36, OutputImg3_35, OutputImg3_34, OutputImg3_33, 
      OutputImg3_32, OutputImg3_31, OutputImg3_30, OutputImg3_29, 
      OutputImg3_28, OutputImg3_27, OutputImg3_26, OutputImg3_25, 
      OutputImg3_24, OutputImg3_23, OutputImg3_22, OutputImg3_21, 
      OutputImg3_20, OutputImg3_19, OutputImg3_18, OutputImg3_17, 
      OutputImg3_16, OutputImg3_15, OutputImg3_14, OutputImg3_13, 
      OutputImg3_12, OutputImg3_11, OutputImg3_10, OutputImg3_9, 
      OutputImg3_8, OutputImg3_7, OutputImg3_6, OutputImg3_5, OutputImg3_4, 
      OutputImg3_3, OutputImg3_2, OutputImg3_1, OutputImg3_0, OutputImg4_79, 
      OutputImg4_78, OutputImg4_77, OutputImg4_76, OutputImg4_75, 
      OutputImg4_74, OutputImg4_73, OutputImg4_72, OutputImg4_71, 
      OutputImg4_70, OutputImg4_69, OutputImg4_68, OutputImg4_67, 
      OutputImg4_66, OutputImg4_65, OutputImg4_64, OutputImg4_63, 
      OutputImg4_62, OutputImg4_61, OutputImg4_60, OutputImg4_59, 
      OutputImg4_58, OutputImg4_57, OutputImg4_56, OutputImg4_55, 
      OutputImg4_54, OutputImg4_53, OutputImg4_52, OutputImg4_51, 
      OutputImg4_50, OutputImg4_49, OutputImg4_48, OutputImg4_47, 
      OutputImg4_46, OutputImg4_45, OutputImg4_44, OutputImg4_43, 
      OutputImg4_42, OutputImg4_41, OutputImg4_40, OutputImg4_39, 
      OutputImg4_38, OutputImg4_37, OutputImg4_36, OutputImg4_35, 
      OutputImg4_34, OutputImg4_33, OutputImg4_32, OutputImg4_31, 
      OutputImg4_30, OutputImg4_29, OutputImg4_28, OutputImg4_27, 
      OutputImg4_26, OutputImg4_25, OutputImg4_24, OutputImg4_23, 
      OutputImg4_22, OutputImg4_21, OutputImg4_20, OutputImg4_19, 
      OutputImg4_18, OutputImg4_17, OutputImg4_16, OutputImg4_15, 
      OutputImg4_14, OutputImg4_13, OutputImg4_12, OutputImg4_11, 
      OutputImg4_10, OutputImg4_9, OutputImg4_8, OutputImg4_7, OutputImg4_6, 
      OutputImg4_5, OutputImg4_4, OutputImg4_3, OutputImg4_2, OutputImg4_1, 
      OutputImg4_0, ConvOuput_15, ConvOuput_14, ConvOuput_13, ConvOuput_12, 
      ConvOuput_11, ConvOuput_10, ConvOuput_9, ConvOuput_8, ConvOuput_7, 
      ConvOuput_6, ConvOuput_5, ConvOuput_4, ConvOuput_3, ConvOuput_2, 
      ConvOuput_1, ConvOuput_0, ShiftLeftCounterOutput_4, 
      ShiftLeftCounterOutput_3, ShiftLeftCounterOutput_2, 
      ShiftLeftCounterOutput_1, ShiftLeftCounterOutput_0, 
      RealOutputCounter_12, RealOutputCounter_11, RealOutputCounter_10, 
      RealOutputCounter_9, RealOutputCounter_8, RealOutputCounter_7, 
      RealOutputCounter_6, RealOutputCounter_5, RealOutputCounter_4, 
      RealOutputCounter_3, RealOutputCounter_2, RealOutputCounter_1, 
      RealOutputCounter_0, OutputCounterLoad_12, OutputCounterLoad_11, 
      OutputCounterLoad_10, OutputCounterLoad_9, OutputCounterLoad_8, 
      OutputCounterLoad_7, OutputCounterLoad_6, OutputCounterLoad_5, 
      OutputCounterLoad_4, OutputCounterLoad_3, OutputCounterLoad_2, 
      OutputCounterLoad_1, OutputCounterLoad_0, Q, NumOfFilters_3, 
      NumOfFilters_2, NumOfFilters_1, NumOfFilters_0, NumOfHeight_4, 
      NumOfHeight_3, NumOfHeight_2, NumOfHeight_1, NumOfHeight_0, X, Y, K, L, 
      D, CNDepthoutput_3, CNDepthoutput_2, CNDepthoutput_1, CNDepthoutput_0, 
      SwitchMEM_0, SwitchBar_0, CLK, DontRstIndicator, lastFilter, 
      lastDepthOut, SwitchClk, TriStateCounterEN, FilterAddressEN, 
      ImgAddRegEN, ShiftCounterRst, AddressChangerEN, TriChnagerToaddEN, 
      ImgAddRST, ramSelector, zero_11, PWR, next_state_5, next_state_14, 
      next_state_dup_134, NOT_L, next_state_13, next_state_12, next_state_11, 
      nx18, nx20, next_state_10, next_state_9, next_state_dup_124, 
      next_state_8, next_state_7, next_state_dup_96, nx48, next_state_6, 
      nx9711, nx66, next_state_3, next_state_2, next_state_dup_26, NOT_nx0, 
      next_state_1, next_state_dup_147, nx100, nx112, nx130, nx142, nx154, 
      SaveAckLatch, nx180, nx186, nx9063, nx210, nx224, nx240, nx256, nx270, 
      nx300, next_state_4, next_state_dup_24, nx322, nx350, nx382, nx416, 
      nx418, nx456, nx466, nx478, nx480, nx482, nx494, nx9718, nx9728, 
      nx9738, nx9748, nx9760, nx9765, nx9768, nx9780, nx9792, nx9796, nx9814, 
      nx9822, nx9824, nx9826, nx9833, nx9835, nx9849, nx9854, nx9856, nx9858, 
      nx9866, nx9870, nx9875, nx9879, nx9881, nx9883, nx9885, nx9887, nx9889, 
      nx9891, nx9893, nx9899, nx9901, nx9903, nx9905, nx9908, nx9911, nx9913, 
      nx9916, nx9921, nx9923, nx9925, nx9932, nx9934, nx9937, nx9939, nx9941, 
      nx9950, nx9952, nx9954, nx9956, nx9958, nx9960, nx9962, nx9964, nx9966, 
      nx9968, nx9970, nx9972, nx9974, nx9976, nx9978, nx9980, nx9982, nx9984, 
      nx9986, nx9988, nx9990, nx9992, nx9994, nx9996, nx9998, nx10000, 
      nx10002, nx10004, nx10006, nx10008, nx10010, nx10012, nx10014, nx10016, 
      nx10018, nx10020, nx10022, nx10024, nx10026, nx10028, nx10032, nx10034, 
      nx10036, nx10038, nx10040, nx10042, nx10044, nx10046, nx10048, nx10050, 
      nx10052, nx10054, nx10056, nx10058, nx10060, nx10062, nx10064, nx10066, 
      nx10068, nx10070, nx10072, nx10074, nx10076, nx10078, nx10080, nx10082, 
      nx10084, nx10086, nx10088, nx10090, nx10092, nx10094, nx10096, nx10098, 
      nx10100, nx10102, nx10104, nx10106, nx10108, nx10110, nx10112, nx10114, 
      nx10116, nx10118, nx10120, nx10122, nx10124, nx10126, nx10128, nx10130, 
      nx10132, nx10134, nx10136, nx10138, nx10140, nx10142, nx10144, nx10146, 
      nx10148, nx10150, nx10152, nx10154, nx10156, nx10158, nx10160, nx10162, 
      nx10164, nx10166, nx10168, nx10170, nx10172, nx10174, nx10176, nx10178, 
      nx10180, nx10182, nx10184, nx10186, nx10188, nx10190, nx10192, nx10194, 
      nx10196, nx10198, nx10200, nx10202, nx10204, nx10206, nx10208, nx10210, 
      nx10212, nx10214, nx10216, nx10218, nx10220, nx10222, nx10224, nx10226, 
      nx10228, nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, nx10242, 
      nx10244, nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, 
      nx10260, nx10262, nx10264, nx10266, nx10268, nx10270, nx10272, nx10274, 
      nx10276, nx10278, nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, 
      nx10292, nx10294, nx10296, nx10298, nx10300, nx10302, nx10304, nx10306, 
      nx10308, nx10310, nx10312, nx10314, nx10316, nx10318, nx10320, nx10322, 
      nx10324, nx10326, nx10328, nx10330, nx10332, nx10334, nx10336, nx10338, 
      nx10340, nx10342, nx10344, nx10346, nx10348, nx10350, nx10352, nx10354, 
      nx10356, nx10358, nx10360, nx10362, nx10364, nx10366, nx10368, nx10370, 
      nx10372, nx10374, nx10376, nx10378, nx10380, nx10382, nx10384, nx10386, 
      nx10388, nx10390, nx10392, nx10394, nx10396, nx10398, nx10400, nx10402, 
      nx10404, nx10406, nx10408, nx10410, nx10412, nx10414, nx10416, nx10418, 
      nx10420, nx10422, nx10424, nx10426, nx10428, nx10430, nx10432, nx10434, 
      nx10436, nx10438, nx10440, nx10442, nx10444, nx10446, nx10448, nx10450, 
      nx10452, nx10454, nx10456, nx10458, nx10460, nx10462, nx10464, nx10466, 
      nx10468, nx10470, nx10472, nx10474, nx10476, nx10478, nx10484, nx10486, 
      nx10488, nx10490, nx10496, nx10498, nx5, nx10500, nx10502, nx10504: 
   std_logic ;
   
   signal DANGLING : std_logic_vector (2728 downto 0 );

begin
   done <= done_EXMPLR ;
   DDF0 : nBitRegister_1 port map ( D(0)=>SwitchBar_0, CLK=>SwitchClk, RST=>
      rst, EN=>PWR, Q(0)=>SwitchMEM_0);
   TriStateAddchanger : triStateBuffer_13 port map ( D(12)=>nx9974, D(11)=>
      nx9978, D(10)=>nx9982, D(9)=>nx9986, D(8)=>nx9990, D(7)=>nx9994, D(6)
      =>nx9998, D(5)=>nx10002, D(4)=>nx10006, D(3)=>nx10010, D(2)=>nx10014, 
      D(1)=>nx10018, D(0)=>nx10022, EN=>nx9958, F(12)=>AddressChangerIN_12, 
      F(11)=>AddressChangerIN_11, F(10)=>AddressChangerIN_10, F(9)=>
      AddressChangerIN_9, F(8)=>AddressChangerIN_8, F(7)=>AddressChangerIN_7, 
      F(6)=>AddressChangerIN_6, F(5)=>AddressChangerIN_5, F(4)=>
      AddressChangerIN_4, F(3)=>AddressChangerIN_3, F(2)=>AddressChangerIN_2, 
      F(1)=>AddressChangerIN_1, F(0)=>AddressChangerIN_0);
   TriStateAddgfd : triStateBuffer_13 port map ( D(12)=>AddressChangerOut_12, 
      D(11)=>AddressChangerOut_11, D(10)=>AddressChangerOut_10, D(9)=>
      AddressChangerOut_9, D(8)=>AddressChangerOut_8, D(7)=>
      AddressChangerOut_7, D(6)=>AddressChangerOut_6, D(5)=>
      AddressChangerOut_5, D(4)=>AddressChangerOut_4, D(3)=>
      AddressChangerOut_3, D(2)=>AddressChangerOut_2, D(1)=>
      AddressChangerOut_1, D(0)=>AddressChangerOut_0, EN=>TriChnagerToaddEN, 
      F(12)=>FilterAddressIN_12, F(11)=>FilterAddressIN_11, F(10)=>
      FilterAddressIN_10, F(9)=>FilterAddressIN_9, F(8)=>FilterAddressIN_8, 
      F(7)=>FilterAddressIN_7, F(6)=>FilterAddressIN_6, F(5)=>
      FilterAddressIN_5, F(4)=>FilterAddressIN_4, F(3)=>FilterAddressIN_3, 
      F(2)=>FilterAddressIN_2, F(1)=>FilterAddressIN_1, F(0)=>
      FilterAddressIN_0);
   addChanger : nBitRegister_13 port map ( D(12)=>AddressChangerIN_12, D(11)
      =>AddressChangerIN_11, D(10)=>AddressChangerIN_10, D(9)=>
      AddressChangerIN_9, D(8)=>AddressChangerIN_8, D(7)=>AddressChangerIN_7, 
      D(6)=>AddressChangerIN_6, D(5)=>AddressChangerIN_5, D(4)=>
      AddressChangerIN_4, D(3)=>AddressChangerIN_3, D(2)=>AddressChangerIN_2, 
      D(1)=>AddressChangerIN_1, D(0)=>AddressChangerIN_0, CLK=>nx10414, RST
      =>rst, EN=>AddressChangerEN, Q(12)=>AddressChangerOut_12, Q(11)=>
      AddressChangerOut_11, Q(10)=>AddressChangerOut_10, Q(9)=>
      AddressChangerOut_9, Q(8)=>AddressChangerOut_8, Q(7)=>
      AddressChangerOut_7, Q(6)=>AddressChangerOut_6, Q(5)=>
      AddressChangerOut_5, Q(4)=>AddressChangerOut_4, Q(3)=>
      AddressChangerOut_3, Q(2)=>AddressChangerOut_2, Q(1)=>
      AddressChangerOut_1, Q(0)=>AddressChangerOut_0);
   FilterMem : RAM_25 port map ( reset=>rst, CLK=>nx10414, W=>zero_11, R=>
      ReadF, address(12)=>AddressF_12, address(11)=>AddressF_11, address(10)
      =>AddressF_10, address(9)=>AddressF_9, address(8)=>AddressF_8, 
      address(7)=>AddressF_7, address(6)=>AddressF_6, address(5)=>AddressF_5, 
      address(4)=>AddressF_4, address(3)=>AddressF_3, address(2)=>AddressF_2, 
      address(1)=>AddressF_1, address(0)=>AddressF_0, dataIn(15)=>zero_11, 
      dataIn(14)=>zero_11, dataIn(13)=>zero_11, dataIn(12)=>zero_11, 
      dataIn(11)=>zero_11, dataIn(10)=>zero_11, dataIn(9)=>zero_11, 
      dataIn(8)=>zero_11, dataIn(7)=>zero_11, dataIn(6)=>zero_11, dataIn(5)
      =>zero_11, dataIn(4)=>zero_11, dataIn(3)=>zero_11, dataIn(2)=>zero_11, 
      dataIn(1)=>zero_11, dataIn(0)=>zero_11, dataOut(399)=>DataFOut_399, 
      dataOut(398)=>DANGLING(0), dataOut(397)=>DANGLING(1), dataOut(396)=>
      DANGLING(2), dataOut(395)=>DANGLING(3), dataOut(394)=>DANGLING(4), 
      dataOut(393)=>DANGLING(5), dataOut(392)=>DANGLING(6), dataOut(391)=>
      DANGLING(7), dataOut(390)=>DANGLING(8), dataOut(389)=>DANGLING(9), 
      dataOut(388)=>DANGLING(10), dataOut(387)=>DANGLING(11), dataOut(386)=>
      DANGLING(12), dataOut(385)=>DANGLING(13), dataOut(384)=>DANGLING(14), 
      dataOut(383)=>DANGLING(15), dataOut(382)=>DANGLING(16), dataOut(381)=>
      DANGLING(17), dataOut(380)=>DANGLING(18), dataOut(379)=>DANGLING(19), 
      dataOut(378)=>DANGLING(20), dataOut(377)=>DANGLING(21), dataOut(376)=>
      DANGLING(22), dataOut(375)=>DANGLING(23), dataOut(374)=>DANGLING(24), 
      dataOut(373)=>DANGLING(25), dataOut(372)=>DANGLING(26), dataOut(371)=>
      DANGLING(27), dataOut(370)=>DANGLING(28), dataOut(369)=>DANGLING(29), 
      dataOut(368)=>DANGLING(30), dataOut(367)=>DANGLING(31), dataOut(366)=>
      DANGLING(32), dataOut(365)=>DANGLING(33), dataOut(364)=>DANGLING(34), 
      dataOut(363)=>DANGLING(35), dataOut(362)=>DANGLING(36), dataOut(361)=>
      DANGLING(37), dataOut(360)=>DANGLING(38), dataOut(359)=>DANGLING(39), 
      dataOut(358)=>DANGLING(40), dataOut(357)=>DANGLING(41), dataOut(356)=>
      DANGLING(42), dataOut(355)=>DANGLING(43), dataOut(354)=>DANGLING(44), 
      dataOut(353)=>DANGLING(45), dataOut(352)=>DANGLING(46), dataOut(351)=>
      DANGLING(47), dataOut(350)=>DANGLING(48), dataOut(349)=>DANGLING(49), 
      dataOut(348)=>DANGLING(50), dataOut(347)=>DANGLING(51), dataOut(346)=>
      DANGLING(52), dataOut(345)=>DANGLING(53), dataOut(344)=>DANGLING(54), 
      dataOut(343)=>DANGLING(55), dataOut(342)=>DANGLING(56), dataOut(341)=>
      DANGLING(57), dataOut(340)=>DANGLING(58), dataOut(339)=>DANGLING(59), 
      dataOut(338)=>DANGLING(60), dataOut(337)=>DANGLING(61), dataOut(336)=>
      DANGLING(62), dataOut(335)=>DANGLING(63), dataOut(334)=>DANGLING(64), 
      dataOut(333)=>DANGLING(65), dataOut(332)=>DANGLING(66), dataOut(331)=>
      DANGLING(67), dataOut(330)=>DANGLING(68), dataOut(329)=>DANGLING(69), 
      dataOut(328)=>DANGLING(70), dataOut(327)=>DANGLING(71), dataOut(326)=>
      DANGLING(72), dataOut(325)=>DANGLING(73), dataOut(324)=>DANGLING(74), 
      dataOut(323)=>DANGLING(75), dataOut(322)=>DANGLING(76), dataOut(321)=>
      DANGLING(77), dataOut(320)=>DANGLING(78), dataOut(319)=>DANGLING(79), 
      dataOut(318)=>DANGLING(80), dataOut(317)=>DANGLING(81), dataOut(316)=>
      DANGLING(82), dataOut(315)=>DANGLING(83), dataOut(314)=>DANGLING(84), 
      dataOut(313)=>DANGLING(85), dataOut(312)=>DANGLING(86), dataOut(311)=>
      DANGLING(87), dataOut(310)=>DANGLING(88), dataOut(309)=>DANGLING(89), 
      dataOut(308)=>DANGLING(90), dataOut(307)=>DANGLING(91), dataOut(306)=>
      DANGLING(92), dataOut(305)=>DANGLING(93), dataOut(304)=>DANGLING(94), 
      dataOut(303)=>DANGLING(95), dataOut(302)=>DANGLING(96), dataOut(301)=>
      DANGLING(97), dataOut(300)=>DANGLING(98), dataOut(299)=>DANGLING(99), 
      dataOut(298)=>DANGLING(100), dataOut(297)=>DANGLING(101), dataOut(296)
      =>DANGLING(102), dataOut(295)=>DANGLING(103), dataOut(294)=>DANGLING(
      104), dataOut(293)=>DANGLING(105), dataOut(292)=>DANGLING(106), 
      dataOut(291)=>DANGLING(107), dataOut(290)=>DANGLING(108), dataOut(289)
      =>DANGLING(109), dataOut(288)=>DANGLING(110), dataOut(287)=>DANGLING(
      111), dataOut(286)=>DANGLING(112), dataOut(285)=>DANGLING(113), 
      dataOut(284)=>DANGLING(114), dataOut(283)=>DANGLING(115), dataOut(282)
      =>DANGLING(116), dataOut(281)=>DANGLING(117), dataOut(280)=>DANGLING(
      118), dataOut(279)=>DANGLING(119), dataOut(278)=>DANGLING(120), 
      dataOut(277)=>DANGLING(121), dataOut(276)=>DANGLING(122), dataOut(275)
      =>DANGLING(123), dataOut(274)=>DANGLING(124), dataOut(273)=>DANGLING(
      125), dataOut(272)=>DANGLING(126), dataOut(271)=>DANGLING(127), 
      dataOut(270)=>DANGLING(128), dataOut(269)=>DANGLING(129), dataOut(268)
      =>DANGLING(130), dataOut(267)=>DANGLING(131), dataOut(266)=>DANGLING(
      132), dataOut(265)=>DANGLING(133), dataOut(264)=>DANGLING(134), 
      dataOut(263)=>DANGLING(135), dataOut(262)=>DANGLING(136), dataOut(261)
      =>DANGLING(137), dataOut(260)=>DANGLING(138), dataOut(259)=>DANGLING(
      139), dataOut(258)=>DANGLING(140), dataOut(257)=>DANGLING(141), 
      dataOut(256)=>DANGLING(142), dataOut(255)=>DANGLING(143), dataOut(254)
      =>DANGLING(144), dataOut(253)=>DANGLING(145), dataOut(252)=>DANGLING(
      146), dataOut(251)=>DANGLING(147), dataOut(250)=>DANGLING(148), 
      dataOut(249)=>DANGLING(149), dataOut(248)=>DANGLING(150), dataOut(247)
      =>DANGLING(151), dataOut(246)=>DANGLING(152), dataOut(245)=>DANGLING(
      153), dataOut(244)=>DANGLING(154), dataOut(243)=>DANGLING(155), 
      dataOut(242)=>DANGLING(156), dataOut(241)=>DANGLING(157), dataOut(240)
      =>DANGLING(158), dataOut(239)=>DANGLING(159), dataOut(238)=>DANGLING(
      160), dataOut(237)=>DANGLING(161), dataOut(236)=>DANGLING(162), 
      dataOut(235)=>DANGLING(163), dataOut(234)=>DANGLING(164), dataOut(233)
      =>DANGLING(165), dataOut(232)=>DANGLING(166), dataOut(231)=>DANGLING(
      167), dataOut(230)=>DANGLING(168), dataOut(229)=>DANGLING(169), 
      dataOut(228)=>DANGLING(170), dataOut(227)=>DANGLING(171), dataOut(226)
      =>DANGLING(172), dataOut(225)=>DANGLING(173), dataOut(224)=>DANGLING(
      174), dataOut(223)=>DANGLING(175), dataOut(222)=>DANGLING(176), 
      dataOut(221)=>DANGLING(177), dataOut(220)=>DANGLING(178), dataOut(219)
      =>DANGLING(179), dataOut(218)=>DANGLING(180), dataOut(217)=>DANGLING(
      181), dataOut(216)=>DANGLING(182), dataOut(215)=>DANGLING(183), 
      dataOut(214)=>DANGLING(184), dataOut(213)=>DANGLING(185), dataOut(212)
      =>DANGLING(186), dataOut(211)=>DANGLING(187), dataOut(210)=>DANGLING(
      188), dataOut(209)=>DANGLING(189), dataOut(208)=>DANGLING(190), 
      dataOut(207)=>DANGLING(191), dataOut(206)=>DANGLING(192), dataOut(205)
      =>DANGLING(193), dataOut(204)=>DANGLING(194), dataOut(203)=>DANGLING(
      195), dataOut(202)=>DANGLING(196), dataOut(201)=>DANGLING(197), 
      dataOut(200)=>DANGLING(198), dataOut(199)=>DANGLING(199), dataOut(198)
      =>DANGLING(200), dataOut(197)=>DANGLING(201), dataOut(196)=>DANGLING(
      202), dataOut(195)=>DANGLING(203), dataOut(194)=>DANGLING(204), 
      dataOut(193)=>DANGLING(205), dataOut(192)=>DANGLING(206), dataOut(191)
      =>DANGLING(207), dataOut(190)=>DANGLING(208), dataOut(189)=>DANGLING(
      209), dataOut(188)=>DANGLING(210), dataOut(187)=>DANGLING(211), 
      dataOut(186)=>DANGLING(212), dataOut(185)=>DANGLING(213), dataOut(184)
      =>DANGLING(214), dataOut(183)=>DANGLING(215), dataOut(182)=>DANGLING(
      216), dataOut(181)=>DANGLING(217), dataOut(180)=>DANGLING(218), 
      dataOut(179)=>DANGLING(219), dataOut(178)=>DANGLING(220), dataOut(177)
      =>DANGLING(221), dataOut(176)=>DANGLING(222), dataOut(175)=>DANGLING(
      223), dataOut(174)=>DANGLING(224), dataOut(173)=>DANGLING(225), 
      dataOut(172)=>DANGLING(226), dataOut(171)=>DANGLING(227), dataOut(170)
      =>DANGLING(228), dataOut(169)=>DANGLING(229), dataOut(168)=>DANGLING(
      230), dataOut(167)=>DANGLING(231), dataOut(166)=>DANGLING(232), 
      dataOut(165)=>DANGLING(233), dataOut(164)=>DANGLING(234), dataOut(163)
      =>DANGLING(235), dataOut(162)=>DANGLING(236), dataOut(161)=>DANGLING(
      237), dataOut(160)=>DANGLING(238), dataOut(159)=>DANGLING(239), 
      dataOut(158)=>DANGLING(240), dataOut(157)=>DANGLING(241), dataOut(156)
      =>DANGLING(242), dataOut(155)=>DANGLING(243), dataOut(154)=>DANGLING(
      244), dataOut(153)=>DANGLING(245), dataOut(152)=>DANGLING(246), 
      dataOut(151)=>DANGLING(247), dataOut(150)=>DANGLING(248), dataOut(149)
      =>DANGLING(249), dataOut(148)=>DANGLING(250), dataOut(147)=>DANGLING(
      251), dataOut(146)=>DANGLING(252), dataOut(145)=>DANGLING(253), 
      dataOut(144)=>DANGLING(254), dataOut(143)=>DANGLING(255), dataOut(142)
      =>DANGLING(256), dataOut(141)=>DANGLING(257), dataOut(140)=>DANGLING(
      258), dataOut(139)=>DANGLING(259), dataOut(138)=>DANGLING(260), 
      dataOut(137)=>DANGLING(261), dataOut(136)=>DANGLING(262), dataOut(135)
      =>DANGLING(263), dataOut(134)=>DANGLING(264), dataOut(133)=>DANGLING(
      265), dataOut(132)=>DANGLING(266), dataOut(131)=>DANGLING(267), 
      dataOut(130)=>DANGLING(268), dataOut(129)=>DANGLING(269), dataOut(128)
      =>DANGLING(270), dataOut(127)=>DANGLING(271), dataOut(126)=>DANGLING(
      272), dataOut(125)=>DANGLING(273), dataOut(124)=>DANGLING(274), 
      dataOut(123)=>DANGLING(275), dataOut(122)=>DANGLING(276), dataOut(121)
      =>DANGLING(277), dataOut(120)=>DANGLING(278), dataOut(119)=>DANGLING(
      279), dataOut(118)=>DANGLING(280), dataOut(117)=>DANGLING(281), 
      dataOut(116)=>DANGLING(282), dataOut(115)=>DANGLING(283), dataOut(114)
      =>DANGLING(284), dataOut(113)=>DANGLING(285), dataOut(112)=>DANGLING(
      286), dataOut(111)=>DANGLING(287), dataOut(110)=>DANGLING(288), 
      dataOut(109)=>DANGLING(289), dataOut(108)=>DANGLING(290), dataOut(107)
      =>DANGLING(291), dataOut(106)=>DANGLING(292), dataOut(105)=>DANGLING(
      293), dataOut(104)=>DANGLING(294), dataOut(103)=>DANGLING(295), 
      dataOut(102)=>DANGLING(296), dataOut(101)=>DANGLING(297), dataOut(100)
      =>DANGLING(298), dataOut(99)=>DANGLING(299), dataOut(98)=>DANGLING(300
      ), dataOut(97)=>DANGLING(301), dataOut(96)=>DANGLING(302), dataOut(95)
      =>DANGLING(303), dataOut(94)=>DANGLING(304), dataOut(93)=>DANGLING(305
      ), dataOut(92)=>DANGLING(306), dataOut(91)=>DANGLING(307), dataOut(90)
      =>DANGLING(308), dataOut(89)=>DANGLING(309), dataOut(88)=>DANGLING(310
      ), dataOut(87)=>DANGLING(311), dataOut(86)=>DANGLING(312), dataOut(85)
      =>DANGLING(313), dataOut(84)=>DANGLING(314), dataOut(83)=>DANGLING(315
      ), dataOut(82)=>DANGLING(316), dataOut(81)=>DANGLING(317), dataOut(80)
      =>DANGLING(318), dataOut(79)=>DANGLING(319), dataOut(78)=>DANGLING(320
      ), dataOut(77)=>DANGLING(321), dataOut(76)=>DANGLING(322), dataOut(75)
      =>DANGLING(323), dataOut(74)=>DANGLING(324), dataOut(73)=>DANGLING(325
      ), dataOut(72)=>DANGLING(326), dataOut(71)=>DANGLING(327), dataOut(70)
      =>DANGLING(328), dataOut(69)=>DANGLING(329), dataOut(68)=>DANGLING(330
      ), dataOut(67)=>DANGLING(331), dataOut(66)=>DANGLING(332), dataOut(65)
      =>DANGLING(333), dataOut(64)=>DANGLING(334), dataOut(63)=>DANGLING(335
      ), dataOut(62)=>DANGLING(336), dataOut(61)=>DANGLING(337), dataOut(60)
      =>DANGLING(338), dataOut(59)=>DANGLING(339), dataOut(58)=>DANGLING(340
      ), dataOut(57)=>DANGLING(341), dataOut(56)=>DANGLING(342), dataOut(55)
      =>DANGLING(343), dataOut(54)=>DANGLING(344), dataOut(53)=>DANGLING(345
      ), dataOut(52)=>DANGLING(346), dataOut(51)=>DANGLING(347), dataOut(50)
      =>DANGLING(348), dataOut(49)=>DANGLING(349), dataOut(48)=>DANGLING(350
      ), dataOut(47)=>DANGLING(351), dataOut(46)=>DANGLING(352), dataOut(45)
      =>DANGLING(353), dataOut(44)=>DANGLING(354), dataOut(43)=>DANGLING(355
      ), dataOut(42)=>DANGLING(356), dataOut(41)=>DANGLING(357), dataOut(40)
      =>DANGLING(358), dataOut(39)=>DANGLING(359), dataOut(38)=>DANGLING(360
      ), dataOut(37)=>DANGLING(361), dataOut(36)=>DANGLING(362), dataOut(35)
      =>DANGLING(363), dataOut(34)=>DANGLING(364), dataOut(33)=>DANGLING(365
      ), dataOut(32)=>DANGLING(366), dataOut(31)=>DANGLING(367), dataOut(30)
      =>DANGLING(368), dataOut(29)=>DANGLING(369), dataOut(28)=>DANGLING(370
      ), dataOut(27)=>DANGLING(371), dataOut(26)=>DANGLING(372), dataOut(25)
      =>DANGLING(373), dataOut(24)=>DANGLING(374), dataOut(23)=>DANGLING(375
      ), dataOut(22)=>DANGLING(376), dataOut(21)=>DANGLING(377), dataOut(20)
      =>DANGLING(378), dataOut(19)=>DANGLING(379), dataOut(18)=>DANGLING(380
      ), dataOut(17)=>DANGLING(381), dataOut(16)=>DANGLING(382), dataOut(15)
      =>DANGLING(383), dataOut(14)=>DANGLING(384), dataOut(13)=>DANGLING(385
      ), dataOut(12)=>DANGLING(386), dataOut(11)=>DANGLING(387), dataOut(10)
      =>DANGLING(388), dataOut(9)=>DANGLING(389), dataOut(8)=>DANGLING(390), 
      dataOut(7)=>DANGLING(391), dataOut(6)=>DANGLING(392), dataOut(5)=>
      DANGLING(393), dataOut(4)=>DANGLING(394), dataOut(3)=>DANGLING(395), 
      dataOut(2)=>DANGLING(396), dataOut(1)=>DANGLING(397), dataOut(0)=>
      DANGLING(398), MFC=>ACKF, counterOut(3)=>DANGLING(399), counterOut(2)
      =>DANGLING(400), counterOut(1)=>DANGLING(401), counterOut(0)=>DANGLING
      (402));
   ImgMem : memoryDMA port map ( resetEN=>rst, AddressIn(12)=>AddressI_12, 
      AddressIn(11)=>AddressI_11, AddressIn(10)=>AddressI_10, AddressIn(9)=>
      AddressI_9, AddressIn(8)=>AddressI_8, AddressIn(7)=>AddressI_7, 
      AddressIn(6)=>AddressI_6, AddressIn(5)=>AddressI_5, AddressIn(4)=>
      AddressI_4, AddressIn(3)=>AddressI_3, AddressIn(2)=>AddressI_2, 
      AddressIn(1)=>AddressI_1, AddressIn(0)=>AddressI_0, dataIn(15)=>
      DataIIn_15, dataIn(14)=>DataIIn_14, dataIn(13)=>DataIIn_13, dataIn(12)
      =>DataIIn_12, dataIn(11)=>DataIIn_11, dataIn(10)=>DataIIn_10, 
      dataIn(9)=>DataIIn_9, dataIn(8)=>DataIIn_8, dataIn(7)=>DataIIn_7, 
      dataIn(6)=>DataIIn_6, dataIn(5)=>DataIIn_5, dataIn(4)=>DataIIn_4, 
      dataIn(3)=>DataIIn_3, dataIn(2)=>DataIIn_2, dataIn(1)=>DataIIn_1, 
      dataIn(0)=>DataIIn_0, switcherEN=>SwitchMEM_0, ramSelector=>
      ramSelector, readEn=>ReadI, writeEn=>WriteI, CLK=>nx10416, Normal=>
      zero_11, MFC=>ImgAddACKTriIN_0, counterOut(3)=>DANGLING(403), 
      counterOut(2)=>DANGLING(404), counterOut(1)=>DANGLING(405), 
      counterOut(0)=>DANGLING(406), dataOut(447)=>DataIOut_447, dataOut(446)
      =>DataIOut_446, dataOut(445)=>DataIOut_445, dataOut(444)=>DataIOut_444, 
      dataOut(443)=>DataIOut_443, dataOut(442)=>DataIOut_442, dataOut(441)=>
      DataIOut_441, dataOut(440)=>DataIOut_440, dataOut(439)=>DataIOut_439, 
      dataOut(438)=>DataIOut_438, dataOut(437)=>DataIOut_437, dataOut(436)=>
      DataIOut_436, dataOut(435)=>DataIOut_435, dataOut(434)=>DataIOut_434, 
      dataOut(433)=>DataIOut_433, dataOut(432)=>DataIOut_432, dataOut(431)=>
      DataIOut_431, dataOut(430)=>DataIOut_430, dataOut(429)=>DataIOut_429, 
      dataOut(428)=>DataIOut_428, dataOut(427)=>DataIOut_427, dataOut(426)=>
      DataIOut_426, dataOut(425)=>DataIOut_425, dataOut(424)=>DataIOut_424, 
      dataOut(423)=>DataIOut_423, dataOut(422)=>DataIOut_422, dataOut(421)=>
      DataIOut_421, dataOut(420)=>DataIOut_420, dataOut(419)=>DataIOut_419, 
      dataOut(418)=>DataIOut_418, dataOut(417)=>DataIOut_417, dataOut(416)=>
      DataIOut_416, dataOut(415)=>DataIOut_415, dataOut(414)=>DataIOut_414, 
      dataOut(413)=>DataIOut_413, dataOut(412)=>DataIOut_412, dataOut(411)=>
      DataIOut_411, dataOut(410)=>DataIOut_410, dataOut(409)=>DataIOut_409, 
      dataOut(408)=>DataIOut_408, dataOut(407)=>DataIOut_407, dataOut(406)=>
      DataIOut_406, dataOut(405)=>DataIOut_405, dataOut(404)=>DataIOut_404, 
      dataOut(403)=>DataIOut_403, dataOut(402)=>DataIOut_402, dataOut(401)=>
      DataIOut_401, dataOut(400)=>DataIOut_400, dataOut(399)=>DataIOut_399, 
      dataOut(398)=>DataIOut_398, dataOut(397)=>DataIOut_397, dataOut(396)=>
      DataIOut_396, dataOut(395)=>DataIOut_395, dataOut(394)=>DataIOut_394, 
      dataOut(393)=>DataIOut_393, dataOut(392)=>DataIOut_392, dataOut(391)=>
      DataIOut_391, dataOut(390)=>DataIOut_390, dataOut(389)=>DataIOut_389, 
      dataOut(388)=>DataIOut_388, dataOut(387)=>DataIOut_387, dataOut(386)=>
      DataIOut_386, dataOut(385)=>DataIOut_385, dataOut(384)=>DataIOut_384, 
      dataOut(383)=>DataIOut_383, dataOut(382)=>DataIOut_382, dataOut(381)=>
      DataIOut_381, dataOut(380)=>DataIOut_380, dataOut(379)=>DataIOut_379, 
      dataOut(378)=>DataIOut_378, dataOut(377)=>DataIOut_377, dataOut(376)=>
      DataIOut_376, dataOut(375)=>DataIOut_375, dataOut(374)=>DataIOut_374, 
      dataOut(373)=>DataIOut_373, dataOut(372)=>DataIOut_372, dataOut(371)=>
      DataIOut_371, dataOut(370)=>DataIOut_370, dataOut(369)=>DataIOut_369, 
      dataOut(368)=>DataIOut_368, dataOut(367)=>DataIOut_367, dataOut(366)=>
      DataIOut_366, dataOut(365)=>DataIOut_365, dataOut(364)=>DataIOut_364, 
      dataOut(363)=>DataIOut_363, dataOut(362)=>DataIOut_362, dataOut(361)=>
      DataIOut_361, dataOut(360)=>DataIOut_360, dataOut(359)=>DataIOut_359, 
      dataOut(358)=>DataIOut_358, dataOut(357)=>DataIOut_357, dataOut(356)=>
      DataIOut_356, dataOut(355)=>DataIOut_355, dataOut(354)=>DataIOut_354, 
      dataOut(353)=>DataIOut_353, dataOut(352)=>DataIOut_352, dataOut(351)=>
      DataIOut_351, dataOut(350)=>DataIOut_350, dataOut(349)=>DataIOut_349, 
      dataOut(348)=>DataIOut_348, dataOut(347)=>DataIOut_347, dataOut(346)=>
      DataIOut_346, dataOut(345)=>DataIOut_345, dataOut(344)=>DataIOut_344, 
      dataOut(343)=>DataIOut_343, dataOut(342)=>DataIOut_342, dataOut(341)=>
      DataIOut_341, dataOut(340)=>DataIOut_340, dataOut(339)=>DataIOut_339, 
      dataOut(338)=>DataIOut_338, dataOut(337)=>DataIOut_337, dataOut(336)=>
      DataIOut_336, dataOut(335)=>DataIOut_335, dataOut(334)=>DataIOut_334, 
      dataOut(333)=>DataIOut_333, dataOut(332)=>DataIOut_332, dataOut(331)=>
      DataIOut_331, dataOut(330)=>DataIOut_330, dataOut(329)=>DataIOut_329, 
      dataOut(328)=>DataIOut_328, dataOut(327)=>DataIOut_327, dataOut(326)=>
      DataIOut_326, dataOut(325)=>DataIOut_325, dataOut(324)=>DataIOut_324, 
      dataOut(323)=>DataIOut_323, dataOut(322)=>DataIOut_322, dataOut(321)=>
      DataIOut_321, dataOut(320)=>DataIOut_320, dataOut(319)=>DataIOut_319, 
      dataOut(318)=>DataIOut_318, dataOut(317)=>DataIOut_317, dataOut(316)=>
      DataIOut_316, dataOut(315)=>DataIOut_315, dataOut(314)=>DataIOut_314, 
      dataOut(313)=>DataIOut_313, dataOut(312)=>DataIOut_312, dataOut(311)=>
      DataIOut_311, dataOut(310)=>DataIOut_310, dataOut(309)=>DataIOut_309, 
      dataOut(308)=>DataIOut_308, dataOut(307)=>DataIOut_307, dataOut(306)=>
      DataIOut_306, dataOut(305)=>DataIOut_305, dataOut(304)=>DataIOut_304, 
      dataOut(303)=>DataIOut_303, dataOut(302)=>DataIOut_302, dataOut(301)=>
      DataIOut_301, dataOut(300)=>DataIOut_300, dataOut(299)=>DataIOut_299, 
      dataOut(298)=>DataIOut_298, dataOut(297)=>DataIOut_297, dataOut(296)=>
      DataIOut_296, dataOut(295)=>DataIOut_295, dataOut(294)=>DataIOut_294, 
      dataOut(293)=>DataIOut_293, dataOut(292)=>DataIOut_292, dataOut(291)=>
      DataIOut_291, dataOut(290)=>DataIOut_290, dataOut(289)=>DataIOut_289, 
      dataOut(288)=>DataIOut_288, dataOut(287)=>DataIOut_287, dataOut(286)=>
      DataIOut_286, dataOut(285)=>DataIOut_285, dataOut(284)=>DataIOut_284, 
      dataOut(283)=>DataIOut_283, dataOut(282)=>DataIOut_282, dataOut(281)=>
      DataIOut_281, dataOut(280)=>DataIOut_280, dataOut(279)=>DataIOut_279, 
      dataOut(278)=>DataIOut_278, dataOut(277)=>DataIOut_277, dataOut(276)=>
      DataIOut_276, dataOut(275)=>DataIOut_275, dataOut(274)=>DataIOut_274, 
      dataOut(273)=>DataIOut_273, dataOut(272)=>DataIOut_272, dataOut(271)=>
      DataIOut_271, dataOut(270)=>DataIOut_270, dataOut(269)=>DataIOut_269, 
      dataOut(268)=>DataIOut_268, dataOut(267)=>DataIOut_267, dataOut(266)=>
      DataIOut_266, dataOut(265)=>DataIOut_265, dataOut(264)=>DataIOut_264, 
      dataOut(263)=>DataIOut_263, dataOut(262)=>DataIOut_262, dataOut(261)=>
      DataIOut_261, dataOut(260)=>DataIOut_260, dataOut(259)=>DataIOut_259, 
      dataOut(258)=>DataIOut_258, dataOut(257)=>DataIOut_257, dataOut(256)=>
      DataIOut_256, dataOut(255)=>DataIOut_255, dataOut(254)=>DataIOut_254, 
      dataOut(253)=>DataIOut_253, dataOut(252)=>DataIOut_252, dataOut(251)=>
      DataIOut_251, dataOut(250)=>DataIOut_250, dataOut(249)=>DataIOut_249, 
      dataOut(248)=>DataIOut_248, dataOut(247)=>DataIOut_247, dataOut(246)=>
      DataIOut_246, dataOut(245)=>DataIOut_245, dataOut(244)=>DataIOut_244, 
      dataOut(243)=>DataIOut_243, dataOut(242)=>DataIOut_242, dataOut(241)=>
      DataIOut_241, dataOut(240)=>DataIOut_240, dataOut(239)=>DataIOut_239, 
      dataOut(238)=>DataIOut_238, dataOut(237)=>DataIOut_237, dataOut(236)=>
      DataIOut_236, dataOut(235)=>DataIOut_235, dataOut(234)=>DataIOut_234, 
      dataOut(233)=>DataIOut_233, dataOut(232)=>DataIOut_232, dataOut(231)=>
      DataIOut_231, dataOut(230)=>DataIOut_230, dataOut(229)=>DataIOut_229, 
      dataOut(228)=>DataIOut_228, dataOut(227)=>DataIOut_227, dataOut(226)=>
      DataIOut_226, dataOut(225)=>DataIOut_225, dataOut(224)=>DataIOut_224, 
      dataOut(223)=>DataIOut_223, dataOut(222)=>DataIOut_222, dataOut(221)=>
      DataIOut_221, dataOut(220)=>DataIOut_220, dataOut(219)=>DataIOut_219, 
      dataOut(218)=>DataIOut_218, dataOut(217)=>DataIOut_217, dataOut(216)=>
      DataIOut_216, dataOut(215)=>DataIOut_215, dataOut(214)=>DataIOut_214, 
      dataOut(213)=>DataIOut_213, dataOut(212)=>DataIOut_212, dataOut(211)=>
      DataIOut_211, dataOut(210)=>DataIOut_210, dataOut(209)=>DataIOut_209, 
      dataOut(208)=>DataIOut_208, dataOut(207)=>DataIOut_207, dataOut(206)=>
      DataIOut_206, dataOut(205)=>DataIOut_205, dataOut(204)=>DataIOut_204, 
      dataOut(203)=>DataIOut_203, dataOut(202)=>DataIOut_202, dataOut(201)=>
      DataIOut_201, dataOut(200)=>DataIOut_200, dataOut(199)=>DataIOut_199, 
      dataOut(198)=>DataIOut_198, dataOut(197)=>DataIOut_197, dataOut(196)=>
      DataIOut_196, dataOut(195)=>DataIOut_195, dataOut(194)=>DataIOut_194, 
      dataOut(193)=>DataIOut_193, dataOut(192)=>DataIOut_192, dataOut(191)=>
      DataIOut_191, dataOut(190)=>DataIOut_190, dataOut(189)=>DataIOut_189, 
      dataOut(188)=>DataIOut_188, dataOut(187)=>DataIOut_187, dataOut(186)=>
      DataIOut_186, dataOut(185)=>DataIOut_185, dataOut(184)=>DataIOut_184, 
      dataOut(183)=>DataIOut_183, dataOut(182)=>DataIOut_182, dataOut(181)=>
      DataIOut_181, dataOut(180)=>DataIOut_180, dataOut(179)=>DataIOut_179, 
      dataOut(178)=>DataIOut_178, dataOut(177)=>DataIOut_177, dataOut(176)=>
      DataIOut_176, dataOut(175)=>DataIOut_175, dataOut(174)=>DataIOut_174, 
      dataOut(173)=>DataIOut_173, dataOut(172)=>DataIOut_172, dataOut(171)=>
      DataIOut_171, dataOut(170)=>DataIOut_170, dataOut(169)=>DataIOut_169, 
      dataOut(168)=>DataIOut_168, dataOut(167)=>DataIOut_167, dataOut(166)=>
      DataIOut_166, dataOut(165)=>DataIOut_165, dataOut(164)=>DataIOut_164, 
      dataOut(163)=>DataIOut_163, dataOut(162)=>DataIOut_162, dataOut(161)=>
      DataIOut_161, dataOut(160)=>DataIOut_160, dataOut(159)=>DataIOut_159, 
      dataOut(158)=>DataIOut_158, dataOut(157)=>DataIOut_157, dataOut(156)=>
      DataIOut_156, dataOut(155)=>DataIOut_155, dataOut(154)=>DataIOut_154, 
      dataOut(153)=>DataIOut_153, dataOut(152)=>DataIOut_152, dataOut(151)=>
      DataIOut_151, dataOut(150)=>DataIOut_150, dataOut(149)=>DataIOut_149, 
      dataOut(148)=>DataIOut_148, dataOut(147)=>DataIOut_147, dataOut(146)=>
      DataIOut_146, dataOut(145)=>DataIOut_145, dataOut(144)=>DataIOut_144, 
      dataOut(143)=>DataIOut_143, dataOut(142)=>DataIOut_142, dataOut(141)=>
      DataIOut_141, dataOut(140)=>DataIOut_140, dataOut(139)=>DataIOut_139, 
      dataOut(138)=>DataIOut_138, dataOut(137)=>DataIOut_137, dataOut(136)=>
      DataIOut_136, dataOut(135)=>DataIOut_135, dataOut(134)=>DataIOut_134, 
      dataOut(133)=>DataIOut_133, dataOut(132)=>DataIOut_132, dataOut(131)=>
      DataIOut_131, dataOut(130)=>DataIOut_130, dataOut(129)=>DataIOut_129, 
      dataOut(128)=>DataIOut_128, dataOut(127)=>DataIOut_127, dataOut(126)=>
      DataIOut_126, dataOut(125)=>DataIOut_125, dataOut(124)=>DataIOut_124, 
      dataOut(123)=>DataIOut_123, dataOut(122)=>DataIOut_122, dataOut(121)=>
      DataIOut_121, dataOut(120)=>DataIOut_120, dataOut(119)=>DataIOut_119, 
      dataOut(118)=>DataIOut_118, dataOut(117)=>DataIOut_117, dataOut(116)=>
      DataIOut_116, dataOut(115)=>DataIOut_115, dataOut(114)=>DataIOut_114, 
      dataOut(113)=>DataIOut_113, dataOut(112)=>DataIOut_112, dataOut(111)=>
      DataIOut_111, dataOut(110)=>DataIOut_110, dataOut(109)=>DataIOut_109, 
      dataOut(108)=>DataIOut_108, dataOut(107)=>DataIOut_107, dataOut(106)=>
      DataIOut_106, dataOut(105)=>DataIOut_105, dataOut(104)=>DataIOut_104, 
      dataOut(103)=>DataIOut_103, dataOut(102)=>DataIOut_102, dataOut(101)=>
      DataIOut_101, dataOut(100)=>DataIOut_100, dataOut(99)=>DataIOut_99, 
      dataOut(98)=>DataIOut_98, dataOut(97)=>DataIOut_97, dataOut(96)=>
      DataIOut_96, dataOut(95)=>DataIOut_95, dataOut(94)=>DataIOut_94, 
      dataOut(93)=>DataIOut_93, dataOut(92)=>DataIOut_92, dataOut(91)=>
      DataIOut_91, dataOut(90)=>DataIOut_90, dataOut(89)=>DataIOut_89, 
      dataOut(88)=>DataIOut_88, dataOut(87)=>DataIOut_87, dataOut(86)=>
      DataIOut_86, dataOut(85)=>DataIOut_85, dataOut(84)=>DataIOut_84, 
      dataOut(83)=>DataIOut_83, dataOut(82)=>DataIOut_82, dataOut(81)=>
      DataIOut_81, dataOut(80)=>DataIOut_80, dataOut(79)=>DataIOut_79, 
      dataOut(78)=>DataIOut_78, dataOut(77)=>DataIOut_77, dataOut(76)=>
      DataIOut_76, dataOut(75)=>DataIOut_75, dataOut(74)=>DataIOut_74, 
      dataOut(73)=>DataIOut_73, dataOut(72)=>DataIOut_72, dataOut(71)=>
      DataIOut_71, dataOut(70)=>DataIOut_70, dataOut(69)=>DataIOut_69, 
      dataOut(68)=>DataIOut_68, dataOut(67)=>DataIOut_67, dataOut(66)=>
      DataIOut_66, dataOut(65)=>DataIOut_65, dataOut(64)=>DataIOut_64, 
      dataOut(63)=>DataIOut_63, dataOut(62)=>DataIOut_62, dataOut(61)=>
      DataIOut_61, dataOut(60)=>DataIOut_60, dataOut(59)=>DataIOut_59, 
      dataOut(58)=>DataIOut_58, dataOut(57)=>DataIOut_57, dataOut(56)=>
      DataIOut_56, dataOut(55)=>DataIOut_55, dataOut(54)=>DataIOut_54, 
      dataOut(53)=>DataIOut_53, dataOut(52)=>DataIOut_52, dataOut(51)=>
      DataIOut_51, dataOut(50)=>DataIOut_50, dataOut(49)=>DataIOut_49, 
      dataOut(48)=>DataIOut_48, dataOut(47)=>DataIOut_47, dataOut(46)=>
      DataIOut_46, dataOut(45)=>DataIOut_45, dataOut(44)=>DataIOut_44, 
      dataOut(43)=>DataIOut_43, dataOut(42)=>DataIOut_42, dataOut(41)=>
      DataIOut_41, dataOut(40)=>DataIOut_40, dataOut(39)=>DataIOut_39, 
      dataOut(38)=>DataIOut_38, dataOut(37)=>DataIOut_37, dataOut(36)=>
      DataIOut_36, dataOut(35)=>DataIOut_35, dataOut(34)=>DataIOut_34, 
      dataOut(33)=>DataIOut_33, dataOut(32)=>DataIOut_32, dataOut(31)=>
      DataIOut_31, dataOut(30)=>DataIOut_30, dataOut(29)=>DataIOut_29, 
      dataOut(28)=>DataIOut_28, dataOut(27)=>DataIOut_27, dataOut(26)=>
      DataIOut_26, dataOut(25)=>DataIOut_25, dataOut(24)=>DataIOut_24, 
      dataOut(23)=>DataIOut_23, dataOut(22)=>DataIOut_22, dataOut(21)=>
      DataIOut_21, dataOut(20)=>DataIOut_20, dataOut(19)=>DataIOut_19, 
      dataOut(18)=>DataIOut_18, dataOut(17)=>DataIOut_17, dataOut(16)=>
      DataIOut_16, dataOut(15)=>DataIOut_15, dataOut(14)=>DataIOut_14, 
      dataOut(13)=>DataIOut_13, dataOut(12)=>DataIOut_12, dataOut(11)=>
      DataIOut_11, dataOut(10)=>DataIOut_10, dataOut(9)=>DataIOut_9, 
      dataOut(8)=>DataIOut_8, dataOut(7)=>DataIOut_7, dataOut(6)=>DataIOut_6, 
      dataOut(5)=>DataIOut_5, dataOut(4)=>DataIOut_4, dataOut(3)=>DataIOut_3, 
      dataOut(2)=>DataIOut_2, dataOut(1)=>DataIOut_1, dataOut(0)=>DataIOut_0
   );
   ReadInf : ReadInfoState port map ( CLK=>nx10418, S(14)=>zero_11, S(13)=>
      zero_11, S(12)=>zero_11, S(11)=>zero_11, S(10)=>zero_11, S(9)=>zero_11, 
      S(8)=>zero_11, S(7)=>zero_11, S(6)=>zero_11, S(5)=>zero_11, S(4)=>
      zero_11, S(3)=>zero_11, S(2)=>zero_11, S(1)=>zero_11, S(0)=>
      current_state_0, reset=>rst, MFC=>zero_11, filterAddressReg_out(12)=>
      nx9974, filterAddressReg_out(11)=>nx9978, filterAddressReg_out(10)=>
      nx9982, filterAddressReg_out(9)=>nx9986, filterAddressReg_out(8)=>
      nx9990, filterAddressReg_out(7)=>nx9994, filterAddressReg_out(6)=>
      nx9998, filterAddressReg_out(5)=>nx10002, filterAddressReg_out(4)=>
      nx10006, filterAddressReg_out(3)=>nx10010, filterAddressReg_out(2)=>
      nx10014, filterAddressReg_out(1)=>nx10018, filterAddressReg_out(0)=>
      nx10022, filterRamData(15)=>nx10256, filterRamData(14)=>nx10262, 
      filterRamData(13)=>nx10268, filterRamData(12)=>nx10274, 
      filterRamData(11)=>nx10280, filterRamData(10)=>nx10286, 
      filterRamData(9)=>nx10292, filterRamData(8)=>nx10292, filterRamData(7)
      =>nx10294, filterRamData(6)=>nx10294, filterRamData(5)=>nx10296, 
      filterRamData(4)=>nx10298, filterRamData(3)=>nx10300, filterRamData(2)
      =>nx10302, filterRamData(1)=>nx10302, filterRamData(0)=>nx10304, 
      noOfLayersReg_out(15)=>DANGLING(407), noOfLayersReg_out(14)=>DANGLING(
      408), noOfLayersReg_out(13)=>DANGLING(409), noOfLayersReg_out(12)=>
      DANGLING(410), noOfLayersReg_out(11)=>DANGLING(411), 
      noOfLayersReg_out(10)=>DANGLING(412), noOfLayersReg_out(9)=>DANGLING(
      413), noOfLayersReg_out(8)=>DANGLING(414), noOfLayersReg_out(7)=>
      DANGLING(415), noOfLayersReg_out(6)=>DANGLING(416), 
      noOfLayersReg_out(5)=>DANGLING(417), noOfLayersReg_out(4)=>DANGLING(
      418), noOfLayersReg_out(3)=>DANGLING(419), noOfLayersReg_out(2)=>
      DANGLING(420), noOfLayersReg_out(1)=>NoOfLayers_1, 
      noOfLayersReg_out(0)=>NoOfLayers_0, filterRamAddress(12)=>AddressF_12, 
      filterRamAddress(11)=>AddressF_11, filterRamAddress(10)=>AddressF_10, 
      filterRamAddress(9)=>AddressF_9, filterRamAddress(8)=>AddressF_8, 
      filterRamAddress(7)=>AddressF_7, filterRamAddress(6)=>AddressF_6, 
      filterRamAddress(5)=>AddressF_5, filterRamAddress(4)=>AddressF_4, 
      filterRamAddress(3)=>AddressF_3, filterRamAddress(2)=>AddressF_2, 
      filterRamAddress(1)=>AddressF_1, filterRamAddress(0)=>AddressF_0);
   FilterAddress : nBitRegister_13 port map ( D(12)=>FilterAddressIN_12, 
      D(11)=>FilterAddressIN_11, D(10)=>FilterAddressIN_10, D(9)=>
      FilterAddressIN_9, D(8)=>FilterAddressIN_8, D(7)=>FilterAddressIN_7, 
      D(6)=>FilterAddressIN_6, D(5)=>FilterAddressIN_5, D(4)=>
      FilterAddressIN_4, D(3)=>FilterAddressIN_3, D(2)=>FilterAddressIN_2, 
      D(1)=>FilterAddressIN_1, D(0)=>FilterAddressIN_0, CLK=>nx10414, RST=>
      rst, EN=>FilterAddressEN, Q(12)=>FilterAddressOut_12, Q(11)=>
      FilterAddressOut_11, Q(10)=>FilterAddressOut_10, Q(9)=>
      FilterAddressOut_9, Q(8)=>FilterAddressOut_8, Q(7)=>FilterAddressOut_7, 
      Q(6)=>FilterAddressOut_6, Q(5)=>FilterAddressOut_5, Q(4)=>
      FilterAddressOut_4, Q(3)=>FilterAddressOut_3, Q(2)=>FilterAddressOut_2, 
      Q(1)=>FilterAddressOut_1, Q(0)=>FilterAddressOut_0);
   AdderTryState : triStateBuffer_13 port map ( D(12)=>TriStateCounterOUT_12, 
      D(11)=>TriStateCounterOUT_11, D(10)=>TriStateCounterOUT_10, D(9)=>
      TriStateCounterOUT_9, D(8)=>TriStateCounterOUT_8, D(7)=>
      TriStateCounterOUT_7, D(6)=>TriStateCounterOUT_6, D(5)=>
      TriStateCounterOUT_5, D(4)=>TriStateCounterOUT_4, D(3)=>
      TriStateCounterOUT_3, D(2)=>TriStateCounterOUT_2, D(1)=>
      TriStateCounterOUT_1, D(0)=>TriStateCounterOUT_0, EN=>
      TriStateCounterEN, F(12)=>FilterAddressIN_12, F(11)=>
      FilterAddressIN_11, F(10)=>FilterAddressIN_10, F(9)=>FilterAddressIN_9, 
      F(8)=>FilterAddressIN_8, F(7)=>FilterAddressIN_7, F(6)=>
      FilterAddressIN_6, F(5)=>FilterAddressIN_5, F(4)=>FilterAddressIN_4, 
      F(3)=>FilterAddressIN_3, F(2)=>FilterAddressIN_2, F(1)=>
      FilterAddressIN_1, F(0)=>FilterAddressIN_0);
   FilterAddressAdder : my_nadder_13 port map ( a(12)=>nx9974, a(11)=>nx9978, 
      a(10)=>nx9982, a(9)=>nx9986, a(8)=>nx9990, a(7)=>nx9994, a(6)=>nx9998, 
      a(5)=>nx10002, a(4)=>nx10006, a(3)=>nx10010, a(2)=>nx10014, a(1)=>
      nx10018, a(0)=>nx10022, b(12)=>zero_11, b(11)=>zero_11, b(10)=>zero_11, 
      b(9)=>zero_11, b(8)=>zero_11, b(7)=>zero_11, b(6)=>zero_11, b(5)=>
      zero_11, b(4)=>zero_11, b(3)=>zero_11, b(2)=>zero_11, b(1)=>zero_11, 
      b(0)=>zero_11, cin=>PWR, s(12)=>TriStateCounterOUT_12, s(11)=>
      TriStateCounterOUT_11, s(10)=>TriStateCounterOUT_10, s(9)=>
      TriStateCounterOUT_9, s(8)=>TriStateCounterOUT_8, s(7)=>
      TriStateCounterOUT_7, s(6)=>TriStateCounterOUT_6, s(5)=>
      TriStateCounterOUT_5, s(4)=>TriStateCounterOUT_4, s(3)=>
      TriStateCounterOUT_3, s(2)=>TriStateCounterOUT_2, s(1)=>
      TriStateCounterOUT_1, s(0)=>TriStateCounterOUT_0, cout=>DANGLING(421)
   );
   ImgAddReg : nBitRegister_13 port map ( D(12)=>ImgAddRegIN_12, D(11)=>
      ImgAddRegIN_11, D(10)=>ImgAddRegIN_10, D(9)=>ImgAddRegIN_9, D(8)=>
      ImgAddRegIN_8, D(7)=>ImgAddRegIN_7, D(6)=>ImgAddRegIN_6, D(5)=>
      ImgAddRegIN_5, D(4)=>ImgAddRegIN_4, D(3)=>ImgAddRegIN_3, D(2)=>
      ImgAddRegIN_2, D(1)=>ImgAddRegIN_1, D(0)=>ImgAddRegIN_0, CLK=>nx10418, 
      RST=>ImgAddRST, EN=>ImgAddRegEN, Q(12)=>ImgAddRegOut_12, Q(11)=>
      ImgAddRegOut_11, Q(10)=>ImgAddRegOut_10, Q(9)=>ImgAddRegOut_9, Q(8)=>
      ImgAddRegOut_8, Q(7)=>ImgAddRegOut_7, Q(6)=>ImgAddRegOut_6, Q(5)=>
      ImgAddRegOut_5, Q(4)=>ImgAddRegOut_4, Q(3)=>ImgAddRegOut_3, Q(2)=>
      ImgAddRegOut_2, Q(1)=>ImgAddRegOut_1, Q(0)=>ImgAddRegOut_0);
   ImgAddACKTri : triStateBuffer_13 port map ( D(12)=>zero_11, D(11)=>
      zero_11, D(10)=>zero_11, D(9)=>zero_11, D(8)=>zero_11, D(7)=>zero_11, 
      D(6)=>zero_11, D(5)=>zero_11, D(4)=>zero_11, D(3)=>zero_11, D(2)=>
      zero_11, D(1)=>zero_11, D(0)=>nx10026, EN=>nx9972, F(12)=>
      ImgAddRegIN_12, F(11)=>ImgAddRegIN_11, F(10)=>ImgAddRegIN_10, F(9)=>
      ImgAddRegIN_9, F(8)=>ImgAddRegIN_8, F(7)=>ImgAddRegIN_7, F(6)=>
      ImgAddRegIN_6, F(5)=>ImgAddRegIN_5, F(4)=>ImgAddRegIN_4, F(3)=>
      ImgAddRegIN_3, F(2)=>ImgAddRegIN_2, F(1)=>ImgAddRegIN_1, F(0)=>
      ImgAddRegIN_0);
   ReadLayerInfo_EXMPLR : ReadLayerInfo port map ( LayerInfoIn(15)=>nx10258, 
      LayerInfoIn(14)=>nx10264, LayerInfoIn(13)=>nx10270, LayerInfoIn(12)=>
      nx10276, LayerInfoIn(11)=>nx10282, LayerInfoIn(10)=>nx10288, 
      LayerInfoIn(9)=>nx10292, LayerInfoIn(8)=>nx10292, LayerInfoIn(7)=>
      nx10294, LayerInfoIn(6)=>nx10296, LayerInfoIn(5)=>nx10298, 
      LayerInfoIn(4)=>nx10298, LayerInfoIn(3)=>nx10300, LayerInfoIn(2)=>
      nx10302, LayerInfoIn(1)=>nx10302, LayerInfoIn(0)=>nx10304, 
      ImgWidthIn(15)=>nx10312, ImgWidthIn(14)=>nx10316, ImgWidthIn(13)=>
      nx10320, ImgWidthIn(12)=>nx10324, ImgWidthIn(11)=>nx10328, 
      ImgWidthIn(10)=>nx10332, ImgWidthIn(9)=>nx10336, ImgWidthIn(8)=>
      nx10340, ImgWidthIn(7)=>nx10344, ImgWidthIn(6)=>nx10348, ImgWidthIn(5)
      =>nx10352, ImgWidthIn(4)=>nx10356, ImgWidthIn(3)=>nx10360, 
      ImgWidthIn(2)=>nx10364, ImgWidthIn(1)=>nx10368, ImgWidthIn(0)=>nx10372, 
      FilterAdd(12)=>nx9974, FilterAdd(11)=>nx9978, FilterAdd(10)=>nx9982, 
      FilterAdd(9)=>nx9986, FilterAdd(8)=>nx9990, FilterAdd(7)=>nx9994, 
      FilterAdd(6)=>nx9998, FilterAdd(5)=>nx10002, FilterAdd(4)=>nx10006, 
      FilterAdd(3)=>nx10010, FilterAdd(2)=>nx10014, FilterAdd(1)=>nx10018, 
      FilterAdd(0)=>nx10022, ImgAdd(12)=>ImgAddRegOut_12, ImgAdd(11)=>
      ImgAddRegOut_11, ImgAdd(10)=>ImgAddRegOut_10, ImgAdd(9)=>
      ImgAddRegOut_9, ImgAdd(8)=>ImgAddRegOut_8, ImgAdd(7)=>ImgAddRegOut_7, 
      ImgAdd(6)=>ImgAddRegOut_6, ImgAdd(5)=>ImgAddRegOut_5, ImgAdd(4)=>
      ImgAddRegOut_4, ImgAdd(3)=>ImgAddRegOut_3, ImgAdd(2)=>ImgAddRegOut_2, 
      ImgAdd(1)=>ImgAddRegOut_1, ImgAdd(0)=>ImgAddRegOut_0, clk=>nx10420, 
      rst=>rst, ACKF=>nx10308, ACKI=>nx10026, current_state(14)=>zero_11, 
      current_state(13)=>zero_11, current_state(12)=>zero_11, 
      current_state(11)=>zero_11, current_state(10)=>zero_11, 
      current_state(9)=>zero_11, current_state(8)=>zero_11, current_state(7)
      =>zero_11, current_state(6)=>zero_11, current_state(5)=>zero_11, 
      current_state(4)=>zero_11, current_state(3)=>zero_11, current_state(2)
      =>zero_11, current_state(1)=>nx9970, current_state(0)=>zero_11, 
      LayerInfoOut(15)=>LayerInfoOut_15, LayerInfoOut(14)=>LayerInfoOut_14, 
      LayerInfoOut(13)=>DANGLING(422), LayerInfoOut(12)=>LayerInfoOut_12, 
      LayerInfoOut(11)=>LayerInfoOut_11, LayerInfoOut(10)=>LayerInfoOut_10, 
      LayerInfoOut(9)=>LayerInfoOut_9, LayerInfoOut(8)=>LayerInfoOut_8, 
      LayerInfoOut(7)=>LayerInfoOut_7, LayerInfoOut(6)=>LayerInfoOut_6, 
      LayerInfoOut(5)=>LayerInfoOut_5, LayerInfoOut(4)=>LayerInfoOut_4, 
      LayerInfoOut(3)=>LayerInfoOut_3, LayerInfoOut(2)=>LayerInfoOut_2, 
      LayerInfoOut(1)=>LayerInfoOut_1, LayerInfoOut(0)=>LayerInfoOut_0, 
      ImgWidthOut(15)=>ImgWidthOut_15, ImgWidthOut(14)=>ImgWidthOut_14, 
      ImgWidthOut(13)=>ImgWidthOut_13, ImgWidthOut(12)=>ImgWidthOut_12, 
      ImgWidthOut(11)=>ImgWidthOut_11, ImgWidthOut(10)=>ImgWidthOut_10, 
      ImgWidthOut(9)=>ImgWidthOut_9, ImgWidthOut(8)=>ImgWidthOut_8, 
      ImgWidthOut(7)=>ImgWidthOut_7, ImgWidthOut(6)=>ImgWidthOut_6, 
      ImgWidthOut(5)=>ImgWidthOut_5, ImgWidthOut(4)=>ImgWidthOut_4, 
      ImgWidthOut(3)=>ImgWidthOut_3, ImgWidthOut(2)=>ImgWidthOut_2, 
      ImgWidthOut(1)=>ImgWidthOut_1, ImgWidthOut(0)=>ImgWidthOut_0, 
      FilterAddToDMA(12)=>AddressF_12, FilterAddToDMA(11)=>AddressF_11, 
      FilterAddToDMA(10)=>AddressF_10, FilterAddToDMA(9)=>AddressF_9, 
      FilterAddToDMA(8)=>AddressF_8, FilterAddToDMA(7)=>AddressF_7, 
      FilterAddToDMA(6)=>AddressF_6, FilterAddToDMA(5)=>AddressF_5, 
      FilterAddToDMA(4)=>AddressF_4, FilterAddToDMA(3)=>AddressF_3, 
      FilterAddToDMA(2)=>AddressF_2, FilterAddToDMA(1)=>AddressF_1, 
      FilterAddToDMA(0)=>AddressF_0, ImgAddToDMA(12)=>AddressI_12, 
      ImgAddToDMA(11)=>AddressI_11, ImgAddToDMA(10)=>AddressI_10, 
      ImgAddToDMA(9)=>AddressI_9, ImgAddToDMA(8)=>AddressI_8, ImgAddToDMA(7)
      =>AddressI_7, ImgAddToDMA(6)=>AddressI_6, ImgAddToDMA(5)=>AddressI_5, 
      ImgAddToDMA(4)=>AddressI_4, ImgAddToDMA(3)=>AddressI_3, ImgAddToDMA(2)
      =>AddressI_2, ImgAddToDMA(1)=>AddressI_1, ImgAddToDMA(0)=>AddressI_0);
   ClacInfo : CalculateInfo port map ( WSquareOut(9)=>WidthSquareOut_9, 
      WSquareOut(8)=>WidthSquareOut_8, WSquareOut(7)=>WidthSquareOut_7, 
      WSquareOut(6)=>WidthSquareOut_6, WSquareOut(5)=>WidthSquareOut_5, 
      WSquareOut(4)=>WidthSquareOut_4, WSquareOut(3)=>WidthSquareOut_3, 
      WSquareOut(2)=>WidthSquareOut_2, WSquareOut(1)=>WidthSquareOut_1, 
      WSquareOut(0)=>WidthSquareOut_0, CounOut(1)=>DANGLING(423), CounOut(0)
      =>DANGLING(424), LayerInfoIn(15)=>zero_11, LayerInfoIn(14)=>zero_11, 
      LayerInfoIn(13)=>zero_11, LayerInfoIn(12)=>zero_11, LayerInfoIn(11)=>
      zero_11, LayerInfoIn(10)=>zero_11, LayerInfoIn(9)=>zero_11, 
      LayerInfoIn(8)=>nx10376, LayerInfoIn(7)=>nx10380, LayerInfoIn(6)=>
      nx10384, LayerInfoIn(5)=>nx10388, LayerInfoIn(4)=>nx10392, 
      LayerInfoIn(3)=>zero_11, LayerInfoIn(2)=>zero_11, LayerInfoIn(1)=>
      zero_11, LayerInfoIn(0)=>zero_11, clk=>nx10504, rst=>rst, 
      current_state(14)=>zero_11, current_state(13)=>zero_11, 
      current_state(12)=>zero_11, current_state(11)=>zero_11, 
      current_state(10)=>zero_11, current_state(9)=>zero_11, 
      current_state(8)=>zero_11, current_state(7)=>zero_11, current_state(6)
      =>zero_11, current_state(5)=>zero_11, current_state(4)=>nx9966, 
      current_state(3)=>zero_11, current_state(2)=>current_state_2, 
      current_state(1)=>zero_11, current_state(0)=>zero_11, ACK=>DANGLING(
      425), ACKI=>nx10026, Wmin1(4)=>DANGLING(426), Wmin1(3)=>DANGLING(427), 
      Wmin1(2)=>DANGLING(428), Wmin1(1)=>DANGLING(429), Wmin1(0)=>DANGLING(
      430));
   RBias : ReadBias port map ( current_state(14)=>zero_11, current_state(13)
      =>zero_11, current_state(12)=>zero_11, current_state(11)=>zero_11, 
      current_state(10)=>zero_11, current_state(9)=>zero_11, 
      current_state(8)=>zero_11, current_state(7)=>zero_11, current_state(6)
      =>zero_11, current_state(5)=>zero_11, current_state(4)=>nx9968, 
      current_state(3)=>zero_11, current_state(2)=>zero_11, current_state(1)
      =>zero_11, current_state(0)=>zero_11, BIAS(399)=>zero_11, BIAS(398)=>
      zero_11, BIAS(397)=>zero_11, BIAS(396)=>zero_11, BIAS(395)=>zero_11, 
      BIAS(394)=>zero_11, BIAS(393)=>zero_11, BIAS(392)=>zero_11, BIAS(391)
      =>zero_11, BIAS(390)=>zero_11, BIAS(389)=>zero_11, BIAS(388)=>zero_11, 
      BIAS(387)=>zero_11, BIAS(386)=>zero_11, BIAS(385)=>zero_11, BIAS(384)
      =>zero_11, BIAS(383)=>zero_11, BIAS(382)=>zero_11, BIAS(381)=>zero_11, 
      BIAS(380)=>zero_11, BIAS(379)=>zero_11, BIAS(378)=>zero_11, BIAS(377)
      =>zero_11, BIAS(376)=>zero_11, BIAS(375)=>zero_11, BIAS(374)=>zero_11, 
      BIAS(373)=>zero_11, BIAS(372)=>zero_11, BIAS(371)=>zero_11, BIAS(370)
      =>zero_11, BIAS(369)=>zero_11, BIAS(368)=>zero_11, BIAS(367)=>zero_11, 
      BIAS(366)=>zero_11, BIAS(365)=>zero_11, BIAS(364)=>zero_11, BIAS(363)
      =>zero_11, BIAS(362)=>zero_11, BIAS(361)=>zero_11, BIAS(360)=>zero_11, 
      BIAS(359)=>zero_11, BIAS(358)=>zero_11, BIAS(357)=>zero_11, BIAS(356)
      =>zero_11, BIAS(355)=>zero_11, BIAS(354)=>zero_11, BIAS(353)=>zero_11, 
      BIAS(352)=>zero_11, BIAS(351)=>zero_11, BIAS(350)=>zero_11, BIAS(349)
      =>zero_11, BIAS(348)=>zero_11, BIAS(347)=>zero_11, BIAS(346)=>zero_11, 
      BIAS(345)=>zero_11, BIAS(344)=>zero_11, BIAS(343)=>zero_11, BIAS(342)
      =>zero_11, BIAS(341)=>zero_11, BIAS(340)=>zero_11, BIAS(339)=>zero_11, 
      BIAS(338)=>zero_11, BIAS(337)=>zero_11, BIAS(336)=>zero_11, BIAS(335)
      =>zero_11, BIAS(334)=>zero_11, BIAS(333)=>zero_11, BIAS(332)=>zero_11, 
      BIAS(331)=>zero_11, BIAS(330)=>zero_11, BIAS(329)=>zero_11, BIAS(328)
      =>zero_11, BIAS(327)=>zero_11, BIAS(326)=>zero_11, BIAS(325)=>zero_11, 
      BIAS(324)=>zero_11, BIAS(323)=>zero_11, BIAS(322)=>zero_11, BIAS(321)
      =>zero_11, BIAS(320)=>zero_11, BIAS(319)=>zero_11, BIAS(318)=>zero_11, 
      BIAS(317)=>zero_11, BIAS(316)=>zero_11, BIAS(315)=>zero_11, BIAS(314)
      =>zero_11, BIAS(313)=>zero_11, BIAS(312)=>zero_11, BIAS(311)=>zero_11, 
      BIAS(310)=>zero_11, BIAS(309)=>zero_11, BIAS(308)=>zero_11, BIAS(307)
      =>zero_11, BIAS(306)=>zero_11, BIAS(305)=>zero_11, BIAS(304)=>zero_11, 
      BIAS(303)=>zero_11, BIAS(302)=>zero_11, BIAS(301)=>zero_11, BIAS(300)
      =>zero_11, BIAS(299)=>zero_11, BIAS(298)=>zero_11, BIAS(297)=>zero_11, 
      BIAS(296)=>zero_11, BIAS(295)=>zero_11, BIAS(294)=>zero_11, BIAS(293)
      =>zero_11, BIAS(292)=>zero_11, BIAS(291)=>zero_11, BIAS(290)=>zero_11, 
      BIAS(289)=>zero_11, BIAS(288)=>zero_11, BIAS(287)=>zero_11, BIAS(286)
      =>zero_11, BIAS(285)=>zero_11, BIAS(284)=>zero_11, BIAS(283)=>zero_11, 
      BIAS(282)=>zero_11, BIAS(281)=>zero_11, BIAS(280)=>zero_11, BIAS(279)
      =>zero_11, BIAS(278)=>zero_11, BIAS(277)=>zero_11, BIAS(276)=>zero_11, 
      BIAS(275)=>zero_11, BIAS(274)=>zero_11, BIAS(273)=>zero_11, BIAS(272)
      =>zero_11, BIAS(271)=>zero_11, BIAS(270)=>zero_11, BIAS(269)=>zero_11, 
      BIAS(268)=>zero_11, BIAS(267)=>zero_11, BIAS(266)=>zero_11, BIAS(265)
      =>zero_11, BIAS(264)=>zero_11, BIAS(263)=>zero_11, BIAS(262)=>zero_11, 
      BIAS(261)=>zero_11, BIAS(260)=>zero_11, BIAS(259)=>zero_11, BIAS(258)
      =>zero_11, BIAS(257)=>zero_11, BIAS(256)=>zero_11, BIAS(255)=>zero_11, 
      BIAS(254)=>zero_11, BIAS(253)=>zero_11, BIAS(252)=>zero_11, BIAS(251)
      =>zero_11, BIAS(250)=>zero_11, BIAS(249)=>zero_11, BIAS(248)=>zero_11, 
      BIAS(247)=>zero_11, BIAS(246)=>zero_11, BIAS(245)=>zero_11, BIAS(244)
      =>zero_11, BIAS(243)=>zero_11, BIAS(242)=>zero_11, BIAS(241)=>zero_11, 
      BIAS(240)=>zero_11, BIAS(239)=>zero_11, BIAS(238)=>zero_11, BIAS(237)
      =>zero_11, BIAS(236)=>zero_11, BIAS(235)=>zero_11, BIAS(234)=>zero_11, 
      BIAS(233)=>zero_11, BIAS(232)=>zero_11, BIAS(231)=>zero_11, BIAS(230)
      =>zero_11, BIAS(229)=>zero_11, BIAS(228)=>zero_11, BIAS(227)=>zero_11, 
      BIAS(226)=>zero_11, BIAS(225)=>zero_11, BIAS(224)=>zero_11, BIAS(223)
      =>zero_11, BIAS(222)=>zero_11, BIAS(221)=>zero_11, BIAS(220)=>zero_11, 
      BIAS(219)=>zero_11, BIAS(218)=>zero_11, BIAS(217)=>zero_11, BIAS(216)
      =>zero_11, BIAS(215)=>zero_11, BIAS(214)=>zero_11, BIAS(213)=>zero_11, 
      BIAS(212)=>zero_11, BIAS(211)=>zero_11, BIAS(210)=>zero_11, BIAS(209)
      =>zero_11, BIAS(208)=>zero_11, BIAS(207)=>zero_11, BIAS(206)=>zero_11, 
      BIAS(205)=>zero_11, BIAS(204)=>zero_11, BIAS(203)=>zero_11, BIAS(202)
      =>zero_11, BIAS(201)=>zero_11, BIAS(200)=>zero_11, BIAS(199)=>zero_11, 
      BIAS(198)=>zero_11, BIAS(197)=>zero_11, BIAS(196)=>zero_11, BIAS(195)
      =>zero_11, BIAS(194)=>zero_11, BIAS(193)=>zero_11, BIAS(192)=>zero_11, 
      BIAS(191)=>zero_11, BIAS(190)=>zero_11, BIAS(189)=>zero_11, BIAS(188)
      =>zero_11, BIAS(187)=>zero_11, BIAS(186)=>zero_11, BIAS(185)=>zero_11, 
      BIAS(184)=>zero_11, BIAS(183)=>zero_11, BIAS(182)=>zero_11, BIAS(181)
      =>zero_11, BIAS(180)=>zero_11, BIAS(179)=>zero_11, BIAS(178)=>zero_11, 
      BIAS(177)=>zero_11, BIAS(176)=>zero_11, BIAS(175)=>zero_11, BIAS(174)
      =>zero_11, BIAS(173)=>zero_11, BIAS(172)=>zero_11, BIAS(171)=>zero_11, 
      BIAS(170)=>zero_11, BIAS(169)=>zero_11, BIAS(168)=>zero_11, BIAS(167)
      =>zero_11, BIAS(166)=>zero_11, BIAS(165)=>zero_11, BIAS(164)=>zero_11, 
      BIAS(163)=>zero_11, BIAS(162)=>zero_11, BIAS(161)=>zero_11, BIAS(160)
      =>zero_11, BIAS(159)=>zero_11, BIAS(158)=>zero_11, BIAS(157)=>zero_11, 
      BIAS(156)=>zero_11, BIAS(155)=>zero_11, BIAS(154)=>zero_11, BIAS(153)
      =>zero_11, BIAS(152)=>zero_11, BIAS(151)=>zero_11, BIAS(150)=>zero_11, 
      BIAS(149)=>zero_11, BIAS(148)=>zero_11, BIAS(147)=>zero_11, BIAS(146)
      =>zero_11, BIAS(145)=>zero_11, BIAS(144)=>zero_11, BIAS(143)=>zero_11, 
      BIAS(142)=>zero_11, BIAS(141)=>zero_11, BIAS(140)=>zero_11, BIAS(139)
      =>zero_11, BIAS(138)=>zero_11, BIAS(137)=>zero_11, BIAS(136)=>zero_11, 
      BIAS(135)=>zero_11, BIAS(134)=>zero_11, BIAS(133)=>zero_11, BIAS(132)
      =>zero_11, BIAS(131)=>zero_11, BIAS(130)=>zero_11, BIAS(129)=>zero_11, 
      BIAS(128)=>zero_11, BIAS(127)=>nx10032, BIAS(126)=>nx10034, BIAS(125)
      =>nx10036, BIAS(124)=>nx10038, BIAS(123)=>nx10040, BIAS(122)=>nx10042, 
      BIAS(121)=>nx10044, BIAS(120)=>nx10046, BIAS(119)=>nx10048, BIAS(118)
      =>nx10050, BIAS(117)=>nx10052, BIAS(116)=>nx10054, BIAS(115)=>nx10056, 
      BIAS(114)=>nx10058, BIAS(113)=>nx10060, BIAS(112)=>nx10062, BIAS(111)
      =>nx10064, BIAS(110)=>nx10066, BIAS(109)=>nx10068, BIAS(108)=>nx10070, 
      BIAS(107)=>nx10072, BIAS(106)=>nx10074, BIAS(105)=>nx10076, BIAS(104)
      =>nx10078, BIAS(103)=>nx10080, BIAS(102)=>nx10082, BIAS(101)=>nx10084, 
      BIAS(100)=>nx10086, BIAS(99)=>nx10088, BIAS(98)=>nx10090, BIAS(97)=>
      nx10092, BIAS(96)=>nx10094, BIAS(95)=>nx10096, BIAS(94)=>nx10098, 
      BIAS(93)=>nx10100, BIAS(92)=>nx10102, BIAS(91)=>nx10104, BIAS(90)=>
      nx10106, BIAS(89)=>nx10108, BIAS(88)=>nx10110, BIAS(87)=>nx10112, 
      BIAS(86)=>nx10114, BIAS(85)=>nx10116, BIAS(84)=>nx10118, BIAS(83)=>
      nx10120, BIAS(82)=>nx10122, BIAS(81)=>nx10124, BIAS(80)=>nx10126, 
      BIAS(79)=>nx10128, BIAS(78)=>nx10130, BIAS(77)=>nx10132, BIAS(76)=>
      nx10134, BIAS(75)=>nx10136, BIAS(74)=>nx10138, BIAS(73)=>nx10140, 
      BIAS(72)=>nx10142, BIAS(71)=>nx10144, BIAS(70)=>nx10146, BIAS(69)=>
      nx10148, BIAS(68)=>nx10150, BIAS(67)=>nx10152, BIAS(66)=>nx10154, 
      BIAS(65)=>nx10156, BIAS(64)=>nx10158, BIAS(63)=>nx10160, BIAS(62)=>
      nx10162, BIAS(61)=>nx10164, BIAS(60)=>nx10166, BIAS(59)=>nx10168, 
      BIAS(58)=>nx10170, BIAS(57)=>nx10172, BIAS(56)=>nx10174, BIAS(55)=>
      nx10176, BIAS(54)=>nx10178, BIAS(53)=>nx10180, BIAS(52)=>nx10182, 
      BIAS(51)=>nx10184, BIAS(50)=>nx10186, BIAS(49)=>nx10188, BIAS(48)=>
      nx10190, BIAS(47)=>nx10192, BIAS(46)=>nx10194, BIAS(45)=>nx10196, 
      BIAS(44)=>nx10198, BIAS(43)=>nx10200, BIAS(42)=>nx10202, BIAS(41)=>
      nx10204, BIAS(40)=>nx10206, BIAS(39)=>nx10208, BIAS(38)=>nx10210, 
      BIAS(37)=>nx10212, BIAS(36)=>nx10214, BIAS(35)=>nx10216, BIAS(34)=>
      nx10218, BIAS(33)=>nx10220, BIAS(32)=>nx10222, BIAS(31)=>nx10224, 
      BIAS(30)=>nx10226, BIAS(29)=>nx10228, BIAS(28)=>nx10230, BIAS(27)=>
      nx10232, BIAS(26)=>nx10234, BIAS(25)=>nx10236, BIAS(24)=>nx10238, 
      BIAS(23)=>nx10240, BIAS(22)=>nx10242, BIAS(21)=>nx10244, BIAS(20)=>
      nx10246, BIAS(19)=>nx10248, BIAS(18)=>nx10250, BIAS(17)=>nx10252, 
      BIAS(16)=>nx10254, BIAS(15)=>nx10260, BIAS(14)=>nx10266, BIAS(13)=>
      nx10272, BIAS(12)=>nx10278, BIAS(11)=>nx10284, BIAS(10)=>nx10290, 
      BIAS(9)=>nx10292, BIAS(8)=>nx10294, BIAS(7)=>nx10294, BIAS(6)=>nx10296, 
      BIAS(5)=>nx10298, BIAS(4)=>nx10298, BIAS(3)=>nx10300, BIAS(2)=>nx10302, 
      BIAS(1)=>nx10304, BIAS(0)=>nx10304, FilterAddress(12)=>nx9976, 
      FilterAddress(11)=>nx9980, FilterAddress(10)=>nx9984, FilterAddress(9)
      =>nx9988, FilterAddress(8)=>nx9992, FilterAddress(7)=>nx9996, 
      FilterAddress(6)=>nx10000, FilterAddress(5)=>nx10004, FilterAddress(4)
      =>nx10008, FilterAddress(3)=>nx10012, FilterAddress(2)=>nx10016, 
      FilterAddress(1)=>nx10020, FilterAddress(0)=>nx10024, 
      DMAAddressToFilter(12)=>AddressF_12, DMAAddressToFilter(11)=>
      AddressF_11, DMAAddressToFilter(10)=>AddressF_10, 
      DMAAddressToFilter(9)=>AddressF_9, DMAAddressToFilter(8)=>AddressF_8, 
      DMAAddressToFilter(7)=>AddressF_7, DMAAddressToFilter(6)=>AddressF_6, 
      DMAAddressToFilter(5)=>AddressF_5, DMAAddressToFilter(4)=>AddressF_4, 
      DMAAddressToFilter(3)=>AddressF_3, DMAAddressToFilter(2)=>AddressF_2, 
      DMAAddressToFilter(1)=>AddressF_1, DMAAddressToFilter(0)=>AddressF_0, 
      UpdatedAddress(12)=>FilterAddressIN_12, UpdatedAddress(11)=>
      FilterAddressIN_11, UpdatedAddress(10)=>FilterAddressIN_10, 
      UpdatedAddress(9)=>FilterAddressIN_9, UpdatedAddress(8)=>
      FilterAddressIN_8, UpdatedAddress(7)=>FilterAddressIN_7, 
      UpdatedAddress(6)=>FilterAddressIN_6, UpdatedAddress(5)=>
      FilterAddressIN_5, UpdatedAddress(4)=>FilterAddressIN_4, 
      UpdatedAddress(3)=>FilterAddressIN_3, UpdatedAddress(2)=>
      FilterAddressIN_2, UpdatedAddress(1)=>FilterAddressIN_1, 
      UpdatedAddress(0)=>FilterAddressIN_0, changerAdd(12)=>
      AddressChangerIN_12, changerAdd(11)=>AddressChangerIN_11, 
      changerAdd(10)=>AddressChangerIN_10, changerAdd(9)=>AddressChangerIN_9, 
      changerAdd(8)=>AddressChangerIN_8, changerAdd(7)=>AddressChangerIN_7, 
      changerAdd(6)=>AddressChangerIN_6, changerAdd(5)=>AddressChangerIN_5, 
      changerAdd(4)=>AddressChangerIN_4, changerAdd(3)=>AddressChangerIN_3, 
      changerAdd(2)=>AddressChangerIN_2, changerAdd(1)=>AddressChangerIN_1, 
      changerAdd(0)=>AddressChangerIN_0, CLK=>nx10416, RST=>rst, 
      LayerInfo(15)=>zero_11, LayerInfo(14)=>zero_11, LayerInfo(13)=>zero_11, 
      LayerInfo(12)=>zero_11, LayerInfo(11)=>zero_11, LayerInfo(10)=>zero_11, 
      LayerInfo(9)=>zero_11, LayerInfo(8)=>zero_11, LayerInfo(7)=>zero_11, 
      LayerInfo(6)=>zero_11, LayerInfo(5)=>zero_11, LayerInfo(4)=>zero_11, 
      LayerInfo(3)=>LayerInfoOut_3, LayerInfo(2)=>LayerInfoOut_2, 
      LayerInfo(1)=>LayerInfoOut_1, LayerInfo(0)=>LayerInfoOut_0, 
      outBias0(15)=>Bias0_15, outBias0(14)=>Bias0_14, outBias0(13)=>Bias0_13, 
      outBias0(12)=>Bias0_12, outBias0(11)=>Bias0_11, outBias0(10)=>Bias0_10, 
      outBias0(9)=>Bias0_9, outBias0(8)=>Bias0_8, outBias0(7)=>Bias0_7, 
      outBias0(6)=>Bias0_6, outBias0(5)=>Bias0_5, outBias0(4)=>Bias0_4, 
      outBias0(3)=>Bias0_3, outBias0(2)=>Bias0_2, outBias0(1)=>Bias0_1, 
      outBias0(0)=>Bias0_0, outBias1(15)=>Bias1_15, outBias1(14)=>Bias1_14, 
      outBias1(13)=>Bias1_13, outBias1(12)=>Bias1_12, outBias1(11)=>Bias1_11, 
      outBias1(10)=>Bias1_10, outBias1(9)=>Bias1_9, outBias1(8)=>Bias1_8, 
      outBias1(7)=>Bias1_7, outBias1(6)=>Bias1_6, outBias1(5)=>Bias1_5, 
      outBias1(4)=>Bias1_4, outBias1(3)=>Bias1_3, outBias1(2)=>Bias1_2, 
      outBias1(1)=>Bias1_1, outBias1(0)=>Bias1_0, outBias2(15)=>Bias2_15, 
      outBias2(14)=>Bias2_14, outBias2(13)=>Bias2_13, outBias2(12)=>Bias2_12, 
      outBias2(11)=>Bias2_11, outBias2(10)=>Bias2_10, outBias2(9)=>Bias2_9, 
      outBias2(8)=>Bias2_8, outBias2(7)=>Bias2_7, outBias2(6)=>Bias2_6, 
      outBias2(5)=>Bias2_5, outBias2(4)=>Bias2_4, outBias2(3)=>Bias2_3, 
      outBias2(2)=>Bias2_2, outBias2(1)=>Bias2_1, outBias2(0)=>Bias2_0, 
      outBias3(15)=>Bias3_15, outBias3(14)=>Bias3_14, outBias3(13)=>Bias3_13, 
      outBias3(12)=>Bias3_12, outBias3(11)=>Bias3_11, outBias3(10)=>Bias3_10, 
      outBias3(9)=>Bias3_9, outBias3(8)=>Bias3_8, outBias3(7)=>Bias3_7, 
      outBias3(6)=>Bias3_6, outBias3(5)=>Bias3_5, outBias3(4)=>Bias3_4, 
      outBias3(3)=>Bias3_3, outBias3(2)=>Bias3_2, outBias3(1)=>Bias3_1, 
      outBias3(0)=>Bias3_0, outBias4(15)=>Bias4_15, outBias4(14)=>Bias4_14, 
      outBias4(13)=>Bias4_13, outBias4(12)=>Bias4_12, outBias4(11)=>Bias4_11, 
      outBias4(10)=>Bias4_10, outBias4(9)=>Bias4_9, outBias4(8)=>Bias4_8, 
      outBias4(7)=>Bias4_7, outBias4(6)=>Bias4_6, outBias4(5)=>Bias4_5, 
      outBias4(4)=>Bias4_4, outBias4(3)=>Bias4_3, outBias4(2)=>Bias4_2, 
      outBias4(1)=>Bias4_1, outBias4(0)=>Bias4_0, outBias5(15)=>Bias5_15, 
      outBias5(14)=>Bias5_14, outBias5(13)=>Bias5_13, outBias5(12)=>Bias5_12, 
      outBias5(11)=>Bias5_11, outBias5(10)=>Bias5_10, outBias5(9)=>Bias5_9, 
      outBias5(8)=>Bias5_8, outBias5(7)=>Bias5_7, outBias5(6)=>Bias5_6, 
      outBias5(5)=>Bias5_5, outBias5(4)=>Bias5_4, outBias5(3)=>Bias5_3, 
      outBias5(2)=>Bias5_2, outBias5(1)=>Bias5_1, outBias5(0)=>Bias5_0, 
      outBias6(15)=>Bias6_15, outBias6(14)=>Bias6_14, outBias6(13)=>Bias6_13, 
      outBias6(12)=>Bias6_12, outBias6(11)=>Bias6_11, outBias6(10)=>Bias6_10, 
      outBias6(9)=>Bias6_9, outBias6(8)=>Bias6_8, outBias6(7)=>Bias6_7, 
      outBias6(6)=>Bias6_6, outBias6(5)=>Bias6_5, outBias6(4)=>Bias6_4, 
      outBias6(3)=>Bias6_3, outBias6(2)=>Bias6_2, outBias6(1)=>Bias6_1, 
      outBias6(0)=>Bias6_0, outBias7(15)=>Bias7_15, outBias7(14)=>Bias7_14, 
      outBias7(13)=>Bias7_13, outBias7(12)=>Bias7_12, outBias7(11)=>Bias7_11, 
      outBias7(10)=>Bias7_10, outBias7(9)=>Bias7_9, outBias7(8)=>Bias7_8, 
      outBias7(7)=>Bias7_7, outBias7(6)=>Bias7_6, outBias7(5)=>Bias7_5, 
      outBias7(4)=>Bias7_4, outBias7(3)=>Bias7_3, outBias7(2)=>Bias7_2, 
      outBias7(1)=>Bias7_1, outBias7(0)=>Bias7_0, ACKF=>nx10308);
   Rfilter : ReadFilter port map ( current_state(14)=>zero_11, 
      current_state(13)=>zero_11, current_state(12)=>zero_11, 
      current_state(11)=>zero_11, current_state(10)=>current_state_10, 
      current_state(9)=>zero_11, current_state(8)=>zero_11, current_state(7)
      =>nx9962, current_state(6)=>zero_11, current_state(5)=>current_state_5, 
      current_state(4)=>zero_11, current_state(3)=>zero_11, current_state(2)
      =>zero_11, current_state(1)=>zero_11, current_state(0)=>zero_11, 
      LayerInfo(15)=>zero_11, LayerInfo(14)=>zero_11, LayerInfo(13)=>zero_11, 
      LayerInfo(12)=>LayerInfoOut_12, LayerInfo(11)=>LayerInfoOut_11, 
      LayerInfo(10)=>LayerInfoOut_10, LayerInfo(9)=>LayerInfoOut_9, 
      LayerInfo(8)=>nx10378, LayerInfo(7)=>nx10382, LayerInfo(6)=>nx10386, 
      LayerInfo(5)=>nx10388, LayerInfo(4)=>nx10392, LayerInfo(3)=>
      LayerInfoOut_3, LayerInfo(2)=>LayerInfoOut_2, LayerInfo(1)=>
      LayerInfoOut_1, LayerInfo(0)=>LayerInfoOut_0, depthcounter(3)=>nx10406, 
      depthcounter(2)=>nx10408, depthcounter(1)=>nx10410, depthcounter(0)=>
      nx10412, FilterCounter(3)=>nx10398, FilterCounter(2)=>nx10400, 
      FilterCounter(1)=>nx10402, FilterCounter(0)=>nx10404, Heightcounter(4)
      =>NumOfHeight_4, Heightcounter(3)=>NumOfHeight_3, Heightcounter(2)=>
      NumOfHeight_2, Heightcounter(1)=>NumOfHeight_1, Heightcounter(0)=>
      NumOfHeight_0, FILTER(399)=>nx10032, FILTER(398)=>nx10032, FILTER(397)
      =>nx10032, FILTER(396)=>nx10034, FILTER(395)=>nx10034, FILTER(394)=>
      nx10034, FILTER(393)=>nx10036, FILTER(392)=>nx10036, FILTER(391)=>
      nx10036, FILTER(390)=>nx10038, FILTER(389)=>nx10038, FILTER(388)=>
      nx10038, FILTER(387)=>nx10040, FILTER(386)=>nx10040, FILTER(385)=>
      nx10040, FILTER(384)=>nx10042, FILTER(383)=>nx10042, FILTER(382)=>
      nx10042, FILTER(381)=>nx10044, FILTER(380)=>nx10044, FILTER(379)=>
      nx10044, FILTER(378)=>nx10046, FILTER(377)=>nx10046, FILTER(376)=>
      nx10046, FILTER(375)=>nx10048, FILTER(374)=>nx10048, FILTER(373)=>
      nx10048, FILTER(372)=>nx10050, FILTER(371)=>nx10050, FILTER(370)=>
      nx10050, FILTER(369)=>nx10052, FILTER(368)=>nx10052, FILTER(367)=>
      nx10052, FILTER(366)=>nx10054, FILTER(365)=>nx10054, FILTER(364)=>
      nx10054, FILTER(363)=>nx10056, FILTER(362)=>nx10056, FILTER(361)=>
      nx10056, FILTER(360)=>nx10058, FILTER(359)=>nx10058, FILTER(358)=>
      nx10058, FILTER(357)=>nx10060, FILTER(356)=>nx10060, FILTER(355)=>
      nx10060, FILTER(354)=>nx10062, FILTER(353)=>nx10062, FILTER(352)=>
      nx10062, FILTER(351)=>nx10064, FILTER(350)=>nx10064, FILTER(349)=>
      nx10064, FILTER(348)=>nx10066, FILTER(347)=>nx10066, FILTER(346)=>
      nx10066, FILTER(345)=>nx10068, FILTER(344)=>nx10068, FILTER(343)=>
      nx10068, FILTER(342)=>nx10070, FILTER(341)=>nx10070, FILTER(340)=>
      nx10070, FILTER(339)=>nx10072, FILTER(338)=>nx10072, FILTER(337)=>
      nx10072, FILTER(336)=>nx10074, FILTER(335)=>nx10074, FILTER(334)=>
      nx10074, FILTER(333)=>nx10076, FILTER(332)=>nx10076, FILTER(331)=>
      nx10076, FILTER(330)=>nx10078, FILTER(329)=>nx10078, FILTER(328)=>
      nx10078, FILTER(327)=>nx10080, FILTER(326)=>nx10080, FILTER(325)=>
      nx10080, FILTER(324)=>nx10082, FILTER(323)=>nx10082, FILTER(322)=>
      nx10082, FILTER(321)=>nx10084, FILTER(320)=>nx10084, FILTER(319)=>
      nx10084, FILTER(318)=>nx10086, FILTER(317)=>nx10086, FILTER(316)=>
      nx10086, FILTER(315)=>nx10088, FILTER(314)=>nx10088, FILTER(313)=>
      nx10088, FILTER(312)=>nx10090, FILTER(311)=>nx10090, FILTER(310)=>
      nx10090, FILTER(309)=>nx10092, FILTER(308)=>nx10092, FILTER(307)=>
      nx10092, FILTER(306)=>nx10094, FILTER(305)=>nx10094, FILTER(304)=>
      nx10094, FILTER(303)=>nx10096, FILTER(302)=>nx10096, FILTER(301)=>
      nx10096, FILTER(300)=>nx10098, FILTER(299)=>nx10098, FILTER(298)=>
      nx10098, FILTER(297)=>nx10100, FILTER(296)=>nx10100, FILTER(295)=>
      nx10100, FILTER(294)=>nx10102, FILTER(293)=>nx10102, FILTER(292)=>
      nx10102, FILTER(291)=>nx10104, FILTER(290)=>nx10104, FILTER(289)=>
      nx10104, FILTER(288)=>nx10106, FILTER(287)=>nx10106, FILTER(286)=>
      nx10106, FILTER(285)=>nx10108, FILTER(284)=>nx10108, FILTER(283)=>
      nx10108, FILTER(282)=>nx10110, FILTER(281)=>nx10110, FILTER(280)=>
      nx10110, FILTER(279)=>nx10112, FILTER(278)=>nx10112, FILTER(277)=>
      nx10112, FILTER(276)=>nx10114, FILTER(275)=>nx10114, FILTER(274)=>
      nx10114, FILTER(273)=>nx10116, FILTER(272)=>nx10116, FILTER(271)=>
      nx10116, FILTER(270)=>nx10118, FILTER(269)=>nx10118, FILTER(268)=>
      nx10118, FILTER(267)=>nx10120, FILTER(266)=>nx10120, FILTER(265)=>
      nx10120, FILTER(264)=>nx10122, FILTER(263)=>nx10122, FILTER(262)=>
      nx10122, FILTER(261)=>nx10124, FILTER(260)=>nx10124, FILTER(259)=>
      nx10124, FILTER(258)=>nx10126, FILTER(257)=>nx10126, FILTER(256)=>
      nx10126, FILTER(255)=>nx10128, FILTER(254)=>nx10128, FILTER(253)=>
      nx10128, FILTER(252)=>nx10130, FILTER(251)=>nx10130, FILTER(250)=>
      nx10130, FILTER(249)=>nx10132, FILTER(248)=>nx10132, FILTER(247)=>
      nx10132, FILTER(246)=>nx10134, FILTER(245)=>nx10134, FILTER(244)=>
      nx10134, FILTER(243)=>nx10136, FILTER(242)=>nx10136, FILTER(241)=>
      nx10136, FILTER(240)=>nx10138, FILTER(239)=>nx10138, FILTER(238)=>
      nx10138, FILTER(237)=>nx10140, FILTER(236)=>nx10140, FILTER(235)=>
      nx10140, FILTER(234)=>nx10142, FILTER(233)=>nx10142, FILTER(232)=>
      nx10142, FILTER(231)=>nx10144, FILTER(230)=>nx10144, FILTER(229)=>
      nx10144, FILTER(228)=>nx10146, FILTER(227)=>nx10146, FILTER(226)=>
      nx10146, FILTER(225)=>nx10148, FILTER(224)=>nx10148, FILTER(223)=>
      nx10148, FILTER(222)=>nx10150, FILTER(221)=>nx10150, FILTER(220)=>
      nx10150, FILTER(219)=>nx10152, FILTER(218)=>nx10152, FILTER(217)=>
      nx10152, FILTER(216)=>nx10154, FILTER(215)=>nx10154, FILTER(214)=>
      nx10154, FILTER(213)=>nx10156, FILTER(212)=>nx10156, FILTER(211)=>
      nx10156, FILTER(210)=>nx10158, FILTER(209)=>nx10158, FILTER(208)=>
      nx10158, FILTER(207)=>nx10160, FILTER(206)=>nx10160, FILTER(205)=>
      nx10160, FILTER(204)=>nx10162, FILTER(203)=>nx10162, FILTER(202)=>
      nx10162, FILTER(201)=>nx10164, FILTER(200)=>nx10164, FILTER(199)=>
      nx10164, FILTER(198)=>nx10166, FILTER(197)=>nx10166, FILTER(196)=>
      nx10166, FILTER(195)=>nx10168, FILTER(194)=>nx10168, FILTER(193)=>
      nx10168, FILTER(192)=>nx10170, FILTER(191)=>nx10170, FILTER(190)=>
      nx10170, FILTER(189)=>nx10172, FILTER(188)=>nx10172, FILTER(187)=>
      nx10172, FILTER(186)=>nx10174, FILTER(185)=>nx10174, FILTER(184)=>
      nx10174, FILTER(183)=>nx10176, FILTER(182)=>nx10176, FILTER(181)=>
      nx10176, FILTER(180)=>nx10178, FILTER(179)=>nx10178, FILTER(178)=>
      nx10178, FILTER(177)=>nx10180, FILTER(176)=>nx10180, FILTER(175)=>
      nx10180, FILTER(174)=>nx10182, FILTER(173)=>nx10182, FILTER(172)=>
      nx10182, FILTER(171)=>nx10184, FILTER(170)=>nx10184, FILTER(169)=>
      nx10184, FILTER(168)=>nx10186, FILTER(167)=>nx10186, FILTER(166)=>
      nx10186, FILTER(165)=>nx10188, FILTER(164)=>nx10188, FILTER(163)=>
      nx10188, FILTER(162)=>nx10190, FILTER(161)=>nx10190, FILTER(160)=>
      nx10190, FILTER(159)=>nx10192, FILTER(158)=>nx10192, FILTER(157)=>
      nx10192, FILTER(156)=>nx10194, FILTER(155)=>nx10194, FILTER(154)=>
      nx10194, FILTER(153)=>nx10196, FILTER(152)=>nx10196, FILTER(151)=>
      nx10196, FILTER(150)=>nx10198, FILTER(149)=>nx10198, FILTER(148)=>
      nx10198, FILTER(147)=>nx10200, FILTER(146)=>nx10200, FILTER(145)=>
      nx10200, FILTER(144)=>nx10202, FILTER(143)=>nx10202, FILTER(142)=>
      nx10202, FILTER(141)=>nx10204, FILTER(140)=>nx10204, FILTER(139)=>
      nx10204, FILTER(138)=>nx10206, FILTER(137)=>nx10206, FILTER(136)=>
      nx10206, FILTER(135)=>nx10208, FILTER(134)=>nx10208, FILTER(133)=>
      nx10208, FILTER(132)=>nx10210, FILTER(131)=>nx10210, FILTER(130)=>
      nx10210, FILTER(129)=>nx10212, FILTER(128)=>nx10212, FILTER(127)=>
      nx10212, FILTER(126)=>nx10214, FILTER(125)=>nx10214, FILTER(124)=>
      nx10214, FILTER(123)=>nx10216, FILTER(122)=>nx10216, FILTER(121)=>
      nx10216, FILTER(120)=>nx10218, FILTER(119)=>nx10218, FILTER(118)=>
      nx10218, FILTER(117)=>nx10220, FILTER(116)=>nx10220, FILTER(115)=>
      nx10220, FILTER(114)=>nx10222, FILTER(113)=>nx10222, FILTER(112)=>
      nx10222, FILTER(111)=>nx10224, FILTER(110)=>nx10224, FILTER(109)=>
      nx10224, FILTER(108)=>nx10226, FILTER(107)=>nx10226, FILTER(106)=>
      nx10226, FILTER(105)=>nx10228, FILTER(104)=>nx10228, FILTER(103)=>
      nx10228, FILTER(102)=>nx10230, FILTER(101)=>nx10230, FILTER(100)=>
      nx10230, FILTER(99)=>nx10232, FILTER(98)=>nx10232, FILTER(97)=>nx10232, 
      FILTER(96)=>nx10234, FILTER(95)=>nx10234, FILTER(94)=>nx10234, 
      FILTER(93)=>nx10236, FILTER(92)=>nx10236, FILTER(91)=>nx10236, 
      FILTER(90)=>nx10238, FILTER(89)=>nx10238, FILTER(88)=>nx10238, 
      FILTER(87)=>nx10240, FILTER(86)=>nx10240, FILTER(85)=>nx10240, 
      FILTER(84)=>nx10242, FILTER(83)=>nx10242, FILTER(82)=>nx10242, 
      FILTER(81)=>nx10244, FILTER(80)=>nx10244, FILTER(79)=>nx10244, 
      FILTER(78)=>nx10246, FILTER(77)=>nx10246, FILTER(76)=>nx10246, 
      FILTER(75)=>nx10248, FILTER(74)=>nx10248, FILTER(73)=>nx10248, 
      FILTER(72)=>nx10250, FILTER(71)=>nx10250, FILTER(70)=>nx10250, 
      FILTER(69)=>nx10252, FILTER(68)=>nx10252, FILTER(67)=>nx10252, 
      FILTER(66)=>nx10254, FILTER(65)=>nx10254, FILTER(64)=>nx10254, 
      FILTER(63)=>nx10256, FILTER(62)=>nx10256, FILTER(61)=>nx10256, 
      FILTER(60)=>nx10258, FILTER(59)=>nx10258, FILTER(58)=>nx10258, 
      FILTER(57)=>nx10260, FILTER(56)=>nx10260, FILTER(55)=>nx10260, 
      FILTER(54)=>nx10262, FILTER(53)=>nx10262, FILTER(52)=>nx10262, 
      FILTER(51)=>nx10264, FILTER(50)=>nx10264, FILTER(49)=>nx10264, 
      FILTER(48)=>nx10266, FILTER(47)=>nx10266, FILTER(46)=>nx10266, 
      FILTER(45)=>nx10268, FILTER(44)=>nx10268, FILTER(43)=>nx10268, 
      FILTER(42)=>nx10270, FILTER(41)=>nx10270, FILTER(40)=>nx10270, 
      FILTER(39)=>nx10272, FILTER(38)=>nx10272, FILTER(37)=>nx10272, 
      FILTER(36)=>nx10274, FILTER(35)=>nx10274, FILTER(34)=>nx10274, 
      FILTER(33)=>nx10276, FILTER(32)=>nx10276, FILTER(31)=>nx10276, 
      FILTER(30)=>nx10278, FILTER(29)=>nx10278, FILTER(28)=>nx10278, 
      FILTER(27)=>nx10280, FILTER(26)=>nx10280, FILTER(25)=>nx10280, 
      FILTER(24)=>nx10282, FILTER(23)=>nx10282, FILTER(22)=>nx10282, 
      FILTER(21)=>nx10284, FILTER(20)=>nx10284, FILTER(19)=>nx10284, 
      FILTER(18)=>nx10286, FILTER(17)=>nx10286, FILTER(16)=>nx10286, 
      FILTER(15)=>nx10288, FILTER(14)=>nx10288, FILTER(13)=>nx10288, 
      FILTER(12)=>nx10290, FILTER(11)=>nx10290, FILTER(10)=>nx10290, 
      FILTER(9)=>nx10292, FILTER(8)=>nx10294, FILTER(7)=>nx10296, FILTER(6)
      =>nx10296, FILTER(5)=>nx10298, FILTER(4)=>nx10300, FILTER(3)=>nx10300, 
      FILTER(2)=>nx10302, FILTER(1)=>nx10304, FILTER(0)=>nx10306, 
      FilterAddress(12)=>nx9976, FilterAddress(11)=>nx9980, 
      FilterAddress(10)=>nx9984, FilterAddress(9)=>nx9988, FilterAddress(8)
      =>nx9992, FilterAddress(7)=>nx9996, FilterAddress(6)=>nx10000, 
      FilterAddress(5)=>nx10004, FilterAddress(4)=>nx10008, FilterAddress(3)
      =>nx10012, FilterAddress(2)=>nx10016, FilterAddress(1)=>nx10020, 
      FilterAddress(0)=>nx10024, msbNoOfFilters=>nx10500, CLK=>nx10422, RST
      =>rst, QImgStat=>Q, ACKF=>nx10308, IndicatorFilter(0)=>IndicatorF_0, 
      DMAAddress(12)=>AddressF_12, DMAAddress(11)=>AddressF_11, 
      DMAAddress(10)=>AddressF_10, DMAAddress(9)=>AddressF_9, DMAAddress(8)
      =>AddressF_8, DMAAddress(7)=>AddressF_7, DMAAddress(6)=>AddressF_6, 
      DMAAddress(5)=>AddressF_5, DMAAddress(4)=>AddressF_4, DMAAddress(3)=>
      AddressF_3, DMAAddress(2)=>AddressF_2, DMAAddress(1)=>AddressF_1, 
      DMAAddress(0)=>AddressF_0, UpdatedAddress(12)=>FilterAddressIN_12, 
      UpdatedAddress(11)=>FilterAddressIN_11, UpdatedAddress(10)=>
      FilterAddressIN_10, UpdatedAddress(9)=>FilterAddressIN_9, 
      UpdatedAddress(8)=>FilterAddressIN_8, UpdatedAddress(7)=>
      FilterAddressIN_7, UpdatedAddress(6)=>FilterAddressIN_6, 
      UpdatedAddress(5)=>FilterAddressIN_5, UpdatedAddress(4)=>
      FilterAddressIN_4, UpdatedAddress(3)=>FilterAddressIN_3, 
      UpdatedAddress(2)=>FilterAddressIN_2, UpdatedAddress(1)=>
      FilterAddressIN_1, UpdatedAddress(0)=>FilterAddressIN_0, 
      outFilter0(399)=>Filter1_399, outFilter0(398)=>Filter1_398, 
      outFilter0(397)=>Filter1_397, outFilter0(396)=>Filter1_396, 
      outFilter0(395)=>Filter1_395, outFilter0(394)=>Filter1_394, 
      outFilter0(393)=>Filter1_393, outFilter0(392)=>Filter1_392, 
      outFilter0(391)=>Filter1_391, outFilter0(390)=>Filter1_390, 
      outFilter0(389)=>Filter1_389, outFilter0(388)=>Filter1_388, 
      outFilter0(387)=>Filter1_387, outFilter0(386)=>Filter1_386, 
      outFilter0(385)=>Filter1_385, outFilter0(384)=>Filter1_384, 
      outFilter0(383)=>Filter1_383, outFilter0(382)=>Filter1_382, 
      outFilter0(381)=>Filter1_381, outFilter0(380)=>Filter1_380, 
      outFilter0(379)=>Filter1_379, outFilter0(378)=>Filter1_378, 
      outFilter0(377)=>Filter1_377, outFilter0(376)=>Filter1_376, 
      outFilter0(375)=>Filter1_375, outFilter0(374)=>Filter1_374, 
      outFilter0(373)=>Filter1_373, outFilter0(372)=>Filter1_372, 
      outFilter0(371)=>Filter1_371, outFilter0(370)=>Filter1_370, 
      outFilter0(369)=>Filter1_369, outFilter0(368)=>Filter1_368, 
      outFilter0(367)=>Filter1_367, outFilter0(366)=>Filter1_366, 
      outFilter0(365)=>Filter1_365, outFilter0(364)=>Filter1_364, 
      outFilter0(363)=>Filter1_363, outFilter0(362)=>Filter1_362, 
      outFilter0(361)=>Filter1_361, outFilter0(360)=>Filter1_360, 
      outFilter0(359)=>Filter1_359, outFilter0(358)=>Filter1_358, 
      outFilter0(357)=>Filter1_357, outFilter0(356)=>Filter1_356, 
      outFilter0(355)=>Filter1_355, outFilter0(354)=>Filter1_354, 
      outFilter0(353)=>Filter1_353, outFilter0(352)=>Filter1_352, 
      outFilter0(351)=>Filter1_351, outFilter0(350)=>Filter1_350, 
      outFilter0(349)=>Filter1_349, outFilter0(348)=>Filter1_348, 
      outFilter0(347)=>Filter1_347, outFilter0(346)=>Filter1_346, 
      outFilter0(345)=>Filter1_345, outFilter0(344)=>Filter1_344, 
      outFilter0(343)=>Filter1_343, outFilter0(342)=>Filter1_342, 
      outFilter0(341)=>Filter1_341, outFilter0(340)=>Filter1_340, 
      outFilter0(339)=>Filter1_339, outFilter0(338)=>Filter1_338, 
      outFilter0(337)=>Filter1_337, outFilter0(336)=>Filter1_336, 
      outFilter0(335)=>Filter1_335, outFilter0(334)=>Filter1_334, 
      outFilter0(333)=>Filter1_333, outFilter0(332)=>Filter1_332, 
      outFilter0(331)=>Filter1_331, outFilter0(330)=>Filter1_330, 
      outFilter0(329)=>Filter1_329, outFilter0(328)=>Filter1_328, 
      outFilter0(327)=>Filter1_327, outFilter0(326)=>Filter1_326, 
      outFilter0(325)=>Filter1_325, outFilter0(324)=>Filter1_324, 
      outFilter0(323)=>Filter1_323, outFilter0(322)=>Filter1_322, 
      outFilter0(321)=>Filter1_321, outFilter0(320)=>Filter1_320, 
      outFilter0(319)=>Filter1_319, outFilter0(318)=>Filter1_318, 
      outFilter0(317)=>Filter1_317, outFilter0(316)=>Filter1_316, 
      outFilter0(315)=>Filter1_315, outFilter0(314)=>Filter1_314, 
      outFilter0(313)=>Filter1_313, outFilter0(312)=>Filter1_312, 
      outFilter0(311)=>Filter1_311, outFilter0(310)=>Filter1_310, 
      outFilter0(309)=>Filter1_309, outFilter0(308)=>Filter1_308, 
      outFilter0(307)=>Filter1_307, outFilter0(306)=>Filter1_306, 
      outFilter0(305)=>Filter1_305, outFilter0(304)=>Filter1_304, 
      outFilter0(303)=>Filter1_303, outFilter0(302)=>Filter1_302, 
      outFilter0(301)=>Filter1_301, outFilter0(300)=>Filter1_300, 
      outFilter0(299)=>Filter1_299, outFilter0(298)=>Filter1_298, 
      outFilter0(297)=>Filter1_297, outFilter0(296)=>Filter1_296, 
      outFilter0(295)=>Filter1_295, outFilter0(294)=>Filter1_294, 
      outFilter0(293)=>Filter1_293, outFilter0(292)=>Filter1_292, 
      outFilter0(291)=>Filter1_291, outFilter0(290)=>Filter1_290, 
      outFilter0(289)=>Filter1_289, outFilter0(288)=>Filter1_288, 
      outFilter0(287)=>Filter1_287, outFilter0(286)=>Filter1_286, 
      outFilter0(285)=>Filter1_285, outFilter0(284)=>Filter1_284, 
      outFilter0(283)=>Filter1_283, outFilter0(282)=>Filter1_282, 
      outFilter0(281)=>Filter1_281, outFilter0(280)=>Filter1_280, 
      outFilter0(279)=>Filter1_279, outFilter0(278)=>Filter1_278, 
      outFilter0(277)=>Filter1_277, outFilter0(276)=>Filter1_276, 
      outFilter0(275)=>Filter1_275, outFilter0(274)=>Filter1_274, 
      outFilter0(273)=>Filter1_273, outFilter0(272)=>Filter1_272, 
      outFilter0(271)=>Filter1_271, outFilter0(270)=>Filter1_270, 
      outFilter0(269)=>Filter1_269, outFilter0(268)=>Filter1_268, 
      outFilter0(267)=>Filter1_267, outFilter0(266)=>Filter1_266, 
      outFilter0(265)=>Filter1_265, outFilter0(264)=>Filter1_264, 
      outFilter0(263)=>Filter1_263, outFilter0(262)=>Filter1_262, 
      outFilter0(261)=>Filter1_261, outFilter0(260)=>Filter1_260, 
      outFilter0(259)=>Filter1_259, outFilter0(258)=>Filter1_258, 
      outFilter0(257)=>Filter1_257, outFilter0(256)=>Filter1_256, 
      outFilter0(255)=>Filter1_255, outFilter0(254)=>Filter1_254, 
      outFilter0(253)=>Filter1_253, outFilter0(252)=>Filter1_252, 
      outFilter0(251)=>Filter1_251, outFilter0(250)=>Filter1_250, 
      outFilter0(249)=>Filter1_249, outFilter0(248)=>Filter1_248, 
      outFilter0(247)=>Filter1_247, outFilter0(246)=>Filter1_246, 
      outFilter0(245)=>Filter1_245, outFilter0(244)=>Filter1_244, 
      outFilter0(243)=>Filter1_243, outFilter0(242)=>Filter1_242, 
      outFilter0(241)=>Filter1_241, outFilter0(240)=>Filter1_240, 
      outFilter0(239)=>Filter1_239, outFilter0(238)=>Filter1_238, 
      outFilter0(237)=>Filter1_237, outFilter0(236)=>Filter1_236, 
      outFilter0(235)=>Filter1_235, outFilter0(234)=>Filter1_234, 
      outFilter0(233)=>Filter1_233, outFilter0(232)=>Filter1_232, 
      outFilter0(231)=>Filter1_231, outFilter0(230)=>Filter1_230, 
      outFilter0(229)=>Filter1_229, outFilter0(228)=>Filter1_228, 
      outFilter0(227)=>Filter1_227, outFilter0(226)=>Filter1_226, 
      outFilter0(225)=>Filter1_225, outFilter0(224)=>Filter1_224, 
      outFilter0(223)=>Filter1_223, outFilter0(222)=>Filter1_222, 
      outFilter0(221)=>Filter1_221, outFilter0(220)=>Filter1_220, 
      outFilter0(219)=>Filter1_219, outFilter0(218)=>Filter1_218, 
      outFilter0(217)=>Filter1_217, outFilter0(216)=>Filter1_216, 
      outFilter0(215)=>Filter1_215, outFilter0(214)=>Filter1_214, 
      outFilter0(213)=>Filter1_213, outFilter0(212)=>Filter1_212, 
      outFilter0(211)=>Filter1_211, outFilter0(210)=>Filter1_210, 
      outFilter0(209)=>Filter1_209, outFilter0(208)=>Filter1_208, 
      outFilter0(207)=>Filter1_207, outFilter0(206)=>Filter1_206, 
      outFilter0(205)=>Filter1_205, outFilter0(204)=>Filter1_204, 
      outFilter0(203)=>Filter1_203, outFilter0(202)=>Filter1_202, 
      outFilter0(201)=>Filter1_201, outFilter0(200)=>Filter1_200, 
      outFilter0(199)=>Filter1_199, outFilter0(198)=>Filter1_198, 
      outFilter0(197)=>Filter1_197, outFilter0(196)=>Filter1_196, 
      outFilter0(195)=>Filter1_195, outFilter0(194)=>Filter1_194, 
      outFilter0(193)=>Filter1_193, outFilter0(192)=>Filter1_192, 
      outFilter0(191)=>Filter1_191, outFilter0(190)=>Filter1_190, 
      outFilter0(189)=>Filter1_189, outFilter0(188)=>Filter1_188, 
      outFilter0(187)=>Filter1_187, outFilter0(186)=>Filter1_186, 
      outFilter0(185)=>Filter1_185, outFilter0(184)=>Filter1_184, 
      outFilter0(183)=>Filter1_183, outFilter0(182)=>Filter1_182, 
      outFilter0(181)=>Filter1_181, outFilter0(180)=>Filter1_180, 
      outFilter0(179)=>Filter1_179, outFilter0(178)=>Filter1_178, 
      outFilter0(177)=>Filter1_177, outFilter0(176)=>Filter1_176, 
      outFilter0(175)=>Filter1_175, outFilter0(174)=>Filter1_174, 
      outFilter0(173)=>Filter1_173, outFilter0(172)=>Filter1_172, 
      outFilter0(171)=>Filter1_171, outFilter0(170)=>Filter1_170, 
      outFilter0(169)=>Filter1_169, outFilter0(168)=>Filter1_168, 
      outFilter0(167)=>Filter1_167, outFilter0(166)=>Filter1_166, 
      outFilter0(165)=>Filter1_165, outFilter0(164)=>Filter1_164, 
      outFilter0(163)=>Filter1_163, outFilter0(162)=>Filter1_162, 
      outFilter0(161)=>Filter1_161, outFilter0(160)=>Filter1_160, 
      outFilter0(159)=>Filter1_159, outFilter0(158)=>Filter1_158, 
      outFilter0(157)=>Filter1_157, outFilter0(156)=>Filter1_156, 
      outFilter0(155)=>Filter1_155, outFilter0(154)=>Filter1_154, 
      outFilter0(153)=>Filter1_153, outFilter0(152)=>Filter1_152, 
      outFilter0(151)=>Filter1_151, outFilter0(150)=>Filter1_150, 
      outFilter0(149)=>Filter1_149, outFilter0(148)=>Filter1_148, 
      outFilter0(147)=>Filter1_147, outFilter0(146)=>Filter1_146, 
      outFilter0(145)=>Filter1_145, outFilter0(144)=>Filter1_144, 
      outFilter0(143)=>Filter1_143, outFilter0(142)=>Filter1_142, 
      outFilter0(141)=>Filter1_141, outFilter0(140)=>Filter1_140, 
      outFilter0(139)=>Filter1_139, outFilter0(138)=>Filter1_138, 
      outFilter0(137)=>Filter1_137, outFilter0(136)=>Filter1_136, 
      outFilter0(135)=>Filter1_135, outFilter0(134)=>Filter1_134, 
      outFilter0(133)=>Filter1_133, outFilter0(132)=>Filter1_132, 
      outFilter0(131)=>Filter1_131, outFilter0(130)=>Filter1_130, 
      outFilter0(129)=>Filter1_129, outFilter0(128)=>Filter1_128, 
      outFilter0(127)=>Filter1_127, outFilter0(126)=>Filter1_126, 
      outFilter0(125)=>Filter1_125, outFilter0(124)=>Filter1_124, 
      outFilter0(123)=>Filter1_123, outFilter0(122)=>Filter1_122, 
      outFilter0(121)=>Filter1_121, outFilter0(120)=>Filter1_120, 
      outFilter0(119)=>Filter1_119, outFilter0(118)=>Filter1_118, 
      outFilter0(117)=>Filter1_117, outFilter0(116)=>Filter1_116, 
      outFilter0(115)=>Filter1_115, outFilter0(114)=>Filter1_114, 
      outFilter0(113)=>Filter1_113, outFilter0(112)=>Filter1_112, 
      outFilter0(111)=>Filter1_111, outFilter0(110)=>Filter1_110, 
      outFilter0(109)=>Filter1_109, outFilter0(108)=>Filter1_108, 
      outFilter0(107)=>Filter1_107, outFilter0(106)=>Filter1_106, 
      outFilter0(105)=>Filter1_105, outFilter0(104)=>Filter1_104, 
      outFilter0(103)=>Filter1_103, outFilter0(102)=>Filter1_102, 
      outFilter0(101)=>Filter1_101, outFilter0(100)=>Filter1_100, 
      outFilter0(99)=>Filter1_99, outFilter0(98)=>Filter1_98, outFilter0(97)
      =>Filter1_97, outFilter0(96)=>Filter1_96, outFilter0(95)=>Filter1_95, 
      outFilter0(94)=>Filter1_94, outFilter0(93)=>Filter1_93, outFilter0(92)
      =>Filter1_92, outFilter0(91)=>Filter1_91, outFilter0(90)=>Filter1_90, 
      outFilter0(89)=>Filter1_89, outFilter0(88)=>Filter1_88, outFilter0(87)
      =>Filter1_87, outFilter0(86)=>Filter1_86, outFilter0(85)=>Filter1_85, 
      outFilter0(84)=>Filter1_84, outFilter0(83)=>Filter1_83, outFilter0(82)
      =>Filter1_82, outFilter0(81)=>Filter1_81, outFilter0(80)=>Filter1_80, 
      outFilter0(79)=>Filter1_79, outFilter0(78)=>Filter1_78, outFilter0(77)
      =>Filter1_77, outFilter0(76)=>Filter1_76, outFilter0(75)=>Filter1_75, 
      outFilter0(74)=>Filter1_74, outFilter0(73)=>Filter1_73, outFilter0(72)
      =>Filter1_72, outFilter0(71)=>Filter1_71, outFilter0(70)=>Filter1_70, 
      outFilter0(69)=>Filter1_69, outFilter0(68)=>Filter1_68, outFilter0(67)
      =>Filter1_67, outFilter0(66)=>Filter1_66, outFilter0(65)=>Filter1_65, 
      outFilter0(64)=>Filter1_64, outFilter0(63)=>Filter1_63, outFilter0(62)
      =>Filter1_62, outFilter0(61)=>Filter1_61, outFilter0(60)=>Filter1_60, 
      outFilter0(59)=>Filter1_59, outFilter0(58)=>Filter1_58, outFilter0(57)
      =>Filter1_57, outFilter0(56)=>Filter1_56, outFilter0(55)=>Filter1_55, 
      outFilter0(54)=>Filter1_54, outFilter0(53)=>Filter1_53, outFilter0(52)
      =>Filter1_52, outFilter0(51)=>Filter1_51, outFilter0(50)=>Filter1_50, 
      outFilter0(49)=>Filter1_49, outFilter0(48)=>Filter1_48, outFilter0(47)
      =>Filter1_47, outFilter0(46)=>Filter1_46, outFilter0(45)=>Filter1_45, 
      outFilter0(44)=>Filter1_44, outFilter0(43)=>Filter1_43, outFilter0(42)
      =>Filter1_42, outFilter0(41)=>Filter1_41, outFilter0(40)=>Filter1_40, 
      outFilter0(39)=>Filter1_39, outFilter0(38)=>Filter1_38, outFilter0(37)
      =>Filter1_37, outFilter0(36)=>Filter1_36, outFilter0(35)=>Filter1_35, 
      outFilter0(34)=>Filter1_34, outFilter0(33)=>Filter1_33, outFilter0(32)
      =>Filter1_32, outFilter0(31)=>Filter1_31, outFilter0(30)=>Filter1_30, 
      outFilter0(29)=>Filter1_29, outFilter0(28)=>Filter1_28, outFilter0(27)
      =>Filter1_27, outFilter0(26)=>Filter1_26, outFilter0(25)=>Filter1_25, 
      outFilter0(24)=>Filter1_24, outFilter0(23)=>Filter1_23, outFilter0(22)
      =>Filter1_22, outFilter0(21)=>Filter1_21, outFilter0(20)=>Filter1_20, 
      outFilter0(19)=>Filter1_19, outFilter0(18)=>Filter1_18, outFilter0(17)
      =>Filter1_17, outFilter0(16)=>Filter1_16, outFilter0(15)=>Filter1_15, 
      outFilter0(14)=>Filter1_14, outFilter0(13)=>Filter1_13, outFilter0(12)
      =>Filter1_12, outFilter0(11)=>Filter1_11, outFilter0(10)=>Filter1_10, 
      outFilter0(9)=>Filter1_9, outFilter0(8)=>Filter1_8, outFilter0(7)=>
      Filter1_7, outFilter0(6)=>Filter1_6, outFilter0(5)=>Filter1_5, 
      outFilter0(4)=>Filter1_4, outFilter0(3)=>Filter1_3, outFilter0(2)=>
      Filter1_2, outFilter0(1)=>Filter1_1, outFilter0(0)=>Filter1_0, 
      outFilter1(399)=>Filter2_399, outFilter1(398)=>Filter2_398, 
      outFilter1(397)=>Filter2_397, outFilter1(396)=>Filter2_396, 
      outFilter1(395)=>Filter2_395, outFilter1(394)=>Filter2_394, 
      outFilter1(393)=>Filter2_393, outFilter1(392)=>Filter2_392, 
      outFilter1(391)=>Filter2_391, outFilter1(390)=>Filter2_390, 
      outFilter1(389)=>Filter2_389, outFilter1(388)=>Filter2_388, 
      outFilter1(387)=>Filter2_387, outFilter1(386)=>Filter2_386, 
      outFilter1(385)=>Filter2_385, outFilter1(384)=>Filter2_384, 
      outFilter1(383)=>Filter2_383, outFilter1(382)=>Filter2_382, 
      outFilter1(381)=>Filter2_381, outFilter1(380)=>Filter2_380, 
      outFilter1(379)=>Filter2_379, outFilter1(378)=>Filter2_378, 
      outFilter1(377)=>Filter2_377, outFilter1(376)=>Filter2_376, 
      outFilter1(375)=>Filter2_375, outFilter1(374)=>Filter2_374, 
      outFilter1(373)=>Filter2_373, outFilter1(372)=>Filter2_372, 
      outFilter1(371)=>Filter2_371, outFilter1(370)=>Filter2_370, 
      outFilter1(369)=>Filter2_369, outFilter1(368)=>Filter2_368, 
      outFilter1(367)=>Filter2_367, outFilter1(366)=>Filter2_366, 
      outFilter1(365)=>Filter2_365, outFilter1(364)=>Filter2_364, 
      outFilter1(363)=>Filter2_363, outFilter1(362)=>Filter2_362, 
      outFilter1(361)=>Filter2_361, outFilter1(360)=>Filter2_360, 
      outFilter1(359)=>Filter2_359, outFilter1(358)=>Filter2_358, 
      outFilter1(357)=>Filter2_357, outFilter1(356)=>Filter2_356, 
      outFilter1(355)=>Filter2_355, outFilter1(354)=>Filter2_354, 
      outFilter1(353)=>Filter2_353, outFilter1(352)=>Filter2_352, 
      outFilter1(351)=>Filter2_351, outFilter1(350)=>Filter2_350, 
      outFilter1(349)=>Filter2_349, outFilter1(348)=>Filter2_348, 
      outFilter1(347)=>Filter2_347, outFilter1(346)=>Filter2_346, 
      outFilter1(345)=>Filter2_345, outFilter1(344)=>Filter2_344, 
      outFilter1(343)=>Filter2_343, outFilter1(342)=>Filter2_342, 
      outFilter1(341)=>Filter2_341, outFilter1(340)=>Filter2_340, 
      outFilter1(339)=>Filter2_339, outFilter1(338)=>Filter2_338, 
      outFilter1(337)=>Filter2_337, outFilter1(336)=>Filter2_336, 
      outFilter1(335)=>Filter2_335, outFilter1(334)=>Filter2_334, 
      outFilter1(333)=>Filter2_333, outFilter1(332)=>Filter2_332, 
      outFilter1(331)=>Filter2_331, outFilter1(330)=>Filter2_330, 
      outFilter1(329)=>Filter2_329, outFilter1(328)=>Filter2_328, 
      outFilter1(327)=>Filter2_327, outFilter1(326)=>Filter2_326, 
      outFilter1(325)=>Filter2_325, outFilter1(324)=>Filter2_324, 
      outFilter1(323)=>Filter2_323, outFilter1(322)=>Filter2_322, 
      outFilter1(321)=>Filter2_321, outFilter1(320)=>Filter2_320, 
      outFilter1(319)=>Filter2_319, outFilter1(318)=>Filter2_318, 
      outFilter1(317)=>Filter2_317, outFilter1(316)=>Filter2_316, 
      outFilter1(315)=>Filter2_315, outFilter1(314)=>Filter2_314, 
      outFilter1(313)=>Filter2_313, outFilter1(312)=>Filter2_312, 
      outFilter1(311)=>Filter2_311, outFilter1(310)=>Filter2_310, 
      outFilter1(309)=>Filter2_309, outFilter1(308)=>Filter2_308, 
      outFilter1(307)=>Filter2_307, outFilter1(306)=>Filter2_306, 
      outFilter1(305)=>Filter2_305, outFilter1(304)=>Filter2_304, 
      outFilter1(303)=>Filter2_303, outFilter1(302)=>Filter2_302, 
      outFilter1(301)=>Filter2_301, outFilter1(300)=>Filter2_300, 
      outFilter1(299)=>Filter2_299, outFilter1(298)=>Filter2_298, 
      outFilter1(297)=>Filter2_297, outFilter1(296)=>Filter2_296, 
      outFilter1(295)=>Filter2_295, outFilter1(294)=>Filter2_294, 
      outFilter1(293)=>Filter2_293, outFilter1(292)=>Filter2_292, 
      outFilter1(291)=>Filter2_291, outFilter1(290)=>Filter2_290, 
      outFilter1(289)=>Filter2_289, outFilter1(288)=>Filter2_288, 
      outFilter1(287)=>Filter2_287, outFilter1(286)=>Filter2_286, 
      outFilter1(285)=>Filter2_285, outFilter1(284)=>Filter2_284, 
      outFilter1(283)=>Filter2_283, outFilter1(282)=>Filter2_282, 
      outFilter1(281)=>Filter2_281, outFilter1(280)=>Filter2_280, 
      outFilter1(279)=>Filter2_279, outFilter1(278)=>Filter2_278, 
      outFilter1(277)=>Filter2_277, outFilter1(276)=>Filter2_276, 
      outFilter1(275)=>Filter2_275, outFilter1(274)=>Filter2_274, 
      outFilter1(273)=>Filter2_273, outFilter1(272)=>Filter2_272, 
      outFilter1(271)=>Filter2_271, outFilter1(270)=>Filter2_270, 
      outFilter1(269)=>Filter2_269, outFilter1(268)=>Filter2_268, 
      outFilter1(267)=>Filter2_267, outFilter1(266)=>Filter2_266, 
      outFilter1(265)=>Filter2_265, outFilter1(264)=>Filter2_264, 
      outFilter1(263)=>Filter2_263, outFilter1(262)=>Filter2_262, 
      outFilter1(261)=>Filter2_261, outFilter1(260)=>Filter2_260, 
      outFilter1(259)=>Filter2_259, outFilter1(258)=>Filter2_258, 
      outFilter1(257)=>Filter2_257, outFilter1(256)=>Filter2_256, 
      outFilter1(255)=>Filter2_255, outFilter1(254)=>Filter2_254, 
      outFilter1(253)=>Filter2_253, outFilter1(252)=>Filter2_252, 
      outFilter1(251)=>Filter2_251, outFilter1(250)=>Filter2_250, 
      outFilter1(249)=>Filter2_249, outFilter1(248)=>Filter2_248, 
      outFilter1(247)=>Filter2_247, outFilter1(246)=>Filter2_246, 
      outFilter1(245)=>Filter2_245, outFilter1(244)=>Filter2_244, 
      outFilter1(243)=>Filter2_243, outFilter1(242)=>Filter2_242, 
      outFilter1(241)=>Filter2_241, outFilter1(240)=>Filter2_240, 
      outFilter1(239)=>Filter2_239, outFilter1(238)=>Filter2_238, 
      outFilter1(237)=>Filter2_237, outFilter1(236)=>Filter2_236, 
      outFilter1(235)=>Filter2_235, outFilter1(234)=>Filter2_234, 
      outFilter1(233)=>Filter2_233, outFilter1(232)=>Filter2_232, 
      outFilter1(231)=>Filter2_231, outFilter1(230)=>Filter2_230, 
      outFilter1(229)=>Filter2_229, outFilter1(228)=>Filter2_228, 
      outFilter1(227)=>Filter2_227, outFilter1(226)=>Filter2_226, 
      outFilter1(225)=>Filter2_225, outFilter1(224)=>Filter2_224, 
      outFilter1(223)=>Filter2_223, outFilter1(222)=>Filter2_222, 
      outFilter1(221)=>Filter2_221, outFilter1(220)=>Filter2_220, 
      outFilter1(219)=>Filter2_219, outFilter1(218)=>Filter2_218, 
      outFilter1(217)=>Filter2_217, outFilter1(216)=>Filter2_216, 
      outFilter1(215)=>Filter2_215, outFilter1(214)=>Filter2_214, 
      outFilter1(213)=>Filter2_213, outFilter1(212)=>Filter2_212, 
      outFilter1(211)=>Filter2_211, outFilter1(210)=>Filter2_210, 
      outFilter1(209)=>Filter2_209, outFilter1(208)=>Filter2_208, 
      outFilter1(207)=>Filter2_207, outFilter1(206)=>Filter2_206, 
      outFilter1(205)=>Filter2_205, outFilter1(204)=>Filter2_204, 
      outFilter1(203)=>Filter2_203, outFilter1(202)=>Filter2_202, 
      outFilter1(201)=>Filter2_201, outFilter1(200)=>Filter2_200, 
      outFilter1(199)=>Filter2_199, outFilter1(198)=>Filter2_198, 
      outFilter1(197)=>Filter2_197, outFilter1(196)=>Filter2_196, 
      outFilter1(195)=>Filter2_195, outFilter1(194)=>Filter2_194, 
      outFilter1(193)=>Filter2_193, outFilter1(192)=>Filter2_192, 
      outFilter1(191)=>Filter2_191, outFilter1(190)=>Filter2_190, 
      outFilter1(189)=>Filter2_189, outFilter1(188)=>Filter2_188, 
      outFilter1(187)=>Filter2_187, outFilter1(186)=>Filter2_186, 
      outFilter1(185)=>Filter2_185, outFilter1(184)=>Filter2_184, 
      outFilter1(183)=>Filter2_183, outFilter1(182)=>Filter2_182, 
      outFilter1(181)=>Filter2_181, outFilter1(180)=>Filter2_180, 
      outFilter1(179)=>Filter2_179, outFilter1(178)=>Filter2_178, 
      outFilter1(177)=>Filter2_177, outFilter1(176)=>Filter2_176, 
      outFilter1(175)=>Filter2_175, outFilter1(174)=>Filter2_174, 
      outFilter1(173)=>Filter2_173, outFilter1(172)=>Filter2_172, 
      outFilter1(171)=>Filter2_171, outFilter1(170)=>Filter2_170, 
      outFilter1(169)=>Filter2_169, outFilter1(168)=>Filter2_168, 
      outFilter1(167)=>Filter2_167, outFilter1(166)=>Filter2_166, 
      outFilter1(165)=>Filter2_165, outFilter1(164)=>Filter2_164, 
      outFilter1(163)=>Filter2_163, outFilter1(162)=>Filter2_162, 
      outFilter1(161)=>Filter2_161, outFilter1(160)=>Filter2_160, 
      outFilter1(159)=>Filter2_159, outFilter1(158)=>Filter2_158, 
      outFilter1(157)=>Filter2_157, outFilter1(156)=>Filter2_156, 
      outFilter1(155)=>Filter2_155, outFilter1(154)=>Filter2_154, 
      outFilter1(153)=>Filter2_153, outFilter1(152)=>Filter2_152, 
      outFilter1(151)=>Filter2_151, outFilter1(150)=>Filter2_150, 
      outFilter1(149)=>Filter2_149, outFilter1(148)=>Filter2_148, 
      outFilter1(147)=>Filter2_147, outFilter1(146)=>Filter2_146, 
      outFilter1(145)=>Filter2_145, outFilter1(144)=>Filter2_144, 
      outFilter1(143)=>Filter2_143, outFilter1(142)=>Filter2_142, 
      outFilter1(141)=>Filter2_141, outFilter1(140)=>Filter2_140, 
      outFilter1(139)=>Filter2_139, outFilter1(138)=>Filter2_138, 
      outFilter1(137)=>Filter2_137, outFilter1(136)=>Filter2_136, 
      outFilter1(135)=>Filter2_135, outFilter1(134)=>Filter2_134, 
      outFilter1(133)=>Filter2_133, outFilter1(132)=>Filter2_132, 
      outFilter1(131)=>Filter2_131, outFilter1(130)=>Filter2_130, 
      outFilter1(129)=>Filter2_129, outFilter1(128)=>Filter2_128, 
      outFilter1(127)=>Filter2_127, outFilter1(126)=>Filter2_126, 
      outFilter1(125)=>Filter2_125, outFilter1(124)=>Filter2_124, 
      outFilter1(123)=>Filter2_123, outFilter1(122)=>Filter2_122, 
      outFilter1(121)=>Filter2_121, outFilter1(120)=>Filter2_120, 
      outFilter1(119)=>Filter2_119, outFilter1(118)=>Filter2_118, 
      outFilter1(117)=>Filter2_117, outFilter1(116)=>Filter2_116, 
      outFilter1(115)=>Filter2_115, outFilter1(114)=>Filter2_114, 
      outFilter1(113)=>Filter2_113, outFilter1(112)=>Filter2_112, 
      outFilter1(111)=>Filter2_111, outFilter1(110)=>Filter2_110, 
      outFilter1(109)=>Filter2_109, outFilter1(108)=>Filter2_108, 
      outFilter1(107)=>Filter2_107, outFilter1(106)=>Filter2_106, 
      outFilter1(105)=>Filter2_105, outFilter1(104)=>Filter2_104, 
      outFilter1(103)=>Filter2_103, outFilter1(102)=>Filter2_102, 
      outFilter1(101)=>Filter2_101, outFilter1(100)=>Filter2_100, 
      outFilter1(99)=>Filter2_99, outFilter1(98)=>Filter2_98, outFilter1(97)
      =>Filter2_97, outFilter1(96)=>Filter2_96, outFilter1(95)=>Filter2_95, 
      outFilter1(94)=>Filter2_94, outFilter1(93)=>Filter2_93, outFilter1(92)
      =>Filter2_92, outFilter1(91)=>Filter2_91, outFilter1(90)=>Filter2_90, 
      outFilter1(89)=>Filter2_89, outFilter1(88)=>Filter2_88, outFilter1(87)
      =>Filter2_87, outFilter1(86)=>Filter2_86, outFilter1(85)=>Filter2_85, 
      outFilter1(84)=>Filter2_84, outFilter1(83)=>Filter2_83, outFilter1(82)
      =>Filter2_82, outFilter1(81)=>Filter2_81, outFilter1(80)=>Filter2_80, 
      outFilter1(79)=>Filter2_79, outFilter1(78)=>Filter2_78, outFilter1(77)
      =>Filter2_77, outFilter1(76)=>Filter2_76, outFilter1(75)=>Filter2_75, 
      outFilter1(74)=>Filter2_74, outFilter1(73)=>Filter2_73, outFilter1(72)
      =>Filter2_72, outFilter1(71)=>Filter2_71, outFilter1(70)=>Filter2_70, 
      outFilter1(69)=>Filter2_69, outFilter1(68)=>Filter2_68, outFilter1(67)
      =>Filter2_67, outFilter1(66)=>Filter2_66, outFilter1(65)=>Filter2_65, 
      outFilter1(64)=>Filter2_64, outFilter1(63)=>Filter2_63, outFilter1(62)
      =>Filter2_62, outFilter1(61)=>Filter2_61, outFilter1(60)=>Filter2_60, 
      outFilter1(59)=>Filter2_59, outFilter1(58)=>Filter2_58, outFilter1(57)
      =>Filter2_57, outFilter1(56)=>Filter2_56, outFilter1(55)=>Filter2_55, 
      outFilter1(54)=>Filter2_54, outFilter1(53)=>Filter2_53, outFilter1(52)
      =>Filter2_52, outFilter1(51)=>Filter2_51, outFilter1(50)=>Filter2_50, 
      outFilter1(49)=>Filter2_49, outFilter1(48)=>Filter2_48, outFilter1(47)
      =>Filter2_47, outFilter1(46)=>Filter2_46, outFilter1(45)=>Filter2_45, 
      outFilter1(44)=>Filter2_44, outFilter1(43)=>Filter2_43, outFilter1(42)
      =>Filter2_42, outFilter1(41)=>Filter2_41, outFilter1(40)=>Filter2_40, 
      outFilter1(39)=>Filter2_39, outFilter1(38)=>Filter2_38, outFilter1(37)
      =>Filter2_37, outFilter1(36)=>Filter2_36, outFilter1(35)=>Filter2_35, 
      outFilter1(34)=>Filter2_34, outFilter1(33)=>Filter2_33, outFilter1(32)
      =>Filter2_32, outFilter1(31)=>Filter2_31, outFilter1(30)=>Filter2_30, 
      outFilter1(29)=>Filter2_29, outFilter1(28)=>Filter2_28, outFilter1(27)
      =>Filter2_27, outFilter1(26)=>Filter2_26, outFilter1(25)=>Filter2_25, 
      outFilter1(24)=>Filter2_24, outFilter1(23)=>Filter2_23, outFilter1(22)
      =>Filter2_22, outFilter1(21)=>Filter2_21, outFilter1(20)=>Filter2_20, 
      outFilter1(19)=>Filter2_19, outFilter1(18)=>Filter2_18, outFilter1(17)
      =>Filter2_17, outFilter1(16)=>Filter2_16, outFilter1(15)=>Filter2_15, 
      outFilter1(14)=>Filter2_14, outFilter1(13)=>Filter2_13, outFilter1(12)
      =>Filter2_12, outFilter1(11)=>Filter2_11, outFilter1(10)=>Filter2_10, 
      outFilter1(9)=>Filter2_9, outFilter1(8)=>Filter2_8, outFilter1(7)=>
      Filter2_7, outFilter1(6)=>Filter2_6, outFilter1(5)=>Filter2_5, 
      outFilter1(4)=>Filter2_4, outFilter1(3)=>Filter2_3, outFilter1(2)=>
      Filter2_2, outFilter1(1)=>Filter2_1, outFilter1(0)=>Filter2_0, 
      donttrust=>DontRstIndicator, LastFilterIND=>lastFilter, LastHeightOut
      =>DANGLING(431), lastDepthOut=>lastDepthOut);
   RImg : ReadImage port map ( WI=>WriteI, current_state(14)=>zero_11, 
      current_state(13)=>zero_11, current_state(12)=>nx9954, 
      current_state(11)=>current_state_11, current_state(10)=>
      current_state_10, current_state(9)=>zero_11, current_state(8)=>
      current_state_8, current_state(7)=>nx9962, current_state(6)=>
      current_state_6, current_state(5)=>current_state_5, current_state(4)=>
      nx9966, current_state(3)=>current_state_3, current_state(2)=>
      current_state_2, current_state(1)=>zero_11, current_state(0)=>zero_11, 
      CLK=>nx10418, RST=>rst, ACK=>nx10026, ImgAddress(12)=>ImgAddRegOut_12, 
      ImgAddress(11)=>ImgAddRegOut_11, ImgAddress(10)=>ImgAddRegOut_10, 
      ImgAddress(9)=>ImgAddRegOut_9, ImgAddress(8)=>ImgAddRegOut_8, 
      ImgAddress(7)=>ImgAddRegOut_7, ImgAddress(6)=>ImgAddRegOut_6, 
      ImgAddress(5)=>ImgAddRegOut_5, ImgAddress(4)=>ImgAddRegOut_4, 
      ImgAddress(3)=>ImgAddRegOut_3, ImgAddress(2)=>ImgAddRegOut_2, 
      ImgAddress(1)=>ImgAddRegOut_1, ImgAddress(0)=>ImgAddRegOut_0, 
      ImgWidth(15)=>ImgWidthOut_15, ImgWidth(14)=>ImgWidthOut_14, 
      ImgWidth(13)=>ImgWidthOut_13, ImgWidth(12)=>ImgWidthOut_12, 
      ImgWidth(11)=>ImgWidthOut_11, ImgWidth(10)=>ImgWidthOut_10, 
      ImgWidth(9)=>ImgWidthOut_9, ImgWidth(8)=>ImgWidthOut_8, ImgWidth(7)=>
      ImgWidthOut_7, ImgWidth(6)=>ImgWidthOut_6, ImgWidth(5)=>ImgWidthOut_5, 
      ImgWidth(4)=>ImgWidthOut_4, ImgWidth(3)=>ImgWidthOut_3, ImgWidth(2)=>
      ImgWidthOut_2, ImgWidth(1)=>ImgWidthOut_1, ImgWidth(0)=>ImgWidthOut_0, 
      DATA(447)=>DataIOut_447, DATA(446)=>DataIOut_446, DATA(445)=>
      DataIOut_445, DATA(444)=>DataIOut_444, DATA(443)=>DataIOut_443, 
      DATA(442)=>DataIOut_442, DATA(441)=>DataIOut_441, DATA(440)=>
      DataIOut_440, DATA(439)=>DataIOut_439, DATA(438)=>DataIOut_438, 
      DATA(437)=>DataIOut_437, DATA(436)=>DataIOut_436, DATA(435)=>
      DataIOut_435, DATA(434)=>DataIOut_434, DATA(433)=>DataIOut_433, 
      DATA(432)=>DataIOut_432, DATA(431)=>DataIOut_431, DATA(430)=>
      DataIOut_430, DATA(429)=>DataIOut_429, DATA(428)=>DataIOut_428, 
      DATA(427)=>DataIOut_427, DATA(426)=>DataIOut_426, DATA(425)=>
      DataIOut_425, DATA(424)=>DataIOut_424, DATA(423)=>DataIOut_423, 
      DATA(422)=>DataIOut_422, DATA(421)=>DataIOut_421, DATA(420)=>
      DataIOut_420, DATA(419)=>DataIOut_419, DATA(418)=>DataIOut_418, 
      DATA(417)=>DataIOut_417, DATA(416)=>DataIOut_416, DATA(415)=>
      DataIOut_415, DATA(414)=>DataIOut_414, DATA(413)=>DataIOut_413, 
      DATA(412)=>DataIOut_412, DATA(411)=>DataIOut_411, DATA(410)=>
      DataIOut_410, DATA(409)=>DataIOut_409, DATA(408)=>DataIOut_408, 
      DATA(407)=>DataIOut_407, DATA(406)=>DataIOut_406, DATA(405)=>
      DataIOut_405, DATA(404)=>DataIOut_404, DATA(403)=>DataIOut_403, 
      DATA(402)=>DataIOut_402, DATA(401)=>DataIOut_401, DATA(400)=>
      DataIOut_400, DATA(399)=>DataIOut_399, DATA(398)=>DataIOut_398, 
      DATA(397)=>DataIOut_397, DATA(396)=>DataIOut_396, DATA(395)=>
      DataIOut_395, DATA(394)=>DataIOut_394, DATA(393)=>DataIOut_393, 
      DATA(392)=>DataIOut_392, DATA(391)=>DataIOut_391, DATA(390)=>
      DataIOut_390, DATA(389)=>DataIOut_389, DATA(388)=>DataIOut_388, 
      DATA(387)=>DataIOut_387, DATA(386)=>DataIOut_386, DATA(385)=>
      DataIOut_385, DATA(384)=>DataIOut_384, DATA(383)=>DataIOut_383, 
      DATA(382)=>DataIOut_382, DATA(381)=>DataIOut_381, DATA(380)=>
      DataIOut_380, DATA(379)=>DataIOut_379, DATA(378)=>DataIOut_378, 
      DATA(377)=>DataIOut_377, DATA(376)=>DataIOut_376, DATA(375)=>
      DataIOut_375, DATA(374)=>DataIOut_374, DATA(373)=>DataIOut_373, 
      DATA(372)=>DataIOut_372, DATA(371)=>DataIOut_371, DATA(370)=>
      DataIOut_370, DATA(369)=>DataIOut_369, DATA(368)=>DataIOut_368, 
      DATA(367)=>DataIOut_367, DATA(366)=>DataIOut_366, DATA(365)=>
      DataIOut_365, DATA(364)=>DataIOut_364, DATA(363)=>DataIOut_363, 
      DATA(362)=>DataIOut_362, DATA(361)=>DataIOut_361, DATA(360)=>
      DataIOut_360, DATA(359)=>DataIOut_359, DATA(358)=>DataIOut_358, 
      DATA(357)=>DataIOut_357, DATA(356)=>DataIOut_356, DATA(355)=>
      DataIOut_355, DATA(354)=>DataIOut_354, DATA(353)=>DataIOut_353, 
      DATA(352)=>DataIOut_352, DATA(351)=>DataIOut_351, DATA(350)=>
      DataIOut_350, DATA(349)=>DataIOut_349, DATA(348)=>DataIOut_348, 
      DATA(347)=>DataIOut_347, DATA(346)=>DataIOut_346, DATA(345)=>
      DataIOut_345, DATA(344)=>DataIOut_344, DATA(343)=>DataIOut_343, 
      DATA(342)=>DataIOut_342, DATA(341)=>DataIOut_341, DATA(340)=>
      DataIOut_340, DATA(339)=>DataIOut_339, DATA(338)=>DataIOut_338, 
      DATA(337)=>DataIOut_337, DATA(336)=>DataIOut_336, DATA(335)=>
      DataIOut_335, DATA(334)=>DataIOut_334, DATA(333)=>DataIOut_333, 
      DATA(332)=>DataIOut_332, DATA(331)=>DataIOut_331, DATA(330)=>
      DataIOut_330, DATA(329)=>DataIOut_329, DATA(328)=>DataIOut_328, 
      DATA(327)=>DataIOut_327, DATA(326)=>DataIOut_326, DATA(325)=>
      DataIOut_325, DATA(324)=>DataIOut_324, DATA(323)=>DataIOut_323, 
      DATA(322)=>DataIOut_322, DATA(321)=>DataIOut_321, DATA(320)=>
      DataIOut_320, DATA(319)=>DataIOut_319, DATA(318)=>DataIOut_318, 
      DATA(317)=>DataIOut_317, DATA(316)=>DataIOut_316, DATA(315)=>
      DataIOut_315, DATA(314)=>DataIOut_314, DATA(313)=>DataIOut_313, 
      DATA(312)=>DataIOut_312, DATA(311)=>DataIOut_311, DATA(310)=>
      DataIOut_310, DATA(309)=>DataIOut_309, DATA(308)=>DataIOut_308, 
      DATA(307)=>DataIOut_307, DATA(306)=>DataIOut_306, DATA(305)=>
      DataIOut_305, DATA(304)=>DataIOut_304, DATA(303)=>DataIOut_303, 
      DATA(302)=>DataIOut_302, DATA(301)=>DataIOut_301, DATA(300)=>
      DataIOut_300, DATA(299)=>DataIOut_299, DATA(298)=>DataIOut_298, 
      DATA(297)=>DataIOut_297, DATA(296)=>DataIOut_296, DATA(295)=>
      DataIOut_295, DATA(294)=>DataIOut_294, DATA(293)=>DataIOut_293, 
      DATA(292)=>DataIOut_292, DATA(291)=>DataIOut_291, DATA(290)=>
      DataIOut_290, DATA(289)=>DataIOut_289, DATA(288)=>DataIOut_288, 
      DATA(287)=>DataIOut_287, DATA(286)=>DataIOut_286, DATA(285)=>
      DataIOut_285, DATA(284)=>DataIOut_284, DATA(283)=>DataIOut_283, 
      DATA(282)=>DataIOut_282, DATA(281)=>DataIOut_281, DATA(280)=>
      DataIOut_280, DATA(279)=>DataIOut_279, DATA(278)=>DataIOut_278, 
      DATA(277)=>DataIOut_277, DATA(276)=>DataIOut_276, DATA(275)=>
      DataIOut_275, DATA(274)=>DataIOut_274, DATA(273)=>DataIOut_273, 
      DATA(272)=>DataIOut_272, DATA(271)=>DataIOut_271, DATA(270)=>
      DataIOut_270, DATA(269)=>DataIOut_269, DATA(268)=>DataIOut_268, 
      DATA(267)=>DataIOut_267, DATA(266)=>DataIOut_266, DATA(265)=>
      DataIOut_265, DATA(264)=>DataIOut_264, DATA(263)=>DataIOut_263, 
      DATA(262)=>DataIOut_262, DATA(261)=>DataIOut_261, DATA(260)=>
      DataIOut_260, DATA(259)=>DataIOut_259, DATA(258)=>DataIOut_258, 
      DATA(257)=>DataIOut_257, DATA(256)=>DataIOut_256, DATA(255)=>
      DataIOut_255, DATA(254)=>DataIOut_254, DATA(253)=>DataIOut_253, 
      DATA(252)=>DataIOut_252, DATA(251)=>DataIOut_251, DATA(250)=>
      DataIOut_250, DATA(249)=>DataIOut_249, DATA(248)=>DataIOut_248, 
      DATA(247)=>DataIOut_247, DATA(246)=>DataIOut_246, DATA(245)=>
      DataIOut_245, DATA(244)=>DataIOut_244, DATA(243)=>DataIOut_243, 
      DATA(242)=>DataIOut_242, DATA(241)=>DataIOut_241, DATA(240)=>
      DataIOut_240, DATA(239)=>DataIOut_239, DATA(238)=>DataIOut_238, 
      DATA(237)=>DataIOut_237, DATA(236)=>DataIOut_236, DATA(235)=>
      DataIOut_235, DATA(234)=>DataIOut_234, DATA(233)=>DataIOut_233, 
      DATA(232)=>DataIOut_232, DATA(231)=>DataIOut_231, DATA(230)=>
      DataIOut_230, DATA(229)=>DataIOut_229, DATA(228)=>DataIOut_228, 
      DATA(227)=>DataIOut_227, DATA(226)=>DataIOut_226, DATA(225)=>
      DataIOut_225, DATA(224)=>DataIOut_224, DATA(223)=>DataIOut_223, 
      DATA(222)=>DataIOut_222, DATA(221)=>DataIOut_221, DATA(220)=>
      DataIOut_220, DATA(219)=>DataIOut_219, DATA(218)=>DataIOut_218, 
      DATA(217)=>DataIOut_217, DATA(216)=>DataIOut_216, DATA(215)=>
      DataIOut_215, DATA(214)=>DataIOut_214, DATA(213)=>DataIOut_213, 
      DATA(212)=>DataIOut_212, DATA(211)=>DataIOut_211, DATA(210)=>
      DataIOut_210, DATA(209)=>DataIOut_209, DATA(208)=>DataIOut_208, 
      DATA(207)=>DataIOut_207, DATA(206)=>DataIOut_206, DATA(205)=>
      DataIOut_205, DATA(204)=>DataIOut_204, DATA(203)=>DataIOut_203, 
      DATA(202)=>DataIOut_202, DATA(201)=>DataIOut_201, DATA(200)=>
      DataIOut_200, DATA(199)=>DataIOut_199, DATA(198)=>DataIOut_198, 
      DATA(197)=>DataIOut_197, DATA(196)=>DataIOut_196, DATA(195)=>
      DataIOut_195, DATA(194)=>DataIOut_194, DATA(193)=>DataIOut_193, 
      DATA(192)=>DataIOut_192, DATA(191)=>DataIOut_191, DATA(190)=>
      DataIOut_190, DATA(189)=>DataIOut_189, DATA(188)=>DataIOut_188, 
      DATA(187)=>DataIOut_187, DATA(186)=>DataIOut_186, DATA(185)=>
      DataIOut_185, DATA(184)=>DataIOut_184, DATA(183)=>DataIOut_183, 
      DATA(182)=>DataIOut_182, DATA(181)=>DataIOut_181, DATA(180)=>
      DataIOut_180, DATA(179)=>DataIOut_179, DATA(178)=>DataIOut_178, 
      DATA(177)=>DataIOut_177, DATA(176)=>DataIOut_176, DATA(175)=>
      DataIOut_175, DATA(174)=>DataIOut_174, DATA(173)=>DataIOut_173, 
      DATA(172)=>DataIOut_172, DATA(171)=>DataIOut_171, DATA(170)=>
      DataIOut_170, DATA(169)=>DataIOut_169, DATA(168)=>DataIOut_168, 
      DATA(167)=>DataIOut_167, DATA(166)=>DataIOut_166, DATA(165)=>
      DataIOut_165, DATA(164)=>DataIOut_164, DATA(163)=>DataIOut_163, 
      DATA(162)=>DataIOut_162, DATA(161)=>DataIOut_161, DATA(160)=>
      DataIOut_160, DATA(159)=>DataIOut_159, DATA(158)=>DataIOut_158, 
      DATA(157)=>DataIOut_157, DATA(156)=>DataIOut_156, DATA(155)=>
      DataIOut_155, DATA(154)=>DataIOut_154, DATA(153)=>DataIOut_153, 
      DATA(152)=>DataIOut_152, DATA(151)=>DataIOut_151, DATA(150)=>
      DataIOut_150, DATA(149)=>DataIOut_149, DATA(148)=>DataIOut_148, 
      DATA(147)=>DataIOut_147, DATA(146)=>DataIOut_146, DATA(145)=>
      DataIOut_145, DATA(144)=>DataIOut_144, DATA(143)=>DataIOut_143, 
      DATA(142)=>DataIOut_142, DATA(141)=>DataIOut_141, DATA(140)=>
      DataIOut_140, DATA(139)=>DataIOut_139, DATA(138)=>DataIOut_138, 
      DATA(137)=>DataIOut_137, DATA(136)=>DataIOut_136, DATA(135)=>
      DataIOut_135, DATA(134)=>DataIOut_134, DATA(133)=>DataIOut_133, 
      DATA(132)=>DataIOut_132, DATA(131)=>DataIOut_131, DATA(130)=>
      DataIOut_130, DATA(129)=>DataIOut_129, DATA(128)=>DataIOut_128, 
      DATA(127)=>DataIOut_127, DATA(126)=>DataIOut_126, DATA(125)=>
      DataIOut_125, DATA(124)=>DataIOut_124, DATA(123)=>DataIOut_123, 
      DATA(122)=>DataIOut_122, DATA(121)=>DataIOut_121, DATA(120)=>
      DataIOut_120, DATA(119)=>DataIOut_119, DATA(118)=>DataIOut_118, 
      DATA(117)=>DataIOut_117, DATA(116)=>DataIOut_116, DATA(115)=>
      DataIOut_115, DATA(114)=>DataIOut_114, DATA(113)=>DataIOut_113, 
      DATA(112)=>DataIOut_112, DATA(111)=>DataIOut_111, DATA(110)=>
      DataIOut_110, DATA(109)=>DataIOut_109, DATA(108)=>DataIOut_108, 
      DATA(107)=>DataIOut_107, DATA(106)=>DataIOut_106, DATA(105)=>
      DataIOut_105, DATA(104)=>DataIOut_104, DATA(103)=>DataIOut_103, 
      DATA(102)=>DataIOut_102, DATA(101)=>DataIOut_101, DATA(100)=>
      DataIOut_100, DATA(99)=>DataIOut_99, DATA(98)=>DataIOut_98, DATA(97)=>
      DataIOut_97, DATA(96)=>DataIOut_96, DATA(95)=>DataIOut_95, DATA(94)=>
      DataIOut_94, DATA(93)=>DataIOut_93, DATA(92)=>DataIOut_92, DATA(91)=>
      DataIOut_91, DATA(90)=>DataIOut_90, DATA(89)=>DataIOut_89, DATA(88)=>
      DataIOut_88, DATA(87)=>DataIOut_87, DATA(86)=>DataIOut_86, DATA(85)=>
      DataIOut_85, DATA(84)=>DataIOut_84, DATA(83)=>DataIOut_83, DATA(82)=>
      DataIOut_82, DATA(81)=>DataIOut_81, DATA(80)=>DataIOut_80, DATA(79)=>
      DataIOut_79, DATA(78)=>DataIOut_78, DATA(77)=>DataIOut_77, DATA(76)=>
      DataIOut_76, DATA(75)=>DataIOut_75, DATA(74)=>DataIOut_74, DATA(73)=>
      DataIOut_73, DATA(72)=>DataIOut_72, DATA(71)=>DataIOut_71, DATA(70)=>
      DataIOut_70, DATA(69)=>DataIOut_69, DATA(68)=>DataIOut_68, DATA(67)=>
      DataIOut_67, DATA(66)=>DataIOut_66, DATA(65)=>DataIOut_65, DATA(64)=>
      DataIOut_64, DATA(63)=>DataIOut_63, DATA(62)=>DataIOut_62, DATA(61)=>
      DataIOut_61, DATA(60)=>DataIOut_60, DATA(59)=>DataIOut_59, DATA(58)=>
      DataIOut_58, DATA(57)=>DataIOut_57, DATA(56)=>DataIOut_56, DATA(55)=>
      DataIOut_55, DATA(54)=>DataIOut_54, DATA(53)=>DataIOut_53, DATA(52)=>
      DataIOut_52, DATA(51)=>DataIOut_51, DATA(50)=>DataIOut_50, DATA(49)=>
      DataIOut_49, DATA(48)=>DataIOut_48, DATA(47)=>DataIOut_47, DATA(46)=>
      DataIOut_46, DATA(45)=>DataIOut_45, DATA(44)=>DataIOut_44, DATA(43)=>
      DataIOut_43, DATA(42)=>DataIOut_42, DATA(41)=>DataIOut_41, DATA(40)=>
      DataIOut_40, DATA(39)=>DataIOut_39, DATA(38)=>DataIOut_38, DATA(37)=>
      DataIOut_37, DATA(36)=>DataIOut_36, DATA(35)=>DataIOut_35, DATA(34)=>
      DataIOut_34, DATA(33)=>DataIOut_33, DATA(32)=>DataIOut_32, DATA(31)=>
      DataIOut_31, DATA(30)=>DataIOut_30, DATA(29)=>DataIOut_29, DATA(28)=>
      DataIOut_28, DATA(27)=>DataIOut_27, DATA(26)=>DataIOut_26, DATA(25)=>
      DataIOut_25, DATA(24)=>DataIOut_24, DATA(23)=>DataIOut_23, DATA(22)=>
      DataIOut_22, DATA(21)=>DataIOut_21, DATA(20)=>DataIOut_20, DATA(19)=>
      DataIOut_19, DATA(18)=>DataIOut_18, DATA(17)=>DataIOut_17, DATA(16)=>
      DataIOut_16, DATA(15)=>nx10312, DATA(14)=>nx10316, DATA(13)=>nx10320, 
      DATA(12)=>nx10324, DATA(11)=>nx10328, DATA(10)=>nx10332, DATA(9)=>
      nx10336, DATA(8)=>nx10340, DATA(7)=>nx10344, DATA(6)=>nx10348, DATA(5)
      =>nx10352, DATA(4)=>nx10356, DATA(3)=>nx10360, DATA(2)=>nx10364, 
      DATA(1)=>nx10368, DATA(0)=>nx10372, OutputImg0(447)=>DANGLING(432), 
      OutputImg0(446)=>DANGLING(433), OutputImg0(445)=>DANGLING(434), 
      OutputImg0(444)=>DANGLING(435), OutputImg0(443)=>DANGLING(436), 
      OutputImg0(442)=>DANGLING(437), OutputImg0(441)=>DANGLING(438), 
      OutputImg0(440)=>DANGLING(439), OutputImg0(439)=>DANGLING(440), 
      OutputImg0(438)=>DANGLING(441), OutputImg0(437)=>DANGLING(442), 
      OutputImg0(436)=>DANGLING(443), OutputImg0(435)=>DANGLING(444), 
      OutputImg0(434)=>DANGLING(445), OutputImg0(433)=>DANGLING(446), 
      OutputImg0(432)=>DANGLING(447), OutputImg0(431)=>DANGLING(448), 
      OutputImg0(430)=>DANGLING(449), OutputImg0(429)=>DANGLING(450), 
      OutputImg0(428)=>DANGLING(451), OutputImg0(427)=>DANGLING(452), 
      OutputImg0(426)=>DANGLING(453), OutputImg0(425)=>DANGLING(454), 
      OutputImg0(424)=>DANGLING(455), OutputImg0(423)=>DANGLING(456), 
      OutputImg0(422)=>DANGLING(457), OutputImg0(421)=>DANGLING(458), 
      OutputImg0(420)=>DANGLING(459), OutputImg0(419)=>DANGLING(460), 
      OutputImg0(418)=>DANGLING(461), OutputImg0(417)=>DANGLING(462), 
      OutputImg0(416)=>DANGLING(463), OutputImg0(415)=>DANGLING(464), 
      OutputImg0(414)=>DANGLING(465), OutputImg0(413)=>DANGLING(466), 
      OutputImg0(412)=>DANGLING(467), OutputImg0(411)=>DANGLING(468), 
      OutputImg0(410)=>DANGLING(469), OutputImg0(409)=>DANGLING(470), 
      OutputImg0(408)=>DANGLING(471), OutputImg0(407)=>DANGLING(472), 
      OutputImg0(406)=>DANGLING(473), OutputImg0(405)=>DANGLING(474), 
      OutputImg0(404)=>DANGLING(475), OutputImg0(403)=>DANGLING(476), 
      OutputImg0(402)=>DANGLING(477), OutputImg0(401)=>DANGLING(478), 
      OutputImg0(400)=>DANGLING(479), OutputImg0(399)=>DANGLING(480), 
      OutputImg0(398)=>DANGLING(481), OutputImg0(397)=>DANGLING(482), 
      OutputImg0(396)=>DANGLING(483), OutputImg0(395)=>DANGLING(484), 
      OutputImg0(394)=>DANGLING(485), OutputImg0(393)=>DANGLING(486), 
      OutputImg0(392)=>DANGLING(487), OutputImg0(391)=>DANGLING(488), 
      OutputImg0(390)=>DANGLING(489), OutputImg0(389)=>DANGLING(490), 
      OutputImg0(388)=>DANGLING(491), OutputImg0(387)=>DANGLING(492), 
      OutputImg0(386)=>DANGLING(493), OutputImg0(385)=>DANGLING(494), 
      OutputImg0(384)=>DANGLING(495), OutputImg0(383)=>DANGLING(496), 
      OutputImg0(382)=>DANGLING(497), OutputImg0(381)=>DANGLING(498), 
      OutputImg0(380)=>DANGLING(499), OutputImg0(379)=>DANGLING(500), 
      OutputImg0(378)=>DANGLING(501), OutputImg0(377)=>DANGLING(502), 
      OutputImg0(376)=>DANGLING(503), OutputImg0(375)=>DANGLING(504), 
      OutputImg0(374)=>DANGLING(505), OutputImg0(373)=>DANGLING(506), 
      OutputImg0(372)=>DANGLING(507), OutputImg0(371)=>DANGLING(508), 
      OutputImg0(370)=>DANGLING(509), OutputImg0(369)=>DANGLING(510), 
      OutputImg0(368)=>DANGLING(511), OutputImg0(367)=>DANGLING(512), 
      OutputImg0(366)=>DANGLING(513), OutputImg0(365)=>DANGLING(514), 
      OutputImg0(364)=>DANGLING(515), OutputImg0(363)=>DANGLING(516), 
      OutputImg0(362)=>DANGLING(517), OutputImg0(361)=>DANGLING(518), 
      OutputImg0(360)=>DANGLING(519), OutputImg0(359)=>DANGLING(520), 
      OutputImg0(358)=>DANGLING(521), OutputImg0(357)=>DANGLING(522), 
      OutputImg0(356)=>DANGLING(523), OutputImg0(355)=>DANGLING(524), 
      OutputImg0(354)=>DANGLING(525), OutputImg0(353)=>DANGLING(526), 
      OutputImg0(352)=>DANGLING(527), OutputImg0(351)=>DANGLING(528), 
      OutputImg0(350)=>DANGLING(529), OutputImg0(349)=>DANGLING(530), 
      OutputImg0(348)=>DANGLING(531), OutputImg0(347)=>DANGLING(532), 
      OutputImg0(346)=>DANGLING(533), OutputImg0(345)=>DANGLING(534), 
      OutputImg0(344)=>DANGLING(535), OutputImg0(343)=>DANGLING(536), 
      OutputImg0(342)=>DANGLING(537), OutputImg0(341)=>DANGLING(538), 
      OutputImg0(340)=>DANGLING(539), OutputImg0(339)=>DANGLING(540), 
      OutputImg0(338)=>DANGLING(541), OutputImg0(337)=>DANGLING(542), 
      OutputImg0(336)=>DANGLING(543), OutputImg0(335)=>DANGLING(544), 
      OutputImg0(334)=>DANGLING(545), OutputImg0(333)=>DANGLING(546), 
      OutputImg0(332)=>DANGLING(547), OutputImg0(331)=>DANGLING(548), 
      OutputImg0(330)=>DANGLING(549), OutputImg0(329)=>DANGLING(550), 
      OutputImg0(328)=>DANGLING(551), OutputImg0(327)=>DANGLING(552), 
      OutputImg0(326)=>DANGLING(553), OutputImg0(325)=>DANGLING(554), 
      OutputImg0(324)=>DANGLING(555), OutputImg0(323)=>DANGLING(556), 
      OutputImg0(322)=>DANGLING(557), OutputImg0(321)=>DANGLING(558), 
      OutputImg0(320)=>DANGLING(559), OutputImg0(319)=>DANGLING(560), 
      OutputImg0(318)=>DANGLING(561), OutputImg0(317)=>DANGLING(562), 
      OutputImg0(316)=>DANGLING(563), OutputImg0(315)=>DANGLING(564), 
      OutputImg0(314)=>DANGLING(565), OutputImg0(313)=>DANGLING(566), 
      OutputImg0(312)=>DANGLING(567), OutputImg0(311)=>DANGLING(568), 
      OutputImg0(310)=>DANGLING(569), OutputImg0(309)=>DANGLING(570), 
      OutputImg0(308)=>DANGLING(571), OutputImg0(307)=>DANGLING(572), 
      OutputImg0(306)=>DANGLING(573), OutputImg0(305)=>DANGLING(574), 
      OutputImg0(304)=>DANGLING(575), OutputImg0(303)=>DANGLING(576), 
      OutputImg0(302)=>DANGLING(577), OutputImg0(301)=>DANGLING(578), 
      OutputImg0(300)=>DANGLING(579), OutputImg0(299)=>DANGLING(580), 
      OutputImg0(298)=>DANGLING(581), OutputImg0(297)=>DANGLING(582), 
      OutputImg0(296)=>DANGLING(583), OutputImg0(295)=>DANGLING(584), 
      OutputImg0(294)=>DANGLING(585), OutputImg0(293)=>DANGLING(586), 
      OutputImg0(292)=>DANGLING(587), OutputImg0(291)=>DANGLING(588), 
      OutputImg0(290)=>DANGLING(589), OutputImg0(289)=>DANGLING(590), 
      OutputImg0(288)=>DANGLING(591), OutputImg0(287)=>DANGLING(592), 
      OutputImg0(286)=>DANGLING(593), OutputImg0(285)=>DANGLING(594), 
      OutputImg0(284)=>DANGLING(595), OutputImg0(283)=>DANGLING(596), 
      OutputImg0(282)=>DANGLING(597), OutputImg0(281)=>DANGLING(598), 
      OutputImg0(280)=>DANGLING(599), OutputImg0(279)=>DANGLING(600), 
      OutputImg0(278)=>DANGLING(601), OutputImg0(277)=>DANGLING(602), 
      OutputImg0(276)=>DANGLING(603), OutputImg0(275)=>DANGLING(604), 
      OutputImg0(274)=>DANGLING(605), OutputImg0(273)=>DANGLING(606), 
      OutputImg0(272)=>DANGLING(607), OutputImg0(271)=>DANGLING(608), 
      OutputImg0(270)=>DANGLING(609), OutputImg0(269)=>DANGLING(610), 
      OutputImg0(268)=>DANGLING(611), OutputImg0(267)=>DANGLING(612), 
      OutputImg0(266)=>DANGLING(613), OutputImg0(265)=>DANGLING(614), 
      OutputImg0(264)=>DANGLING(615), OutputImg0(263)=>DANGLING(616), 
      OutputImg0(262)=>DANGLING(617), OutputImg0(261)=>DANGLING(618), 
      OutputImg0(260)=>DANGLING(619), OutputImg0(259)=>DANGLING(620), 
      OutputImg0(258)=>DANGLING(621), OutputImg0(257)=>DANGLING(622), 
      OutputImg0(256)=>DANGLING(623), OutputImg0(255)=>DANGLING(624), 
      OutputImg0(254)=>DANGLING(625), OutputImg0(253)=>DANGLING(626), 
      OutputImg0(252)=>DANGLING(627), OutputImg0(251)=>DANGLING(628), 
      OutputImg0(250)=>DANGLING(629), OutputImg0(249)=>DANGLING(630), 
      OutputImg0(248)=>DANGLING(631), OutputImg0(247)=>DANGLING(632), 
      OutputImg0(246)=>DANGLING(633), OutputImg0(245)=>DANGLING(634), 
      OutputImg0(244)=>DANGLING(635), OutputImg0(243)=>DANGLING(636), 
      OutputImg0(242)=>DANGLING(637), OutputImg0(241)=>DANGLING(638), 
      OutputImg0(240)=>DANGLING(639), OutputImg0(239)=>DANGLING(640), 
      OutputImg0(238)=>DANGLING(641), OutputImg0(237)=>DANGLING(642), 
      OutputImg0(236)=>DANGLING(643), OutputImg0(235)=>DANGLING(644), 
      OutputImg0(234)=>DANGLING(645), OutputImg0(233)=>DANGLING(646), 
      OutputImg0(232)=>DANGLING(647), OutputImg0(231)=>DANGLING(648), 
      OutputImg0(230)=>DANGLING(649), OutputImg0(229)=>DANGLING(650), 
      OutputImg0(228)=>DANGLING(651), OutputImg0(227)=>DANGLING(652), 
      OutputImg0(226)=>DANGLING(653), OutputImg0(225)=>DANGLING(654), 
      OutputImg0(224)=>DANGLING(655), OutputImg0(223)=>DANGLING(656), 
      OutputImg0(222)=>DANGLING(657), OutputImg0(221)=>DANGLING(658), 
      OutputImg0(220)=>DANGLING(659), OutputImg0(219)=>DANGLING(660), 
      OutputImg0(218)=>DANGLING(661), OutputImg0(217)=>DANGLING(662), 
      OutputImg0(216)=>DANGLING(663), OutputImg0(215)=>DANGLING(664), 
      OutputImg0(214)=>DANGLING(665), OutputImg0(213)=>DANGLING(666), 
      OutputImg0(212)=>DANGLING(667), OutputImg0(211)=>DANGLING(668), 
      OutputImg0(210)=>DANGLING(669), OutputImg0(209)=>DANGLING(670), 
      OutputImg0(208)=>DANGLING(671), OutputImg0(207)=>DANGLING(672), 
      OutputImg0(206)=>DANGLING(673), OutputImg0(205)=>DANGLING(674), 
      OutputImg0(204)=>DANGLING(675), OutputImg0(203)=>DANGLING(676), 
      OutputImg0(202)=>DANGLING(677), OutputImg0(201)=>DANGLING(678), 
      OutputImg0(200)=>DANGLING(679), OutputImg0(199)=>DANGLING(680), 
      OutputImg0(198)=>DANGLING(681), OutputImg0(197)=>DANGLING(682), 
      OutputImg0(196)=>DANGLING(683), OutputImg0(195)=>DANGLING(684), 
      OutputImg0(194)=>DANGLING(685), OutputImg0(193)=>DANGLING(686), 
      OutputImg0(192)=>DANGLING(687), OutputImg0(191)=>DANGLING(688), 
      OutputImg0(190)=>DANGLING(689), OutputImg0(189)=>DANGLING(690), 
      OutputImg0(188)=>DANGLING(691), OutputImg0(187)=>DANGLING(692), 
      OutputImg0(186)=>DANGLING(693), OutputImg0(185)=>DANGLING(694), 
      OutputImg0(184)=>DANGLING(695), OutputImg0(183)=>DANGLING(696), 
      OutputImg0(182)=>DANGLING(697), OutputImg0(181)=>DANGLING(698), 
      OutputImg0(180)=>DANGLING(699), OutputImg0(179)=>DANGLING(700), 
      OutputImg0(178)=>DANGLING(701), OutputImg0(177)=>DANGLING(702), 
      OutputImg0(176)=>DANGLING(703), OutputImg0(175)=>DANGLING(704), 
      OutputImg0(174)=>DANGLING(705), OutputImg0(173)=>DANGLING(706), 
      OutputImg0(172)=>DANGLING(707), OutputImg0(171)=>DANGLING(708), 
      OutputImg0(170)=>DANGLING(709), OutputImg0(169)=>DANGLING(710), 
      OutputImg0(168)=>DANGLING(711), OutputImg0(167)=>DANGLING(712), 
      OutputImg0(166)=>DANGLING(713), OutputImg0(165)=>DANGLING(714), 
      OutputImg0(164)=>DANGLING(715), OutputImg0(163)=>DANGLING(716), 
      OutputImg0(162)=>DANGLING(717), OutputImg0(161)=>DANGLING(718), 
      OutputImg0(160)=>DANGLING(719), OutputImg0(159)=>DANGLING(720), 
      OutputImg0(158)=>DANGLING(721), OutputImg0(157)=>DANGLING(722), 
      OutputImg0(156)=>DANGLING(723), OutputImg0(155)=>DANGLING(724), 
      OutputImg0(154)=>DANGLING(725), OutputImg0(153)=>DANGLING(726), 
      OutputImg0(152)=>DANGLING(727), OutputImg0(151)=>DANGLING(728), 
      OutputImg0(150)=>DANGLING(729), OutputImg0(149)=>DANGLING(730), 
      OutputImg0(148)=>DANGLING(731), OutputImg0(147)=>DANGLING(732), 
      OutputImg0(146)=>DANGLING(733), OutputImg0(145)=>DANGLING(734), 
      OutputImg0(144)=>DANGLING(735), OutputImg0(143)=>DANGLING(736), 
      OutputImg0(142)=>DANGLING(737), OutputImg0(141)=>DANGLING(738), 
      OutputImg0(140)=>DANGLING(739), OutputImg0(139)=>DANGLING(740), 
      OutputImg0(138)=>DANGLING(741), OutputImg0(137)=>DANGLING(742), 
      OutputImg0(136)=>DANGLING(743), OutputImg0(135)=>DANGLING(744), 
      OutputImg0(134)=>DANGLING(745), OutputImg0(133)=>DANGLING(746), 
      OutputImg0(132)=>DANGLING(747), OutputImg0(131)=>DANGLING(748), 
      OutputImg0(130)=>DANGLING(749), OutputImg0(129)=>DANGLING(750), 
      OutputImg0(128)=>DANGLING(751), OutputImg0(127)=>DANGLING(752), 
      OutputImg0(126)=>DANGLING(753), OutputImg0(125)=>DANGLING(754), 
      OutputImg0(124)=>DANGLING(755), OutputImg0(123)=>DANGLING(756), 
      OutputImg0(122)=>DANGLING(757), OutputImg0(121)=>DANGLING(758), 
      OutputImg0(120)=>DANGLING(759), OutputImg0(119)=>DANGLING(760), 
      OutputImg0(118)=>DANGLING(761), OutputImg0(117)=>DANGLING(762), 
      OutputImg0(116)=>DANGLING(763), OutputImg0(115)=>DANGLING(764), 
      OutputImg0(114)=>DANGLING(765), OutputImg0(113)=>DANGLING(766), 
      OutputImg0(112)=>DANGLING(767), OutputImg0(111)=>DANGLING(768), 
      OutputImg0(110)=>DANGLING(769), OutputImg0(109)=>DANGLING(770), 
      OutputImg0(108)=>DANGLING(771), OutputImg0(107)=>DANGLING(772), 
      OutputImg0(106)=>DANGLING(773), OutputImg0(105)=>DANGLING(774), 
      OutputImg0(104)=>DANGLING(775), OutputImg0(103)=>DANGLING(776), 
      OutputImg0(102)=>DANGLING(777), OutputImg0(101)=>DANGLING(778), 
      OutputImg0(100)=>DANGLING(779), OutputImg0(99)=>DANGLING(780), 
      OutputImg0(98)=>DANGLING(781), OutputImg0(97)=>DANGLING(782), 
      OutputImg0(96)=>DANGLING(783), OutputImg0(95)=>DANGLING(784), 
      OutputImg0(94)=>DANGLING(785), OutputImg0(93)=>DANGLING(786), 
      OutputImg0(92)=>DANGLING(787), OutputImg0(91)=>DANGLING(788), 
      OutputImg0(90)=>DANGLING(789), OutputImg0(89)=>DANGLING(790), 
      OutputImg0(88)=>DANGLING(791), OutputImg0(87)=>DANGLING(792), 
      OutputImg0(86)=>DANGLING(793), OutputImg0(85)=>DANGLING(794), 
      OutputImg0(84)=>DANGLING(795), OutputImg0(83)=>DANGLING(796), 
      OutputImg0(82)=>DANGLING(797), OutputImg0(81)=>DANGLING(798), 
      OutputImg0(80)=>DANGLING(799), OutputImg0(79)=>OutputImg0_79, 
      OutputImg0(78)=>OutputImg0_78, OutputImg0(77)=>OutputImg0_77, 
      OutputImg0(76)=>OutputImg0_76, OutputImg0(75)=>OutputImg0_75, 
      OutputImg0(74)=>OutputImg0_74, OutputImg0(73)=>OutputImg0_73, 
      OutputImg0(72)=>OutputImg0_72, OutputImg0(71)=>OutputImg0_71, 
      OutputImg0(70)=>OutputImg0_70, OutputImg0(69)=>OutputImg0_69, 
      OutputImg0(68)=>OutputImg0_68, OutputImg0(67)=>OutputImg0_67, 
      OutputImg0(66)=>OutputImg0_66, OutputImg0(65)=>OutputImg0_65, 
      OutputImg0(64)=>OutputImg0_64, OutputImg0(63)=>OutputImg0_63, 
      OutputImg0(62)=>OutputImg0_62, OutputImg0(61)=>OutputImg0_61, 
      OutputImg0(60)=>OutputImg0_60, OutputImg0(59)=>OutputImg0_59, 
      OutputImg0(58)=>OutputImg0_58, OutputImg0(57)=>OutputImg0_57, 
      OutputImg0(56)=>OutputImg0_56, OutputImg0(55)=>OutputImg0_55, 
      OutputImg0(54)=>OutputImg0_54, OutputImg0(53)=>OutputImg0_53, 
      OutputImg0(52)=>OutputImg0_52, OutputImg0(51)=>OutputImg0_51, 
      OutputImg0(50)=>OutputImg0_50, OutputImg0(49)=>OutputImg0_49, 
      OutputImg0(48)=>OutputImg0_48, OutputImg0(47)=>OutputImg0_47, 
      OutputImg0(46)=>OutputImg0_46, OutputImg0(45)=>OutputImg0_45, 
      OutputImg0(44)=>OutputImg0_44, OutputImg0(43)=>OutputImg0_43, 
      OutputImg0(42)=>OutputImg0_42, OutputImg0(41)=>OutputImg0_41, 
      OutputImg0(40)=>OutputImg0_40, OutputImg0(39)=>OutputImg0_39, 
      OutputImg0(38)=>OutputImg0_38, OutputImg0(37)=>OutputImg0_37, 
      OutputImg0(36)=>OutputImg0_36, OutputImg0(35)=>OutputImg0_35, 
      OutputImg0(34)=>OutputImg0_34, OutputImg0(33)=>OutputImg0_33, 
      OutputImg0(32)=>OutputImg0_32, OutputImg0(31)=>OutputImg0_31, 
      OutputImg0(30)=>OutputImg0_30, OutputImg0(29)=>OutputImg0_29, 
      OutputImg0(28)=>OutputImg0_28, OutputImg0(27)=>OutputImg0_27, 
      OutputImg0(26)=>OutputImg0_26, OutputImg0(25)=>OutputImg0_25, 
      OutputImg0(24)=>OutputImg0_24, OutputImg0(23)=>OutputImg0_23, 
      OutputImg0(22)=>OutputImg0_22, OutputImg0(21)=>OutputImg0_21, 
      OutputImg0(20)=>OutputImg0_20, OutputImg0(19)=>OutputImg0_19, 
      OutputImg0(18)=>OutputImg0_18, OutputImg0(17)=>OutputImg0_17, 
      OutputImg0(16)=>OutputImg0_16, OutputImg0(15)=>OutputImg0_15, 
      OutputImg0(14)=>OutputImg0_14, OutputImg0(13)=>OutputImg0_13, 
      OutputImg0(12)=>OutputImg0_12, OutputImg0(11)=>OutputImg0_11, 
      OutputImg0(10)=>OutputImg0_10, OutputImg0(9)=>OutputImg0_9, 
      OutputImg0(8)=>OutputImg0_8, OutputImg0(7)=>OutputImg0_7, 
      OutputImg0(6)=>OutputImg0_6, OutputImg0(5)=>OutputImg0_5, 
      OutputImg0(4)=>OutputImg0_4, OutputImg0(3)=>OutputImg0_3, 
      OutputImg0(2)=>OutputImg0_2, OutputImg0(1)=>OutputImg0_1, 
      OutputImg0(0)=>OutputImg0_0, OutputImg1(447)=>DANGLING(800), 
      OutputImg1(446)=>DANGLING(801), OutputImg1(445)=>DANGLING(802), 
      OutputImg1(444)=>DANGLING(803), OutputImg1(443)=>DANGLING(804), 
      OutputImg1(442)=>DANGLING(805), OutputImg1(441)=>DANGLING(806), 
      OutputImg1(440)=>DANGLING(807), OutputImg1(439)=>DANGLING(808), 
      OutputImg1(438)=>DANGLING(809), OutputImg1(437)=>DANGLING(810), 
      OutputImg1(436)=>DANGLING(811), OutputImg1(435)=>DANGLING(812), 
      OutputImg1(434)=>DANGLING(813), OutputImg1(433)=>DANGLING(814), 
      OutputImg1(432)=>DANGLING(815), OutputImg1(431)=>DANGLING(816), 
      OutputImg1(430)=>DANGLING(817), OutputImg1(429)=>DANGLING(818), 
      OutputImg1(428)=>DANGLING(819), OutputImg1(427)=>DANGLING(820), 
      OutputImg1(426)=>DANGLING(821), OutputImg1(425)=>DANGLING(822), 
      OutputImg1(424)=>DANGLING(823), OutputImg1(423)=>DANGLING(824), 
      OutputImg1(422)=>DANGLING(825), OutputImg1(421)=>DANGLING(826), 
      OutputImg1(420)=>DANGLING(827), OutputImg1(419)=>DANGLING(828), 
      OutputImg1(418)=>DANGLING(829), OutputImg1(417)=>DANGLING(830), 
      OutputImg1(416)=>DANGLING(831), OutputImg1(415)=>DANGLING(832), 
      OutputImg1(414)=>DANGLING(833), OutputImg1(413)=>DANGLING(834), 
      OutputImg1(412)=>DANGLING(835), OutputImg1(411)=>DANGLING(836), 
      OutputImg1(410)=>DANGLING(837), OutputImg1(409)=>DANGLING(838), 
      OutputImg1(408)=>DANGLING(839), OutputImg1(407)=>DANGLING(840), 
      OutputImg1(406)=>DANGLING(841), OutputImg1(405)=>DANGLING(842), 
      OutputImg1(404)=>DANGLING(843), OutputImg1(403)=>DANGLING(844), 
      OutputImg1(402)=>DANGLING(845), OutputImg1(401)=>DANGLING(846), 
      OutputImg1(400)=>DANGLING(847), OutputImg1(399)=>DANGLING(848), 
      OutputImg1(398)=>DANGLING(849), OutputImg1(397)=>DANGLING(850), 
      OutputImg1(396)=>DANGLING(851), OutputImg1(395)=>DANGLING(852), 
      OutputImg1(394)=>DANGLING(853), OutputImg1(393)=>DANGLING(854), 
      OutputImg1(392)=>DANGLING(855), OutputImg1(391)=>DANGLING(856), 
      OutputImg1(390)=>DANGLING(857), OutputImg1(389)=>DANGLING(858), 
      OutputImg1(388)=>DANGLING(859), OutputImg1(387)=>DANGLING(860), 
      OutputImg1(386)=>DANGLING(861), OutputImg1(385)=>DANGLING(862), 
      OutputImg1(384)=>DANGLING(863), OutputImg1(383)=>DANGLING(864), 
      OutputImg1(382)=>DANGLING(865), OutputImg1(381)=>DANGLING(866), 
      OutputImg1(380)=>DANGLING(867), OutputImg1(379)=>DANGLING(868), 
      OutputImg1(378)=>DANGLING(869), OutputImg1(377)=>DANGLING(870), 
      OutputImg1(376)=>DANGLING(871), OutputImg1(375)=>DANGLING(872), 
      OutputImg1(374)=>DANGLING(873), OutputImg1(373)=>DANGLING(874), 
      OutputImg1(372)=>DANGLING(875), OutputImg1(371)=>DANGLING(876), 
      OutputImg1(370)=>DANGLING(877), OutputImg1(369)=>DANGLING(878), 
      OutputImg1(368)=>DANGLING(879), OutputImg1(367)=>DANGLING(880), 
      OutputImg1(366)=>DANGLING(881), OutputImg1(365)=>DANGLING(882), 
      OutputImg1(364)=>DANGLING(883), OutputImg1(363)=>DANGLING(884), 
      OutputImg1(362)=>DANGLING(885), OutputImg1(361)=>DANGLING(886), 
      OutputImg1(360)=>DANGLING(887), OutputImg1(359)=>DANGLING(888), 
      OutputImg1(358)=>DANGLING(889), OutputImg1(357)=>DANGLING(890), 
      OutputImg1(356)=>DANGLING(891), OutputImg1(355)=>DANGLING(892), 
      OutputImg1(354)=>DANGLING(893), OutputImg1(353)=>DANGLING(894), 
      OutputImg1(352)=>DANGLING(895), OutputImg1(351)=>DANGLING(896), 
      OutputImg1(350)=>DANGLING(897), OutputImg1(349)=>DANGLING(898), 
      OutputImg1(348)=>DANGLING(899), OutputImg1(347)=>DANGLING(900), 
      OutputImg1(346)=>DANGLING(901), OutputImg1(345)=>DANGLING(902), 
      OutputImg1(344)=>DANGLING(903), OutputImg1(343)=>DANGLING(904), 
      OutputImg1(342)=>DANGLING(905), OutputImg1(341)=>DANGLING(906), 
      OutputImg1(340)=>DANGLING(907), OutputImg1(339)=>DANGLING(908), 
      OutputImg1(338)=>DANGLING(909), OutputImg1(337)=>DANGLING(910), 
      OutputImg1(336)=>DANGLING(911), OutputImg1(335)=>DANGLING(912), 
      OutputImg1(334)=>DANGLING(913), OutputImg1(333)=>DANGLING(914), 
      OutputImg1(332)=>DANGLING(915), OutputImg1(331)=>DANGLING(916), 
      OutputImg1(330)=>DANGLING(917), OutputImg1(329)=>DANGLING(918), 
      OutputImg1(328)=>DANGLING(919), OutputImg1(327)=>DANGLING(920), 
      OutputImg1(326)=>DANGLING(921), OutputImg1(325)=>DANGLING(922), 
      OutputImg1(324)=>DANGLING(923), OutputImg1(323)=>DANGLING(924), 
      OutputImg1(322)=>DANGLING(925), OutputImg1(321)=>DANGLING(926), 
      OutputImg1(320)=>DANGLING(927), OutputImg1(319)=>DANGLING(928), 
      OutputImg1(318)=>DANGLING(929), OutputImg1(317)=>DANGLING(930), 
      OutputImg1(316)=>DANGLING(931), OutputImg1(315)=>DANGLING(932), 
      OutputImg1(314)=>DANGLING(933), OutputImg1(313)=>DANGLING(934), 
      OutputImg1(312)=>DANGLING(935), OutputImg1(311)=>DANGLING(936), 
      OutputImg1(310)=>DANGLING(937), OutputImg1(309)=>DANGLING(938), 
      OutputImg1(308)=>DANGLING(939), OutputImg1(307)=>DANGLING(940), 
      OutputImg1(306)=>DANGLING(941), OutputImg1(305)=>DANGLING(942), 
      OutputImg1(304)=>DANGLING(943), OutputImg1(303)=>DANGLING(944), 
      OutputImg1(302)=>DANGLING(945), OutputImg1(301)=>DANGLING(946), 
      OutputImg1(300)=>DANGLING(947), OutputImg1(299)=>DANGLING(948), 
      OutputImg1(298)=>DANGLING(949), OutputImg1(297)=>DANGLING(950), 
      OutputImg1(296)=>DANGLING(951), OutputImg1(295)=>DANGLING(952), 
      OutputImg1(294)=>DANGLING(953), OutputImg1(293)=>DANGLING(954), 
      OutputImg1(292)=>DANGLING(955), OutputImg1(291)=>DANGLING(956), 
      OutputImg1(290)=>DANGLING(957), OutputImg1(289)=>DANGLING(958), 
      OutputImg1(288)=>DANGLING(959), OutputImg1(287)=>DANGLING(960), 
      OutputImg1(286)=>DANGLING(961), OutputImg1(285)=>DANGLING(962), 
      OutputImg1(284)=>DANGLING(963), OutputImg1(283)=>DANGLING(964), 
      OutputImg1(282)=>DANGLING(965), OutputImg1(281)=>DANGLING(966), 
      OutputImg1(280)=>DANGLING(967), OutputImg1(279)=>DANGLING(968), 
      OutputImg1(278)=>DANGLING(969), OutputImg1(277)=>DANGLING(970), 
      OutputImg1(276)=>DANGLING(971), OutputImg1(275)=>DANGLING(972), 
      OutputImg1(274)=>DANGLING(973), OutputImg1(273)=>DANGLING(974), 
      OutputImg1(272)=>DANGLING(975), OutputImg1(271)=>DANGLING(976), 
      OutputImg1(270)=>DANGLING(977), OutputImg1(269)=>DANGLING(978), 
      OutputImg1(268)=>DANGLING(979), OutputImg1(267)=>DANGLING(980), 
      OutputImg1(266)=>DANGLING(981), OutputImg1(265)=>DANGLING(982), 
      OutputImg1(264)=>DANGLING(983), OutputImg1(263)=>DANGLING(984), 
      OutputImg1(262)=>DANGLING(985), OutputImg1(261)=>DANGLING(986), 
      OutputImg1(260)=>DANGLING(987), OutputImg1(259)=>DANGLING(988), 
      OutputImg1(258)=>DANGLING(989), OutputImg1(257)=>DANGLING(990), 
      OutputImg1(256)=>DANGLING(991), OutputImg1(255)=>DANGLING(992), 
      OutputImg1(254)=>DANGLING(993), OutputImg1(253)=>DANGLING(994), 
      OutputImg1(252)=>DANGLING(995), OutputImg1(251)=>DANGLING(996), 
      OutputImg1(250)=>DANGLING(997), OutputImg1(249)=>DANGLING(998), 
      OutputImg1(248)=>DANGLING(999), OutputImg1(247)=>DANGLING(1000), 
      OutputImg1(246)=>DANGLING(1001), OutputImg1(245)=>DANGLING(1002), 
      OutputImg1(244)=>DANGLING(1003), OutputImg1(243)=>DANGLING(1004), 
      OutputImg1(242)=>DANGLING(1005), OutputImg1(241)=>DANGLING(1006), 
      OutputImg1(240)=>DANGLING(1007), OutputImg1(239)=>DANGLING(1008), 
      OutputImg1(238)=>DANGLING(1009), OutputImg1(237)=>DANGLING(1010), 
      OutputImg1(236)=>DANGLING(1011), OutputImg1(235)=>DANGLING(1012), 
      OutputImg1(234)=>DANGLING(1013), OutputImg1(233)=>DANGLING(1014), 
      OutputImg1(232)=>DANGLING(1015), OutputImg1(231)=>DANGLING(1016), 
      OutputImg1(230)=>DANGLING(1017), OutputImg1(229)=>DANGLING(1018), 
      OutputImg1(228)=>DANGLING(1019), OutputImg1(227)=>DANGLING(1020), 
      OutputImg1(226)=>DANGLING(1021), OutputImg1(225)=>DANGLING(1022), 
      OutputImg1(224)=>DANGLING(1023), OutputImg1(223)=>DANGLING(1024), 
      OutputImg1(222)=>DANGLING(1025), OutputImg1(221)=>DANGLING(1026), 
      OutputImg1(220)=>DANGLING(1027), OutputImg1(219)=>DANGLING(1028), 
      OutputImg1(218)=>DANGLING(1029), OutputImg1(217)=>DANGLING(1030), 
      OutputImg1(216)=>DANGLING(1031), OutputImg1(215)=>DANGLING(1032), 
      OutputImg1(214)=>DANGLING(1033), OutputImg1(213)=>DANGLING(1034), 
      OutputImg1(212)=>DANGLING(1035), OutputImg1(211)=>DANGLING(1036), 
      OutputImg1(210)=>DANGLING(1037), OutputImg1(209)=>DANGLING(1038), 
      OutputImg1(208)=>DANGLING(1039), OutputImg1(207)=>DANGLING(1040), 
      OutputImg1(206)=>DANGLING(1041), OutputImg1(205)=>DANGLING(1042), 
      OutputImg1(204)=>DANGLING(1043), OutputImg1(203)=>DANGLING(1044), 
      OutputImg1(202)=>DANGLING(1045), OutputImg1(201)=>DANGLING(1046), 
      OutputImg1(200)=>DANGLING(1047), OutputImg1(199)=>DANGLING(1048), 
      OutputImg1(198)=>DANGLING(1049), OutputImg1(197)=>DANGLING(1050), 
      OutputImg1(196)=>DANGLING(1051), OutputImg1(195)=>DANGLING(1052), 
      OutputImg1(194)=>DANGLING(1053), OutputImg1(193)=>DANGLING(1054), 
      OutputImg1(192)=>DANGLING(1055), OutputImg1(191)=>DANGLING(1056), 
      OutputImg1(190)=>DANGLING(1057), OutputImg1(189)=>DANGLING(1058), 
      OutputImg1(188)=>DANGLING(1059), OutputImg1(187)=>DANGLING(1060), 
      OutputImg1(186)=>DANGLING(1061), OutputImg1(185)=>DANGLING(1062), 
      OutputImg1(184)=>DANGLING(1063), OutputImg1(183)=>DANGLING(1064), 
      OutputImg1(182)=>DANGLING(1065), OutputImg1(181)=>DANGLING(1066), 
      OutputImg1(180)=>DANGLING(1067), OutputImg1(179)=>DANGLING(1068), 
      OutputImg1(178)=>DANGLING(1069), OutputImg1(177)=>DANGLING(1070), 
      OutputImg1(176)=>DANGLING(1071), OutputImg1(175)=>DANGLING(1072), 
      OutputImg1(174)=>DANGLING(1073), OutputImg1(173)=>DANGLING(1074), 
      OutputImg1(172)=>DANGLING(1075), OutputImg1(171)=>DANGLING(1076), 
      OutputImg1(170)=>DANGLING(1077), OutputImg1(169)=>DANGLING(1078), 
      OutputImg1(168)=>DANGLING(1079), OutputImg1(167)=>DANGLING(1080), 
      OutputImg1(166)=>DANGLING(1081), OutputImg1(165)=>DANGLING(1082), 
      OutputImg1(164)=>DANGLING(1083), OutputImg1(163)=>DANGLING(1084), 
      OutputImg1(162)=>DANGLING(1085), OutputImg1(161)=>DANGLING(1086), 
      OutputImg1(160)=>DANGLING(1087), OutputImg1(159)=>DANGLING(1088), 
      OutputImg1(158)=>DANGLING(1089), OutputImg1(157)=>DANGLING(1090), 
      OutputImg1(156)=>DANGLING(1091), OutputImg1(155)=>DANGLING(1092), 
      OutputImg1(154)=>DANGLING(1093), OutputImg1(153)=>DANGLING(1094), 
      OutputImg1(152)=>DANGLING(1095), OutputImg1(151)=>DANGLING(1096), 
      OutputImg1(150)=>DANGLING(1097), OutputImg1(149)=>DANGLING(1098), 
      OutputImg1(148)=>DANGLING(1099), OutputImg1(147)=>DANGLING(1100), 
      OutputImg1(146)=>DANGLING(1101), OutputImg1(145)=>DANGLING(1102), 
      OutputImg1(144)=>DANGLING(1103), OutputImg1(143)=>DANGLING(1104), 
      OutputImg1(142)=>DANGLING(1105), OutputImg1(141)=>DANGLING(1106), 
      OutputImg1(140)=>DANGLING(1107), OutputImg1(139)=>DANGLING(1108), 
      OutputImg1(138)=>DANGLING(1109), OutputImg1(137)=>DANGLING(1110), 
      OutputImg1(136)=>DANGLING(1111), OutputImg1(135)=>DANGLING(1112), 
      OutputImg1(134)=>DANGLING(1113), OutputImg1(133)=>DANGLING(1114), 
      OutputImg1(132)=>DANGLING(1115), OutputImg1(131)=>DANGLING(1116), 
      OutputImg1(130)=>DANGLING(1117), OutputImg1(129)=>DANGLING(1118), 
      OutputImg1(128)=>DANGLING(1119), OutputImg1(127)=>DANGLING(1120), 
      OutputImg1(126)=>DANGLING(1121), OutputImg1(125)=>DANGLING(1122), 
      OutputImg1(124)=>DANGLING(1123), OutputImg1(123)=>DANGLING(1124), 
      OutputImg1(122)=>DANGLING(1125), OutputImg1(121)=>DANGLING(1126), 
      OutputImg1(120)=>DANGLING(1127), OutputImg1(119)=>DANGLING(1128), 
      OutputImg1(118)=>DANGLING(1129), OutputImg1(117)=>DANGLING(1130), 
      OutputImg1(116)=>DANGLING(1131), OutputImg1(115)=>DANGLING(1132), 
      OutputImg1(114)=>DANGLING(1133), OutputImg1(113)=>DANGLING(1134), 
      OutputImg1(112)=>DANGLING(1135), OutputImg1(111)=>DANGLING(1136), 
      OutputImg1(110)=>DANGLING(1137), OutputImg1(109)=>DANGLING(1138), 
      OutputImg1(108)=>DANGLING(1139), OutputImg1(107)=>DANGLING(1140), 
      OutputImg1(106)=>DANGLING(1141), OutputImg1(105)=>DANGLING(1142), 
      OutputImg1(104)=>DANGLING(1143), OutputImg1(103)=>DANGLING(1144), 
      OutputImg1(102)=>DANGLING(1145), OutputImg1(101)=>DANGLING(1146), 
      OutputImg1(100)=>DANGLING(1147), OutputImg1(99)=>DANGLING(1148), 
      OutputImg1(98)=>DANGLING(1149), OutputImg1(97)=>DANGLING(1150), 
      OutputImg1(96)=>DANGLING(1151), OutputImg1(95)=>DANGLING(1152), 
      OutputImg1(94)=>DANGLING(1153), OutputImg1(93)=>DANGLING(1154), 
      OutputImg1(92)=>DANGLING(1155), OutputImg1(91)=>DANGLING(1156), 
      OutputImg1(90)=>DANGLING(1157), OutputImg1(89)=>DANGLING(1158), 
      OutputImg1(88)=>DANGLING(1159), OutputImg1(87)=>DANGLING(1160), 
      OutputImg1(86)=>DANGLING(1161), OutputImg1(85)=>DANGLING(1162), 
      OutputImg1(84)=>DANGLING(1163), OutputImg1(83)=>DANGLING(1164), 
      OutputImg1(82)=>DANGLING(1165), OutputImg1(81)=>DANGLING(1166), 
      OutputImg1(80)=>DANGLING(1167), OutputImg1(79)=>OutputImg1_79, 
      OutputImg1(78)=>OutputImg1_78, OutputImg1(77)=>OutputImg1_77, 
      OutputImg1(76)=>OutputImg1_76, OutputImg1(75)=>OutputImg1_75, 
      OutputImg1(74)=>OutputImg1_74, OutputImg1(73)=>OutputImg1_73, 
      OutputImg1(72)=>OutputImg1_72, OutputImg1(71)=>OutputImg1_71, 
      OutputImg1(70)=>OutputImg1_70, OutputImg1(69)=>OutputImg1_69, 
      OutputImg1(68)=>OutputImg1_68, OutputImg1(67)=>OutputImg1_67, 
      OutputImg1(66)=>OutputImg1_66, OutputImg1(65)=>OutputImg1_65, 
      OutputImg1(64)=>OutputImg1_64, OutputImg1(63)=>OutputImg1_63, 
      OutputImg1(62)=>OutputImg1_62, OutputImg1(61)=>OutputImg1_61, 
      OutputImg1(60)=>OutputImg1_60, OutputImg1(59)=>OutputImg1_59, 
      OutputImg1(58)=>OutputImg1_58, OutputImg1(57)=>OutputImg1_57, 
      OutputImg1(56)=>OutputImg1_56, OutputImg1(55)=>OutputImg1_55, 
      OutputImg1(54)=>OutputImg1_54, OutputImg1(53)=>OutputImg1_53, 
      OutputImg1(52)=>OutputImg1_52, OutputImg1(51)=>OutputImg1_51, 
      OutputImg1(50)=>OutputImg1_50, OutputImg1(49)=>OutputImg1_49, 
      OutputImg1(48)=>OutputImg1_48, OutputImg1(47)=>OutputImg1_47, 
      OutputImg1(46)=>OutputImg1_46, OutputImg1(45)=>OutputImg1_45, 
      OutputImg1(44)=>OutputImg1_44, OutputImg1(43)=>OutputImg1_43, 
      OutputImg1(42)=>OutputImg1_42, OutputImg1(41)=>OutputImg1_41, 
      OutputImg1(40)=>OutputImg1_40, OutputImg1(39)=>OutputImg1_39, 
      OutputImg1(38)=>OutputImg1_38, OutputImg1(37)=>OutputImg1_37, 
      OutputImg1(36)=>OutputImg1_36, OutputImg1(35)=>OutputImg1_35, 
      OutputImg1(34)=>OutputImg1_34, OutputImg1(33)=>OutputImg1_33, 
      OutputImg1(32)=>OutputImg1_32, OutputImg1(31)=>OutputImg1_31, 
      OutputImg1(30)=>OutputImg1_30, OutputImg1(29)=>OutputImg1_29, 
      OutputImg1(28)=>OutputImg1_28, OutputImg1(27)=>OutputImg1_27, 
      OutputImg1(26)=>OutputImg1_26, OutputImg1(25)=>OutputImg1_25, 
      OutputImg1(24)=>OutputImg1_24, OutputImg1(23)=>OutputImg1_23, 
      OutputImg1(22)=>OutputImg1_22, OutputImg1(21)=>OutputImg1_21, 
      OutputImg1(20)=>OutputImg1_20, OutputImg1(19)=>OutputImg1_19, 
      OutputImg1(18)=>OutputImg1_18, OutputImg1(17)=>OutputImg1_17, 
      OutputImg1(16)=>OutputImg1_16, OutputImg1(15)=>OutputImg1_15, 
      OutputImg1(14)=>OutputImg1_14, OutputImg1(13)=>OutputImg1_13, 
      OutputImg1(12)=>OutputImg1_12, OutputImg1(11)=>OutputImg1_11, 
      OutputImg1(10)=>OutputImg1_10, OutputImg1(9)=>OutputImg1_9, 
      OutputImg1(8)=>OutputImg1_8, OutputImg1(7)=>OutputImg1_7, 
      OutputImg1(6)=>OutputImg1_6, OutputImg1(5)=>OutputImg1_5, 
      OutputImg1(4)=>OutputImg1_4, OutputImg1(3)=>OutputImg1_3, 
      OutputImg1(2)=>OutputImg1_2, OutputImg1(1)=>OutputImg1_1, 
      OutputImg1(0)=>OutputImg1_0, OutputImg2(447)=>DANGLING(1168), 
      OutputImg2(446)=>DANGLING(1169), OutputImg2(445)=>DANGLING(1170), 
      OutputImg2(444)=>DANGLING(1171), OutputImg2(443)=>DANGLING(1172), 
      OutputImg2(442)=>DANGLING(1173), OutputImg2(441)=>DANGLING(1174), 
      OutputImg2(440)=>DANGLING(1175), OutputImg2(439)=>DANGLING(1176), 
      OutputImg2(438)=>DANGLING(1177), OutputImg2(437)=>DANGLING(1178), 
      OutputImg2(436)=>DANGLING(1179), OutputImg2(435)=>DANGLING(1180), 
      OutputImg2(434)=>DANGLING(1181), OutputImg2(433)=>DANGLING(1182), 
      OutputImg2(432)=>DANGLING(1183), OutputImg2(431)=>DANGLING(1184), 
      OutputImg2(430)=>DANGLING(1185), OutputImg2(429)=>DANGLING(1186), 
      OutputImg2(428)=>DANGLING(1187), OutputImg2(427)=>DANGLING(1188), 
      OutputImg2(426)=>DANGLING(1189), OutputImg2(425)=>DANGLING(1190), 
      OutputImg2(424)=>DANGLING(1191), OutputImg2(423)=>DANGLING(1192), 
      OutputImg2(422)=>DANGLING(1193), OutputImg2(421)=>DANGLING(1194), 
      OutputImg2(420)=>DANGLING(1195), OutputImg2(419)=>DANGLING(1196), 
      OutputImg2(418)=>DANGLING(1197), OutputImg2(417)=>DANGLING(1198), 
      OutputImg2(416)=>DANGLING(1199), OutputImg2(415)=>DANGLING(1200), 
      OutputImg2(414)=>DANGLING(1201), OutputImg2(413)=>DANGLING(1202), 
      OutputImg2(412)=>DANGLING(1203), OutputImg2(411)=>DANGLING(1204), 
      OutputImg2(410)=>DANGLING(1205), OutputImg2(409)=>DANGLING(1206), 
      OutputImg2(408)=>DANGLING(1207), OutputImg2(407)=>DANGLING(1208), 
      OutputImg2(406)=>DANGLING(1209), OutputImg2(405)=>DANGLING(1210), 
      OutputImg2(404)=>DANGLING(1211), OutputImg2(403)=>DANGLING(1212), 
      OutputImg2(402)=>DANGLING(1213), OutputImg2(401)=>DANGLING(1214), 
      OutputImg2(400)=>DANGLING(1215), OutputImg2(399)=>DANGLING(1216), 
      OutputImg2(398)=>DANGLING(1217), OutputImg2(397)=>DANGLING(1218), 
      OutputImg2(396)=>DANGLING(1219), OutputImg2(395)=>DANGLING(1220), 
      OutputImg2(394)=>DANGLING(1221), OutputImg2(393)=>DANGLING(1222), 
      OutputImg2(392)=>DANGLING(1223), OutputImg2(391)=>DANGLING(1224), 
      OutputImg2(390)=>DANGLING(1225), OutputImg2(389)=>DANGLING(1226), 
      OutputImg2(388)=>DANGLING(1227), OutputImg2(387)=>DANGLING(1228), 
      OutputImg2(386)=>DANGLING(1229), OutputImg2(385)=>DANGLING(1230), 
      OutputImg2(384)=>DANGLING(1231), OutputImg2(383)=>DANGLING(1232), 
      OutputImg2(382)=>DANGLING(1233), OutputImg2(381)=>DANGLING(1234), 
      OutputImg2(380)=>DANGLING(1235), OutputImg2(379)=>DANGLING(1236), 
      OutputImg2(378)=>DANGLING(1237), OutputImg2(377)=>DANGLING(1238), 
      OutputImg2(376)=>DANGLING(1239), OutputImg2(375)=>DANGLING(1240), 
      OutputImg2(374)=>DANGLING(1241), OutputImg2(373)=>DANGLING(1242), 
      OutputImg2(372)=>DANGLING(1243), OutputImg2(371)=>DANGLING(1244), 
      OutputImg2(370)=>DANGLING(1245), OutputImg2(369)=>DANGLING(1246), 
      OutputImg2(368)=>DANGLING(1247), OutputImg2(367)=>DANGLING(1248), 
      OutputImg2(366)=>DANGLING(1249), OutputImg2(365)=>DANGLING(1250), 
      OutputImg2(364)=>DANGLING(1251), OutputImg2(363)=>DANGLING(1252), 
      OutputImg2(362)=>DANGLING(1253), OutputImg2(361)=>DANGLING(1254), 
      OutputImg2(360)=>DANGLING(1255), OutputImg2(359)=>DANGLING(1256), 
      OutputImg2(358)=>DANGLING(1257), OutputImg2(357)=>DANGLING(1258), 
      OutputImg2(356)=>DANGLING(1259), OutputImg2(355)=>DANGLING(1260), 
      OutputImg2(354)=>DANGLING(1261), OutputImg2(353)=>DANGLING(1262), 
      OutputImg2(352)=>DANGLING(1263), OutputImg2(351)=>DANGLING(1264), 
      OutputImg2(350)=>DANGLING(1265), OutputImg2(349)=>DANGLING(1266), 
      OutputImg2(348)=>DANGLING(1267), OutputImg2(347)=>DANGLING(1268), 
      OutputImg2(346)=>DANGLING(1269), OutputImg2(345)=>DANGLING(1270), 
      OutputImg2(344)=>DANGLING(1271), OutputImg2(343)=>DANGLING(1272), 
      OutputImg2(342)=>DANGLING(1273), OutputImg2(341)=>DANGLING(1274), 
      OutputImg2(340)=>DANGLING(1275), OutputImg2(339)=>DANGLING(1276), 
      OutputImg2(338)=>DANGLING(1277), OutputImg2(337)=>DANGLING(1278), 
      OutputImg2(336)=>DANGLING(1279), OutputImg2(335)=>DANGLING(1280), 
      OutputImg2(334)=>DANGLING(1281), OutputImg2(333)=>DANGLING(1282), 
      OutputImg2(332)=>DANGLING(1283), OutputImg2(331)=>DANGLING(1284), 
      OutputImg2(330)=>DANGLING(1285), OutputImg2(329)=>DANGLING(1286), 
      OutputImg2(328)=>DANGLING(1287), OutputImg2(327)=>DANGLING(1288), 
      OutputImg2(326)=>DANGLING(1289), OutputImg2(325)=>DANGLING(1290), 
      OutputImg2(324)=>DANGLING(1291), OutputImg2(323)=>DANGLING(1292), 
      OutputImg2(322)=>DANGLING(1293), OutputImg2(321)=>DANGLING(1294), 
      OutputImg2(320)=>DANGLING(1295), OutputImg2(319)=>DANGLING(1296), 
      OutputImg2(318)=>DANGLING(1297), OutputImg2(317)=>DANGLING(1298), 
      OutputImg2(316)=>DANGLING(1299), OutputImg2(315)=>DANGLING(1300), 
      OutputImg2(314)=>DANGLING(1301), OutputImg2(313)=>DANGLING(1302), 
      OutputImg2(312)=>DANGLING(1303), OutputImg2(311)=>DANGLING(1304), 
      OutputImg2(310)=>DANGLING(1305), OutputImg2(309)=>DANGLING(1306), 
      OutputImg2(308)=>DANGLING(1307), OutputImg2(307)=>DANGLING(1308), 
      OutputImg2(306)=>DANGLING(1309), OutputImg2(305)=>DANGLING(1310), 
      OutputImg2(304)=>DANGLING(1311), OutputImg2(303)=>DANGLING(1312), 
      OutputImg2(302)=>DANGLING(1313), OutputImg2(301)=>DANGLING(1314), 
      OutputImg2(300)=>DANGLING(1315), OutputImg2(299)=>DANGLING(1316), 
      OutputImg2(298)=>DANGLING(1317), OutputImg2(297)=>DANGLING(1318), 
      OutputImg2(296)=>DANGLING(1319), OutputImg2(295)=>DANGLING(1320), 
      OutputImg2(294)=>DANGLING(1321), OutputImg2(293)=>DANGLING(1322), 
      OutputImg2(292)=>DANGLING(1323), OutputImg2(291)=>DANGLING(1324), 
      OutputImg2(290)=>DANGLING(1325), OutputImg2(289)=>DANGLING(1326), 
      OutputImg2(288)=>DANGLING(1327), OutputImg2(287)=>DANGLING(1328), 
      OutputImg2(286)=>DANGLING(1329), OutputImg2(285)=>DANGLING(1330), 
      OutputImg2(284)=>DANGLING(1331), OutputImg2(283)=>DANGLING(1332), 
      OutputImg2(282)=>DANGLING(1333), OutputImg2(281)=>DANGLING(1334), 
      OutputImg2(280)=>DANGLING(1335), OutputImg2(279)=>DANGLING(1336), 
      OutputImg2(278)=>DANGLING(1337), OutputImg2(277)=>DANGLING(1338), 
      OutputImg2(276)=>DANGLING(1339), OutputImg2(275)=>DANGLING(1340), 
      OutputImg2(274)=>DANGLING(1341), OutputImg2(273)=>DANGLING(1342), 
      OutputImg2(272)=>DANGLING(1343), OutputImg2(271)=>DANGLING(1344), 
      OutputImg2(270)=>DANGLING(1345), OutputImg2(269)=>DANGLING(1346), 
      OutputImg2(268)=>DANGLING(1347), OutputImg2(267)=>DANGLING(1348), 
      OutputImg2(266)=>DANGLING(1349), OutputImg2(265)=>DANGLING(1350), 
      OutputImg2(264)=>DANGLING(1351), OutputImg2(263)=>DANGLING(1352), 
      OutputImg2(262)=>DANGLING(1353), OutputImg2(261)=>DANGLING(1354), 
      OutputImg2(260)=>DANGLING(1355), OutputImg2(259)=>DANGLING(1356), 
      OutputImg2(258)=>DANGLING(1357), OutputImg2(257)=>DANGLING(1358), 
      OutputImg2(256)=>DANGLING(1359), OutputImg2(255)=>DANGLING(1360), 
      OutputImg2(254)=>DANGLING(1361), OutputImg2(253)=>DANGLING(1362), 
      OutputImg2(252)=>DANGLING(1363), OutputImg2(251)=>DANGLING(1364), 
      OutputImg2(250)=>DANGLING(1365), OutputImg2(249)=>DANGLING(1366), 
      OutputImg2(248)=>DANGLING(1367), OutputImg2(247)=>DANGLING(1368), 
      OutputImg2(246)=>DANGLING(1369), OutputImg2(245)=>DANGLING(1370), 
      OutputImg2(244)=>DANGLING(1371), OutputImg2(243)=>DANGLING(1372), 
      OutputImg2(242)=>DANGLING(1373), OutputImg2(241)=>DANGLING(1374), 
      OutputImg2(240)=>DANGLING(1375), OutputImg2(239)=>DANGLING(1376), 
      OutputImg2(238)=>DANGLING(1377), OutputImg2(237)=>DANGLING(1378), 
      OutputImg2(236)=>DANGLING(1379), OutputImg2(235)=>DANGLING(1380), 
      OutputImg2(234)=>DANGLING(1381), OutputImg2(233)=>DANGLING(1382), 
      OutputImg2(232)=>DANGLING(1383), OutputImg2(231)=>DANGLING(1384), 
      OutputImg2(230)=>DANGLING(1385), OutputImg2(229)=>DANGLING(1386), 
      OutputImg2(228)=>DANGLING(1387), OutputImg2(227)=>DANGLING(1388), 
      OutputImg2(226)=>DANGLING(1389), OutputImg2(225)=>DANGLING(1390), 
      OutputImg2(224)=>DANGLING(1391), OutputImg2(223)=>DANGLING(1392), 
      OutputImg2(222)=>DANGLING(1393), OutputImg2(221)=>DANGLING(1394), 
      OutputImg2(220)=>DANGLING(1395), OutputImg2(219)=>DANGLING(1396), 
      OutputImg2(218)=>DANGLING(1397), OutputImg2(217)=>DANGLING(1398), 
      OutputImg2(216)=>DANGLING(1399), OutputImg2(215)=>DANGLING(1400), 
      OutputImg2(214)=>DANGLING(1401), OutputImg2(213)=>DANGLING(1402), 
      OutputImg2(212)=>DANGLING(1403), OutputImg2(211)=>DANGLING(1404), 
      OutputImg2(210)=>DANGLING(1405), OutputImg2(209)=>DANGLING(1406), 
      OutputImg2(208)=>DANGLING(1407), OutputImg2(207)=>DANGLING(1408), 
      OutputImg2(206)=>DANGLING(1409), OutputImg2(205)=>DANGLING(1410), 
      OutputImg2(204)=>DANGLING(1411), OutputImg2(203)=>DANGLING(1412), 
      OutputImg2(202)=>DANGLING(1413), OutputImg2(201)=>DANGLING(1414), 
      OutputImg2(200)=>DANGLING(1415), OutputImg2(199)=>DANGLING(1416), 
      OutputImg2(198)=>DANGLING(1417), OutputImg2(197)=>DANGLING(1418), 
      OutputImg2(196)=>DANGLING(1419), OutputImg2(195)=>DANGLING(1420), 
      OutputImg2(194)=>DANGLING(1421), OutputImg2(193)=>DANGLING(1422), 
      OutputImg2(192)=>DANGLING(1423), OutputImg2(191)=>DANGLING(1424), 
      OutputImg2(190)=>DANGLING(1425), OutputImg2(189)=>DANGLING(1426), 
      OutputImg2(188)=>DANGLING(1427), OutputImg2(187)=>DANGLING(1428), 
      OutputImg2(186)=>DANGLING(1429), OutputImg2(185)=>DANGLING(1430), 
      OutputImg2(184)=>DANGLING(1431), OutputImg2(183)=>DANGLING(1432), 
      OutputImg2(182)=>DANGLING(1433), OutputImg2(181)=>DANGLING(1434), 
      OutputImg2(180)=>DANGLING(1435), OutputImg2(179)=>DANGLING(1436), 
      OutputImg2(178)=>DANGLING(1437), OutputImg2(177)=>DANGLING(1438), 
      OutputImg2(176)=>DANGLING(1439), OutputImg2(175)=>DANGLING(1440), 
      OutputImg2(174)=>DANGLING(1441), OutputImg2(173)=>DANGLING(1442), 
      OutputImg2(172)=>DANGLING(1443), OutputImg2(171)=>DANGLING(1444), 
      OutputImg2(170)=>DANGLING(1445), OutputImg2(169)=>DANGLING(1446), 
      OutputImg2(168)=>DANGLING(1447), OutputImg2(167)=>DANGLING(1448), 
      OutputImg2(166)=>DANGLING(1449), OutputImg2(165)=>DANGLING(1450), 
      OutputImg2(164)=>DANGLING(1451), OutputImg2(163)=>DANGLING(1452), 
      OutputImg2(162)=>DANGLING(1453), OutputImg2(161)=>DANGLING(1454), 
      OutputImg2(160)=>DANGLING(1455), OutputImg2(159)=>DANGLING(1456), 
      OutputImg2(158)=>DANGLING(1457), OutputImg2(157)=>DANGLING(1458), 
      OutputImg2(156)=>DANGLING(1459), OutputImg2(155)=>DANGLING(1460), 
      OutputImg2(154)=>DANGLING(1461), OutputImg2(153)=>DANGLING(1462), 
      OutputImg2(152)=>DANGLING(1463), OutputImg2(151)=>DANGLING(1464), 
      OutputImg2(150)=>DANGLING(1465), OutputImg2(149)=>DANGLING(1466), 
      OutputImg2(148)=>DANGLING(1467), OutputImg2(147)=>DANGLING(1468), 
      OutputImg2(146)=>DANGLING(1469), OutputImg2(145)=>DANGLING(1470), 
      OutputImg2(144)=>DANGLING(1471), OutputImg2(143)=>DANGLING(1472), 
      OutputImg2(142)=>DANGLING(1473), OutputImg2(141)=>DANGLING(1474), 
      OutputImg2(140)=>DANGLING(1475), OutputImg2(139)=>DANGLING(1476), 
      OutputImg2(138)=>DANGLING(1477), OutputImg2(137)=>DANGLING(1478), 
      OutputImg2(136)=>DANGLING(1479), OutputImg2(135)=>DANGLING(1480), 
      OutputImg2(134)=>DANGLING(1481), OutputImg2(133)=>DANGLING(1482), 
      OutputImg2(132)=>DANGLING(1483), OutputImg2(131)=>DANGLING(1484), 
      OutputImg2(130)=>DANGLING(1485), OutputImg2(129)=>DANGLING(1486), 
      OutputImg2(128)=>DANGLING(1487), OutputImg2(127)=>DANGLING(1488), 
      OutputImg2(126)=>DANGLING(1489), OutputImg2(125)=>DANGLING(1490), 
      OutputImg2(124)=>DANGLING(1491), OutputImg2(123)=>DANGLING(1492), 
      OutputImg2(122)=>DANGLING(1493), OutputImg2(121)=>DANGLING(1494), 
      OutputImg2(120)=>DANGLING(1495), OutputImg2(119)=>DANGLING(1496), 
      OutputImg2(118)=>DANGLING(1497), OutputImg2(117)=>DANGLING(1498), 
      OutputImg2(116)=>DANGLING(1499), OutputImg2(115)=>DANGLING(1500), 
      OutputImg2(114)=>DANGLING(1501), OutputImg2(113)=>DANGLING(1502), 
      OutputImg2(112)=>DANGLING(1503), OutputImg2(111)=>DANGLING(1504), 
      OutputImg2(110)=>DANGLING(1505), OutputImg2(109)=>DANGLING(1506), 
      OutputImg2(108)=>DANGLING(1507), OutputImg2(107)=>DANGLING(1508), 
      OutputImg2(106)=>DANGLING(1509), OutputImg2(105)=>DANGLING(1510), 
      OutputImg2(104)=>DANGLING(1511), OutputImg2(103)=>DANGLING(1512), 
      OutputImg2(102)=>DANGLING(1513), OutputImg2(101)=>DANGLING(1514), 
      OutputImg2(100)=>DANGLING(1515), OutputImg2(99)=>DANGLING(1516), 
      OutputImg2(98)=>DANGLING(1517), OutputImg2(97)=>DANGLING(1518), 
      OutputImg2(96)=>DANGLING(1519), OutputImg2(95)=>DANGLING(1520), 
      OutputImg2(94)=>DANGLING(1521), OutputImg2(93)=>DANGLING(1522), 
      OutputImg2(92)=>DANGLING(1523), OutputImg2(91)=>DANGLING(1524), 
      OutputImg2(90)=>DANGLING(1525), OutputImg2(89)=>DANGLING(1526), 
      OutputImg2(88)=>DANGLING(1527), OutputImg2(87)=>DANGLING(1528), 
      OutputImg2(86)=>DANGLING(1529), OutputImg2(85)=>DANGLING(1530), 
      OutputImg2(84)=>DANGLING(1531), OutputImg2(83)=>DANGLING(1532), 
      OutputImg2(82)=>DANGLING(1533), OutputImg2(81)=>DANGLING(1534), 
      OutputImg2(80)=>DANGLING(1535), OutputImg2(79)=>OutputImg2_79, 
      OutputImg2(78)=>OutputImg2_78, OutputImg2(77)=>OutputImg2_77, 
      OutputImg2(76)=>OutputImg2_76, OutputImg2(75)=>OutputImg2_75, 
      OutputImg2(74)=>OutputImg2_74, OutputImg2(73)=>OutputImg2_73, 
      OutputImg2(72)=>OutputImg2_72, OutputImg2(71)=>OutputImg2_71, 
      OutputImg2(70)=>OutputImg2_70, OutputImg2(69)=>OutputImg2_69, 
      OutputImg2(68)=>OutputImg2_68, OutputImg2(67)=>OutputImg2_67, 
      OutputImg2(66)=>OutputImg2_66, OutputImg2(65)=>OutputImg2_65, 
      OutputImg2(64)=>OutputImg2_64, OutputImg2(63)=>OutputImg2_63, 
      OutputImg2(62)=>OutputImg2_62, OutputImg2(61)=>OutputImg2_61, 
      OutputImg2(60)=>OutputImg2_60, OutputImg2(59)=>OutputImg2_59, 
      OutputImg2(58)=>OutputImg2_58, OutputImg2(57)=>OutputImg2_57, 
      OutputImg2(56)=>OutputImg2_56, OutputImg2(55)=>OutputImg2_55, 
      OutputImg2(54)=>OutputImg2_54, OutputImg2(53)=>OutputImg2_53, 
      OutputImg2(52)=>OutputImg2_52, OutputImg2(51)=>OutputImg2_51, 
      OutputImg2(50)=>OutputImg2_50, OutputImg2(49)=>OutputImg2_49, 
      OutputImg2(48)=>OutputImg2_48, OutputImg2(47)=>OutputImg2_47, 
      OutputImg2(46)=>OutputImg2_46, OutputImg2(45)=>OutputImg2_45, 
      OutputImg2(44)=>OutputImg2_44, OutputImg2(43)=>OutputImg2_43, 
      OutputImg2(42)=>OutputImg2_42, OutputImg2(41)=>OutputImg2_41, 
      OutputImg2(40)=>OutputImg2_40, OutputImg2(39)=>OutputImg2_39, 
      OutputImg2(38)=>OutputImg2_38, OutputImg2(37)=>OutputImg2_37, 
      OutputImg2(36)=>OutputImg2_36, OutputImg2(35)=>OutputImg2_35, 
      OutputImg2(34)=>OutputImg2_34, OutputImg2(33)=>OutputImg2_33, 
      OutputImg2(32)=>OutputImg2_32, OutputImg2(31)=>OutputImg2_31, 
      OutputImg2(30)=>OutputImg2_30, OutputImg2(29)=>OutputImg2_29, 
      OutputImg2(28)=>OutputImg2_28, OutputImg2(27)=>OutputImg2_27, 
      OutputImg2(26)=>OutputImg2_26, OutputImg2(25)=>OutputImg2_25, 
      OutputImg2(24)=>OutputImg2_24, OutputImg2(23)=>OutputImg2_23, 
      OutputImg2(22)=>OutputImg2_22, OutputImg2(21)=>OutputImg2_21, 
      OutputImg2(20)=>OutputImg2_20, OutputImg2(19)=>OutputImg2_19, 
      OutputImg2(18)=>OutputImg2_18, OutputImg2(17)=>OutputImg2_17, 
      OutputImg2(16)=>OutputImg2_16, OutputImg2(15)=>OutputImg2_15, 
      OutputImg2(14)=>OutputImg2_14, OutputImg2(13)=>OutputImg2_13, 
      OutputImg2(12)=>OutputImg2_12, OutputImg2(11)=>OutputImg2_11, 
      OutputImg2(10)=>OutputImg2_10, OutputImg2(9)=>OutputImg2_9, 
      OutputImg2(8)=>OutputImg2_8, OutputImg2(7)=>OutputImg2_7, 
      OutputImg2(6)=>OutputImg2_6, OutputImg2(5)=>OutputImg2_5, 
      OutputImg2(4)=>OutputImg2_4, OutputImg2(3)=>OutputImg2_3, 
      OutputImg2(2)=>OutputImg2_2, OutputImg2(1)=>OutputImg2_1, 
      OutputImg2(0)=>OutputImg2_0, OutputImg3(447)=>DANGLING(1536), 
      OutputImg3(446)=>DANGLING(1537), OutputImg3(445)=>DANGLING(1538), 
      OutputImg3(444)=>DANGLING(1539), OutputImg3(443)=>DANGLING(1540), 
      OutputImg3(442)=>DANGLING(1541), OutputImg3(441)=>DANGLING(1542), 
      OutputImg3(440)=>DANGLING(1543), OutputImg3(439)=>DANGLING(1544), 
      OutputImg3(438)=>DANGLING(1545), OutputImg3(437)=>DANGLING(1546), 
      OutputImg3(436)=>DANGLING(1547), OutputImg3(435)=>DANGLING(1548), 
      OutputImg3(434)=>DANGLING(1549), OutputImg3(433)=>DANGLING(1550), 
      OutputImg3(432)=>DANGLING(1551), OutputImg3(431)=>DANGLING(1552), 
      OutputImg3(430)=>DANGLING(1553), OutputImg3(429)=>DANGLING(1554), 
      OutputImg3(428)=>DANGLING(1555), OutputImg3(427)=>DANGLING(1556), 
      OutputImg3(426)=>DANGLING(1557), OutputImg3(425)=>DANGLING(1558), 
      OutputImg3(424)=>DANGLING(1559), OutputImg3(423)=>DANGLING(1560), 
      OutputImg3(422)=>DANGLING(1561), OutputImg3(421)=>DANGLING(1562), 
      OutputImg3(420)=>DANGLING(1563), OutputImg3(419)=>DANGLING(1564), 
      OutputImg3(418)=>DANGLING(1565), OutputImg3(417)=>DANGLING(1566), 
      OutputImg3(416)=>DANGLING(1567), OutputImg3(415)=>DANGLING(1568), 
      OutputImg3(414)=>DANGLING(1569), OutputImg3(413)=>DANGLING(1570), 
      OutputImg3(412)=>DANGLING(1571), OutputImg3(411)=>DANGLING(1572), 
      OutputImg3(410)=>DANGLING(1573), OutputImg3(409)=>DANGLING(1574), 
      OutputImg3(408)=>DANGLING(1575), OutputImg3(407)=>DANGLING(1576), 
      OutputImg3(406)=>DANGLING(1577), OutputImg3(405)=>DANGLING(1578), 
      OutputImg3(404)=>DANGLING(1579), OutputImg3(403)=>DANGLING(1580), 
      OutputImg3(402)=>DANGLING(1581), OutputImg3(401)=>DANGLING(1582), 
      OutputImg3(400)=>DANGLING(1583), OutputImg3(399)=>DANGLING(1584), 
      OutputImg3(398)=>DANGLING(1585), OutputImg3(397)=>DANGLING(1586), 
      OutputImg3(396)=>DANGLING(1587), OutputImg3(395)=>DANGLING(1588), 
      OutputImg3(394)=>DANGLING(1589), OutputImg3(393)=>DANGLING(1590), 
      OutputImg3(392)=>DANGLING(1591), OutputImg3(391)=>DANGLING(1592), 
      OutputImg3(390)=>DANGLING(1593), OutputImg3(389)=>DANGLING(1594), 
      OutputImg3(388)=>DANGLING(1595), OutputImg3(387)=>DANGLING(1596), 
      OutputImg3(386)=>DANGLING(1597), OutputImg3(385)=>DANGLING(1598), 
      OutputImg3(384)=>DANGLING(1599), OutputImg3(383)=>DANGLING(1600), 
      OutputImg3(382)=>DANGLING(1601), OutputImg3(381)=>DANGLING(1602), 
      OutputImg3(380)=>DANGLING(1603), OutputImg3(379)=>DANGLING(1604), 
      OutputImg3(378)=>DANGLING(1605), OutputImg3(377)=>DANGLING(1606), 
      OutputImg3(376)=>DANGLING(1607), OutputImg3(375)=>DANGLING(1608), 
      OutputImg3(374)=>DANGLING(1609), OutputImg3(373)=>DANGLING(1610), 
      OutputImg3(372)=>DANGLING(1611), OutputImg3(371)=>DANGLING(1612), 
      OutputImg3(370)=>DANGLING(1613), OutputImg3(369)=>DANGLING(1614), 
      OutputImg3(368)=>DANGLING(1615), OutputImg3(367)=>DANGLING(1616), 
      OutputImg3(366)=>DANGLING(1617), OutputImg3(365)=>DANGLING(1618), 
      OutputImg3(364)=>DANGLING(1619), OutputImg3(363)=>DANGLING(1620), 
      OutputImg3(362)=>DANGLING(1621), OutputImg3(361)=>DANGLING(1622), 
      OutputImg3(360)=>DANGLING(1623), OutputImg3(359)=>DANGLING(1624), 
      OutputImg3(358)=>DANGLING(1625), OutputImg3(357)=>DANGLING(1626), 
      OutputImg3(356)=>DANGLING(1627), OutputImg3(355)=>DANGLING(1628), 
      OutputImg3(354)=>DANGLING(1629), OutputImg3(353)=>DANGLING(1630), 
      OutputImg3(352)=>DANGLING(1631), OutputImg3(351)=>DANGLING(1632), 
      OutputImg3(350)=>DANGLING(1633), OutputImg3(349)=>DANGLING(1634), 
      OutputImg3(348)=>DANGLING(1635), OutputImg3(347)=>DANGLING(1636), 
      OutputImg3(346)=>DANGLING(1637), OutputImg3(345)=>DANGLING(1638), 
      OutputImg3(344)=>DANGLING(1639), OutputImg3(343)=>DANGLING(1640), 
      OutputImg3(342)=>DANGLING(1641), OutputImg3(341)=>DANGLING(1642), 
      OutputImg3(340)=>DANGLING(1643), OutputImg3(339)=>DANGLING(1644), 
      OutputImg3(338)=>DANGLING(1645), OutputImg3(337)=>DANGLING(1646), 
      OutputImg3(336)=>DANGLING(1647), OutputImg3(335)=>DANGLING(1648), 
      OutputImg3(334)=>DANGLING(1649), OutputImg3(333)=>DANGLING(1650), 
      OutputImg3(332)=>DANGLING(1651), OutputImg3(331)=>DANGLING(1652), 
      OutputImg3(330)=>DANGLING(1653), OutputImg3(329)=>DANGLING(1654), 
      OutputImg3(328)=>DANGLING(1655), OutputImg3(327)=>DANGLING(1656), 
      OutputImg3(326)=>DANGLING(1657), OutputImg3(325)=>DANGLING(1658), 
      OutputImg3(324)=>DANGLING(1659), OutputImg3(323)=>DANGLING(1660), 
      OutputImg3(322)=>DANGLING(1661), OutputImg3(321)=>DANGLING(1662), 
      OutputImg3(320)=>DANGLING(1663), OutputImg3(319)=>DANGLING(1664), 
      OutputImg3(318)=>DANGLING(1665), OutputImg3(317)=>DANGLING(1666), 
      OutputImg3(316)=>DANGLING(1667), OutputImg3(315)=>DANGLING(1668), 
      OutputImg3(314)=>DANGLING(1669), OutputImg3(313)=>DANGLING(1670), 
      OutputImg3(312)=>DANGLING(1671), OutputImg3(311)=>DANGLING(1672), 
      OutputImg3(310)=>DANGLING(1673), OutputImg3(309)=>DANGLING(1674), 
      OutputImg3(308)=>DANGLING(1675), OutputImg3(307)=>DANGLING(1676), 
      OutputImg3(306)=>DANGLING(1677), OutputImg3(305)=>DANGLING(1678), 
      OutputImg3(304)=>DANGLING(1679), OutputImg3(303)=>DANGLING(1680), 
      OutputImg3(302)=>DANGLING(1681), OutputImg3(301)=>DANGLING(1682), 
      OutputImg3(300)=>DANGLING(1683), OutputImg3(299)=>DANGLING(1684), 
      OutputImg3(298)=>DANGLING(1685), OutputImg3(297)=>DANGLING(1686), 
      OutputImg3(296)=>DANGLING(1687), OutputImg3(295)=>DANGLING(1688), 
      OutputImg3(294)=>DANGLING(1689), OutputImg3(293)=>DANGLING(1690), 
      OutputImg3(292)=>DANGLING(1691), OutputImg3(291)=>DANGLING(1692), 
      OutputImg3(290)=>DANGLING(1693), OutputImg3(289)=>DANGLING(1694), 
      OutputImg3(288)=>DANGLING(1695), OutputImg3(287)=>DANGLING(1696), 
      OutputImg3(286)=>DANGLING(1697), OutputImg3(285)=>DANGLING(1698), 
      OutputImg3(284)=>DANGLING(1699), OutputImg3(283)=>DANGLING(1700), 
      OutputImg3(282)=>DANGLING(1701), OutputImg3(281)=>DANGLING(1702), 
      OutputImg3(280)=>DANGLING(1703), OutputImg3(279)=>DANGLING(1704), 
      OutputImg3(278)=>DANGLING(1705), OutputImg3(277)=>DANGLING(1706), 
      OutputImg3(276)=>DANGLING(1707), OutputImg3(275)=>DANGLING(1708), 
      OutputImg3(274)=>DANGLING(1709), OutputImg3(273)=>DANGLING(1710), 
      OutputImg3(272)=>DANGLING(1711), OutputImg3(271)=>DANGLING(1712), 
      OutputImg3(270)=>DANGLING(1713), OutputImg3(269)=>DANGLING(1714), 
      OutputImg3(268)=>DANGLING(1715), OutputImg3(267)=>DANGLING(1716), 
      OutputImg3(266)=>DANGLING(1717), OutputImg3(265)=>DANGLING(1718), 
      OutputImg3(264)=>DANGLING(1719), OutputImg3(263)=>DANGLING(1720), 
      OutputImg3(262)=>DANGLING(1721), OutputImg3(261)=>DANGLING(1722), 
      OutputImg3(260)=>DANGLING(1723), OutputImg3(259)=>DANGLING(1724), 
      OutputImg3(258)=>DANGLING(1725), OutputImg3(257)=>DANGLING(1726), 
      OutputImg3(256)=>DANGLING(1727), OutputImg3(255)=>DANGLING(1728), 
      OutputImg3(254)=>DANGLING(1729), OutputImg3(253)=>DANGLING(1730), 
      OutputImg3(252)=>DANGLING(1731), OutputImg3(251)=>DANGLING(1732), 
      OutputImg3(250)=>DANGLING(1733), OutputImg3(249)=>DANGLING(1734), 
      OutputImg3(248)=>DANGLING(1735), OutputImg3(247)=>DANGLING(1736), 
      OutputImg3(246)=>DANGLING(1737), OutputImg3(245)=>DANGLING(1738), 
      OutputImg3(244)=>DANGLING(1739), OutputImg3(243)=>DANGLING(1740), 
      OutputImg3(242)=>DANGLING(1741), OutputImg3(241)=>DANGLING(1742), 
      OutputImg3(240)=>DANGLING(1743), OutputImg3(239)=>DANGLING(1744), 
      OutputImg3(238)=>DANGLING(1745), OutputImg3(237)=>DANGLING(1746), 
      OutputImg3(236)=>DANGLING(1747), OutputImg3(235)=>DANGLING(1748), 
      OutputImg3(234)=>DANGLING(1749), OutputImg3(233)=>DANGLING(1750), 
      OutputImg3(232)=>DANGLING(1751), OutputImg3(231)=>DANGLING(1752), 
      OutputImg3(230)=>DANGLING(1753), OutputImg3(229)=>DANGLING(1754), 
      OutputImg3(228)=>DANGLING(1755), OutputImg3(227)=>DANGLING(1756), 
      OutputImg3(226)=>DANGLING(1757), OutputImg3(225)=>DANGLING(1758), 
      OutputImg3(224)=>DANGLING(1759), OutputImg3(223)=>DANGLING(1760), 
      OutputImg3(222)=>DANGLING(1761), OutputImg3(221)=>DANGLING(1762), 
      OutputImg3(220)=>DANGLING(1763), OutputImg3(219)=>DANGLING(1764), 
      OutputImg3(218)=>DANGLING(1765), OutputImg3(217)=>DANGLING(1766), 
      OutputImg3(216)=>DANGLING(1767), OutputImg3(215)=>DANGLING(1768), 
      OutputImg3(214)=>DANGLING(1769), OutputImg3(213)=>DANGLING(1770), 
      OutputImg3(212)=>DANGLING(1771), OutputImg3(211)=>DANGLING(1772), 
      OutputImg3(210)=>DANGLING(1773), OutputImg3(209)=>DANGLING(1774), 
      OutputImg3(208)=>DANGLING(1775), OutputImg3(207)=>DANGLING(1776), 
      OutputImg3(206)=>DANGLING(1777), OutputImg3(205)=>DANGLING(1778), 
      OutputImg3(204)=>DANGLING(1779), OutputImg3(203)=>DANGLING(1780), 
      OutputImg3(202)=>DANGLING(1781), OutputImg3(201)=>DANGLING(1782), 
      OutputImg3(200)=>DANGLING(1783), OutputImg3(199)=>DANGLING(1784), 
      OutputImg3(198)=>DANGLING(1785), OutputImg3(197)=>DANGLING(1786), 
      OutputImg3(196)=>DANGLING(1787), OutputImg3(195)=>DANGLING(1788), 
      OutputImg3(194)=>DANGLING(1789), OutputImg3(193)=>DANGLING(1790), 
      OutputImg3(192)=>DANGLING(1791), OutputImg3(191)=>DANGLING(1792), 
      OutputImg3(190)=>DANGLING(1793), OutputImg3(189)=>DANGLING(1794), 
      OutputImg3(188)=>DANGLING(1795), OutputImg3(187)=>DANGLING(1796), 
      OutputImg3(186)=>DANGLING(1797), OutputImg3(185)=>DANGLING(1798), 
      OutputImg3(184)=>DANGLING(1799), OutputImg3(183)=>DANGLING(1800), 
      OutputImg3(182)=>DANGLING(1801), OutputImg3(181)=>DANGLING(1802), 
      OutputImg3(180)=>DANGLING(1803), OutputImg3(179)=>DANGLING(1804), 
      OutputImg3(178)=>DANGLING(1805), OutputImg3(177)=>DANGLING(1806), 
      OutputImg3(176)=>DANGLING(1807), OutputImg3(175)=>DANGLING(1808), 
      OutputImg3(174)=>DANGLING(1809), OutputImg3(173)=>DANGLING(1810), 
      OutputImg3(172)=>DANGLING(1811), OutputImg3(171)=>DANGLING(1812), 
      OutputImg3(170)=>DANGLING(1813), OutputImg3(169)=>DANGLING(1814), 
      OutputImg3(168)=>DANGLING(1815), OutputImg3(167)=>DANGLING(1816), 
      OutputImg3(166)=>DANGLING(1817), OutputImg3(165)=>DANGLING(1818), 
      OutputImg3(164)=>DANGLING(1819), OutputImg3(163)=>DANGLING(1820), 
      OutputImg3(162)=>DANGLING(1821), OutputImg3(161)=>DANGLING(1822), 
      OutputImg3(160)=>DANGLING(1823), OutputImg3(159)=>DANGLING(1824), 
      OutputImg3(158)=>DANGLING(1825), OutputImg3(157)=>DANGLING(1826), 
      OutputImg3(156)=>DANGLING(1827), OutputImg3(155)=>DANGLING(1828), 
      OutputImg3(154)=>DANGLING(1829), OutputImg3(153)=>DANGLING(1830), 
      OutputImg3(152)=>DANGLING(1831), OutputImg3(151)=>DANGLING(1832), 
      OutputImg3(150)=>DANGLING(1833), OutputImg3(149)=>DANGLING(1834), 
      OutputImg3(148)=>DANGLING(1835), OutputImg3(147)=>DANGLING(1836), 
      OutputImg3(146)=>DANGLING(1837), OutputImg3(145)=>DANGLING(1838), 
      OutputImg3(144)=>DANGLING(1839), OutputImg3(143)=>DANGLING(1840), 
      OutputImg3(142)=>DANGLING(1841), OutputImg3(141)=>DANGLING(1842), 
      OutputImg3(140)=>DANGLING(1843), OutputImg3(139)=>DANGLING(1844), 
      OutputImg3(138)=>DANGLING(1845), OutputImg3(137)=>DANGLING(1846), 
      OutputImg3(136)=>DANGLING(1847), OutputImg3(135)=>DANGLING(1848), 
      OutputImg3(134)=>DANGLING(1849), OutputImg3(133)=>DANGLING(1850), 
      OutputImg3(132)=>DANGLING(1851), OutputImg3(131)=>DANGLING(1852), 
      OutputImg3(130)=>DANGLING(1853), OutputImg3(129)=>DANGLING(1854), 
      OutputImg3(128)=>DANGLING(1855), OutputImg3(127)=>DANGLING(1856), 
      OutputImg3(126)=>DANGLING(1857), OutputImg3(125)=>DANGLING(1858), 
      OutputImg3(124)=>DANGLING(1859), OutputImg3(123)=>DANGLING(1860), 
      OutputImg3(122)=>DANGLING(1861), OutputImg3(121)=>DANGLING(1862), 
      OutputImg3(120)=>DANGLING(1863), OutputImg3(119)=>DANGLING(1864), 
      OutputImg3(118)=>DANGLING(1865), OutputImg3(117)=>DANGLING(1866), 
      OutputImg3(116)=>DANGLING(1867), OutputImg3(115)=>DANGLING(1868), 
      OutputImg3(114)=>DANGLING(1869), OutputImg3(113)=>DANGLING(1870), 
      OutputImg3(112)=>DANGLING(1871), OutputImg3(111)=>DANGLING(1872), 
      OutputImg3(110)=>DANGLING(1873), OutputImg3(109)=>DANGLING(1874), 
      OutputImg3(108)=>DANGLING(1875), OutputImg3(107)=>DANGLING(1876), 
      OutputImg3(106)=>DANGLING(1877), OutputImg3(105)=>DANGLING(1878), 
      OutputImg3(104)=>DANGLING(1879), OutputImg3(103)=>DANGLING(1880), 
      OutputImg3(102)=>DANGLING(1881), OutputImg3(101)=>DANGLING(1882), 
      OutputImg3(100)=>DANGLING(1883), OutputImg3(99)=>DANGLING(1884), 
      OutputImg3(98)=>DANGLING(1885), OutputImg3(97)=>DANGLING(1886), 
      OutputImg3(96)=>DANGLING(1887), OutputImg3(95)=>DANGLING(1888), 
      OutputImg3(94)=>DANGLING(1889), OutputImg3(93)=>DANGLING(1890), 
      OutputImg3(92)=>DANGLING(1891), OutputImg3(91)=>DANGLING(1892), 
      OutputImg3(90)=>DANGLING(1893), OutputImg3(89)=>DANGLING(1894), 
      OutputImg3(88)=>DANGLING(1895), OutputImg3(87)=>DANGLING(1896), 
      OutputImg3(86)=>DANGLING(1897), OutputImg3(85)=>DANGLING(1898), 
      OutputImg3(84)=>DANGLING(1899), OutputImg3(83)=>DANGLING(1900), 
      OutputImg3(82)=>DANGLING(1901), OutputImg3(81)=>DANGLING(1902), 
      OutputImg3(80)=>DANGLING(1903), OutputImg3(79)=>OutputImg3_79, 
      OutputImg3(78)=>OutputImg3_78, OutputImg3(77)=>OutputImg3_77, 
      OutputImg3(76)=>OutputImg3_76, OutputImg3(75)=>OutputImg3_75, 
      OutputImg3(74)=>OutputImg3_74, OutputImg3(73)=>OutputImg3_73, 
      OutputImg3(72)=>OutputImg3_72, OutputImg3(71)=>OutputImg3_71, 
      OutputImg3(70)=>OutputImg3_70, OutputImg3(69)=>OutputImg3_69, 
      OutputImg3(68)=>OutputImg3_68, OutputImg3(67)=>OutputImg3_67, 
      OutputImg3(66)=>OutputImg3_66, OutputImg3(65)=>OutputImg3_65, 
      OutputImg3(64)=>OutputImg3_64, OutputImg3(63)=>OutputImg3_63, 
      OutputImg3(62)=>OutputImg3_62, OutputImg3(61)=>OutputImg3_61, 
      OutputImg3(60)=>OutputImg3_60, OutputImg3(59)=>OutputImg3_59, 
      OutputImg3(58)=>OutputImg3_58, OutputImg3(57)=>OutputImg3_57, 
      OutputImg3(56)=>OutputImg3_56, OutputImg3(55)=>OutputImg3_55, 
      OutputImg3(54)=>OutputImg3_54, OutputImg3(53)=>OutputImg3_53, 
      OutputImg3(52)=>OutputImg3_52, OutputImg3(51)=>OutputImg3_51, 
      OutputImg3(50)=>OutputImg3_50, OutputImg3(49)=>OutputImg3_49, 
      OutputImg3(48)=>OutputImg3_48, OutputImg3(47)=>OutputImg3_47, 
      OutputImg3(46)=>OutputImg3_46, OutputImg3(45)=>OutputImg3_45, 
      OutputImg3(44)=>OutputImg3_44, OutputImg3(43)=>OutputImg3_43, 
      OutputImg3(42)=>OutputImg3_42, OutputImg3(41)=>OutputImg3_41, 
      OutputImg3(40)=>OutputImg3_40, OutputImg3(39)=>OutputImg3_39, 
      OutputImg3(38)=>OutputImg3_38, OutputImg3(37)=>OutputImg3_37, 
      OutputImg3(36)=>OutputImg3_36, OutputImg3(35)=>OutputImg3_35, 
      OutputImg3(34)=>OutputImg3_34, OutputImg3(33)=>OutputImg3_33, 
      OutputImg3(32)=>OutputImg3_32, OutputImg3(31)=>OutputImg3_31, 
      OutputImg3(30)=>OutputImg3_30, OutputImg3(29)=>OutputImg3_29, 
      OutputImg3(28)=>OutputImg3_28, OutputImg3(27)=>OutputImg3_27, 
      OutputImg3(26)=>OutputImg3_26, OutputImg3(25)=>OutputImg3_25, 
      OutputImg3(24)=>OutputImg3_24, OutputImg3(23)=>OutputImg3_23, 
      OutputImg3(22)=>OutputImg3_22, OutputImg3(21)=>OutputImg3_21, 
      OutputImg3(20)=>OutputImg3_20, OutputImg3(19)=>OutputImg3_19, 
      OutputImg3(18)=>OutputImg3_18, OutputImg3(17)=>OutputImg3_17, 
      OutputImg3(16)=>OutputImg3_16, OutputImg3(15)=>OutputImg3_15, 
      OutputImg3(14)=>OutputImg3_14, OutputImg3(13)=>OutputImg3_13, 
      OutputImg3(12)=>OutputImg3_12, OutputImg3(11)=>OutputImg3_11, 
      OutputImg3(10)=>OutputImg3_10, OutputImg3(9)=>OutputImg3_9, 
      OutputImg3(8)=>OutputImg3_8, OutputImg3(7)=>OutputImg3_7, 
      OutputImg3(6)=>OutputImg3_6, OutputImg3(5)=>OutputImg3_5, 
      OutputImg3(4)=>OutputImg3_4, OutputImg3(3)=>OutputImg3_3, 
      OutputImg3(2)=>OutputImg3_2, OutputImg3(1)=>OutputImg3_1, 
      OutputImg3(0)=>OutputImg3_0, OutputImg4(447)=>DANGLING(1904), 
      OutputImg4(446)=>DANGLING(1905), OutputImg4(445)=>DANGLING(1906), 
      OutputImg4(444)=>DANGLING(1907), OutputImg4(443)=>DANGLING(1908), 
      OutputImg4(442)=>DANGLING(1909), OutputImg4(441)=>DANGLING(1910), 
      OutputImg4(440)=>DANGLING(1911), OutputImg4(439)=>DANGLING(1912), 
      OutputImg4(438)=>DANGLING(1913), OutputImg4(437)=>DANGLING(1914), 
      OutputImg4(436)=>DANGLING(1915), OutputImg4(435)=>DANGLING(1916), 
      OutputImg4(434)=>DANGLING(1917), OutputImg4(433)=>DANGLING(1918), 
      OutputImg4(432)=>DANGLING(1919), OutputImg4(431)=>DANGLING(1920), 
      OutputImg4(430)=>DANGLING(1921), OutputImg4(429)=>DANGLING(1922), 
      OutputImg4(428)=>DANGLING(1923), OutputImg4(427)=>DANGLING(1924), 
      OutputImg4(426)=>DANGLING(1925), OutputImg4(425)=>DANGLING(1926), 
      OutputImg4(424)=>DANGLING(1927), OutputImg4(423)=>DANGLING(1928), 
      OutputImg4(422)=>DANGLING(1929), OutputImg4(421)=>DANGLING(1930), 
      OutputImg4(420)=>DANGLING(1931), OutputImg4(419)=>DANGLING(1932), 
      OutputImg4(418)=>DANGLING(1933), OutputImg4(417)=>DANGLING(1934), 
      OutputImg4(416)=>DANGLING(1935), OutputImg4(415)=>DANGLING(1936), 
      OutputImg4(414)=>DANGLING(1937), OutputImg4(413)=>DANGLING(1938), 
      OutputImg4(412)=>DANGLING(1939), OutputImg4(411)=>DANGLING(1940), 
      OutputImg4(410)=>DANGLING(1941), OutputImg4(409)=>DANGLING(1942), 
      OutputImg4(408)=>DANGLING(1943), OutputImg4(407)=>DANGLING(1944), 
      OutputImg4(406)=>DANGLING(1945), OutputImg4(405)=>DANGLING(1946), 
      OutputImg4(404)=>DANGLING(1947), OutputImg4(403)=>DANGLING(1948), 
      OutputImg4(402)=>DANGLING(1949), OutputImg4(401)=>DANGLING(1950), 
      OutputImg4(400)=>DANGLING(1951), OutputImg4(399)=>DANGLING(1952), 
      OutputImg4(398)=>DANGLING(1953), OutputImg4(397)=>DANGLING(1954), 
      OutputImg4(396)=>DANGLING(1955), OutputImg4(395)=>DANGLING(1956), 
      OutputImg4(394)=>DANGLING(1957), OutputImg4(393)=>DANGLING(1958), 
      OutputImg4(392)=>DANGLING(1959), OutputImg4(391)=>DANGLING(1960), 
      OutputImg4(390)=>DANGLING(1961), OutputImg4(389)=>DANGLING(1962), 
      OutputImg4(388)=>DANGLING(1963), OutputImg4(387)=>DANGLING(1964), 
      OutputImg4(386)=>DANGLING(1965), OutputImg4(385)=>DANGLING(1966), 
      OutputImg4(384)=>DANGLING(1967), OutputImg4(383)=>DANGLING(1968), 
      OutputImg4(382)=>DANGLING(1969), OutputImg4(381)=>DANGLING(1970), 
      OutputImg4(380)=>DANGLING(1971), OutputImg4(379)=>DANGLING(1972), 
      OutputImg4(378)=>DANGLING(1973), OutputImg4(377)=>DANGLING(1974), 
      OutputImg4(376)=>DANGLING(1975), OutputImg4(375)=>DANGLING(1976), 
      OutputImg4(374)=>DANGLING(1977), OutputImg4(373)=>DANGLING(1978), 
      OutputImg4(372)=>DANGLING(1979), OutputImg4(371)=>DANGLING(1980), 
      OutputImg4(370)=>DANGLING(1981), OutputImg4(369)=>DANGLING(1982), 
      OutputImg4(368)=>DANGLING(1983), OutputImg4(367)=>DANGLING(1984), 
      OutputImg4(366)=>DANGLING(1985), OutputImg4(365)=>DANGLING(1986), 
      OutputImg4(364)=>DANGLING(1987), OutputImg4(363)=>DANGLING(1988), 
      OutputImg4(362)=>DANGLING(1989), OutputImg4(361)=>DANGLING(1990), 
      OutputImg4(360)=>DANGLING(1991), OutputImg4(359)=>DANGLING(1992), 
      OutputImg4(358)=>DANGLING(1993), OutputImg4(357)=>DANGLING(1994), 
      OutputImg4(356)=>DANGLING(1995), OutputImg4(355)=>DANGLING(1996), 
      OutputImg4(354)=>DANGLING(1997), OutputImg4(353)=>DANGLING(1998), 
      OutputImg4(352)=>DANGLING(1999), OutputImg4(351)=>DANGLING(2000), 
      OutputImg4(350)=>DANGLING(2001), OutputImg4(349)=>DANGLING(2002), 
      OutputImg4(348)=>DANGLING(2003), OutputImg4(347)=>DANGLING(2004), 
      OutputImg4(346)=>DANGLING(2005), OutputImg4(345)=>DANGLING(2006), 
      OutputImg4(344)=>DANGLING(2007), OutputImg4(343)=>DANGLING(2008), 
      OutputImg4(342)=>DANGLING(2009), OutputImg4(341)=>DANGLING(2010), 
      OutputImg4(340)=>DANGLING(2011), OutputImg4(339)=>DANGLING(2012), 
      OutputImg4(338)=>DANGLING(2013), OutputImg4(337)=>DANGLING(2014), 
      OutputImg4(336)=>DANGLING(2015), OutputImg4(335)=>DANGLING(2016), 
      OutputImg4(334)=>DANGLING(2017), OutputImg4(333)=>DANGLING(2018), 
      OutputImg4(332)=>DANGLING(2019), OutputImg4(331)=>DANGLING(2020), 
      OutputImg4(330)=>DANGLING(2021), OutputImg4(329)=>DANGLING(2022), 
      OutputImg4(328)=>DANGLING(2023), OutputImg4(327)=>DANGLING(2024), 
      OutputImg4(326)=>DANGLING(2025), OutputImg4(325)=>DANGLING(2026), 
      OutputImg4(324)=>DANGLING(2027), OutputImg4(323)=>DANGLING(2028), 
      OutputImg4(322)=>DANGLING(2029), OutputImg4(321)=>DANGLING(2030), 
      OutputImg4(320)=>DANGLING(2031), OutputImg4(319)=>DANGLING(2032), 
      OutputImg4(318)=>DANGLING(2033), OutputImg4(317)=>DANGLING(2034), 
      OutputImg4(316)=>DANGLING(2035), OutputImg4(315)=>DANGLING(2036), 
      OutputImg4(314)=>DANGLING(2037), OutputImg4(313)=>DANGLING(2038), 
      OutputImg4(312)=>DANGLING(2039), OutputImg4(311)=>DANGLING(2040), 
      OutputImg4(310)=>DANGLING(2041), OutputImg4(309)=>DANGLING(2042), 
      OutputImg4(308)=>DANGLING(2043), OutputImg4(307)=>DANGLING(2044), 
      OutputImg4(306)=>DANGLING(2045), OutputImg4(305)=>DANGLING(2046), 
      OutputImg4(304)=>DANGLING(2047), OutputImg4(303)=>DANGLING(2048), 
      OutputImg4(302)=>DANGLING(2049), OutputImg4(301)=>DANGLING(2050), 
      OutputImg4(300)=>DANGLING(2051), OutputImg4(299)=>DANGLING(2052), 
      OutputImg4(298)=>DANGLING(2053), OutputImg4(297)=>DANGLING(2054), 
      OutputImg4(296)=>DANGLING(2055), OutputImg4(295)=>DANGLING(2056), 
      OutputImg4(294)=>DANGLING(2057), OutputImg4(293)=>DANGLING(2058), 
      OutputImg4(292)=>DANGLING(2059), OutputImg4(291)=>DANGLING(2060), 
      OutputImg4(290)=>DANGLING(2061), OutputImg4(289)=>DANGLING(2062), 
      OutputImg4(288)=>DANGLING(2063), OutputImg4(287)=>DANGLING(2064), 
      OutputImg4(286)=>DANGLING(2065), OutputImg4(285)=>DANGLING(2066), 
      OutputImg4(284)=>DANGLING(2067), OutputImg4(283)=>DANGLING(2068), 
      OutputImg4(282)=>DANGLING(2069), OutputImg4(281)=>DANGLING(2070), 
      OutputImg4(280)=>DANGLING(2071), OutputImg4(279)=>DANGLING(2072), 
      OutputImg4(278)=>DANGLING(2073), OutputImg4(277)=>DANGLING(2074), 
      OutputImg4(276)=>DANGLING(2075), OutputImg4(275)=>DANGLING(2076), 
      OutputImg4(274)=>DANGLING(2077), OutputImg4(273)=>DANGLING(2078), 
      OutputImg4(272)=>DANGLING(2079), OutputImg4(271)=>DANGLING(2080), 
      OutputImg4(270)=>DANGLING(2081), OutputImg4(269)=>DANGLING(2082), 
      OutputImg4(268)=>DANGLING(2083), OutputImg4(267)=>DANGLING(2084), 
      OutputImg4(266)=>DANGLING(2085), OutputImg4(265)=>DANGLING(2086), 
      OutputImg4(264)=>DANGLING(2087), OutputImg4(263)=>DANGLING(2088), 
      OutputImg4(262)=>DANGLING(2089), OutputImg4(261)=>DANGLING(2090), 
      OutputImg4(260)=>DANGLING(2091), OutputImg4(259)=>DANGLING(2092), 
      OutputImg4(258)=>DANGLING(2093), OutputImg4(257)=>DANGLING(2094), 
      OutputImg4(256)=>DANGLING(2095), OutputImg4(255)=>DANGLING(2096), 
      OutputImg4(254)=>DANGLING(2097), OutputImg4(253)=>DANGLING(2098), 
      OutputImg4(252)=>DANGLING(2099), OutputImg4(251)=>DANGLING(2100), 
      OutputImg4(250)=>DANGLING(2101), OutputImg4(249)=>DANGLING(2102), 
      OutputImg4(248)=>DANGLING(2103), OutputImg4(247)=>DANGLING(2104), 
      OutputImg4(246)=>DANGLING(2105), OutputImg4(245)=>DANGLING(2106), 
      OutputImg4(244)=>DANGLING(2107), OutputImg4(243)=>DANGLING(2108), 
      OutputImg4(242)=>DANGLING(2109), OutputImg4(241)=>DANGLING(2110), 
      OutputImg4(240)=>DANGLING(2111), OutputImg4(239)=>DANGLING(2112), 
      OutputImg4(238)=>DANGLING(2113), OutputImg4(237)=>DANGLING(2114), 
      OutputImg4(236)=>DANGLING(2115), OutputImg4(235)=>DANGLING(2116), 
      OutputImg4(234)=>DANGLING(2117), OutputImg4(233)=>DANGLING(2118), 
      OutputImg4(232)=>DANGLING(2119), OutputImg4(231)=>DANGLING(2120), 
      OutputImg4(230)=>DANGLING(2121), OutputImg4(229)=>DANGLING(2122), 
      OutputImg4(228)=>DANGLING(2123), OutputImg4(227)=>DANGLING(2124), 
      OutputImg4(226)=>DANGLING(2125), OutputImg4(225)=>DANGLING(2126), 
      OutputImg4(224)=>DANGLING(2127), OutputImg4(223)=>DANGLING(2128), 
      OutputImg4(222)=>DANGLING(2129), OutputImg4(221)=>DANGLING(2130), 
      OutputImg4(220)=>DANGLING(2131), OutputImg4(219)=>DANGLING(2132), 
      OutputImg4(218)=>DANGLING(2133), OutputImg4(217)=>DANGLING(2134), 
      OutputImg4(216)=>DANGLING(2135), OutputImg4(215)=>DANGLING(2136), 
      OutputImg4(214)=>DANGLING(2137), OutputImg4(213)=>DANGLING(2138), 
      OutputImg4(212)=>DANGLING(2139), OutputImg4(211)=>DANGLING(2140), 
      OutputImg4(210)=>DANGLING(2141), OutputImg4(209)=>DANGLING(2142), 
      OutputImg4(208)=>DANGLING(2143), OutputImg4(207)=>DANGLING(2144), 
      OutputImg4(206)=>DANGLING(2145), OutputImg4(205)=>DANGLING(2146), 
      OutputImg4(204)=>DANGLING(2147), OutputImg4(203)=>DANGLING(2148), 
      OutputImg4(202)=>DANGLING(2149), OutputImg4(201)=>DANGLING(2150), 
      OutputImg4(200)=>DANGLING(2151), OutputImg4(199)=>DANGLING(2152), 
      OutputImg4(198)=>DANGLING(2153), OutputImg4(197)=>DANGLING(2154), 
      OutputImg4(196)=>DANGLING(2155), OutputImg4(195)=>DANGLING(2156), 
      OutputImg4(194)=>DANGLING(2157), OutputImg4(193)=>DANGLING(2158), 
      OutputImg4(192)=>DANGLING(2159), OutputImg4(191)=>DANGLING(2160), 
      OutputImg4(190)=>DANGLING(2161), OutputImg4(189)=>DANGLING(2162), 
      OutputImg4(188)=>DANGLING(2163), OutputImg4(187)=>DANGLING(2164), 
      OutputImg4(186)=>DANGLING(2165), OutputImg4(185)=>DANGLING(2166), 
      OutputImg4(184)=>DANGLING(2167), OutputImg4(183)=>DANGLING(2168), 
      OutputImg4(182)=>DANGLING(2169), OutputImg4(181)=>DANGLING(2170), 
      OutputImg4(180)=>DANGLING(2171), OutputImg4(179)=>DANGLING(2172), 
      OutputImg4(178)=>DANGLING(2173), OutputImg4(177)=>DANGLING(2174), 
      OutputImg4(176)=>DANGLING(2175), OutputImg4(175)=>DANGLING(2176), 
      OutputImg4(174)=>DANGLING(2177), OutputImg4(173)=>DANGLING(2178), 
      OutputImg4(172)=>DANGLING(2179), OutputImg4(171)=>DANGLING(2180), 
      OutputImg4(170)=>DANGLING(2181), OutputImg4(169)=>DANGLING(2182), 
      OutputImg4(168)=>DANGLING(2183), OutputImg4(167)=>DANGLING(2184), 
      OutputImg4(166)=>DANGLING(2185), OutputImg4(165)=>DANGLING(2186), 
      OutputImg4(164)=>DANGLING(2187), OutputImg4(163)=>DANGLING(2188), 
      OutputImg4(162)=>DANGLING(2189), OutputImg4(161)=>DANGLING(2190), 
      OutputImg4(160)=>DANGLING(2191), OutputImg4(159)=>DANGLING(2192), 
      OutputImg4(158)=>DANGLING(2193), OutputImg4(157)=>DANGLING(2194), 
      OutputImg4(156)=>DANGLING(2195), OutputImg4(155)=>DANGLING(2196), 
      OutputImg4(154)=>DANGLING(2197), OutputImg4(153)=>DANGLING(2198), 
      OutputImg4(152)=>DANGLING(2199), OutputImg4(151)=>DANGLING(2200), 
      OutputImg4(150)=>DANGLING(2201), OutputImg4(149)=>DANGLING(2202), 
      OutputImg4(148)=>DANGLING(2203), OutputImg4(147)=>DANGLING(2204), 
      OutputImg4(146)=>DANGLING(2205), OutputImg4(145)=>DANGLING(2206), 
      OutputImg4(144)=>DANGLING(2207), OutputImg4(143)=>DANGLING(2208), 
      OutputImg4(142)=>DANGLING(2209), OutputImg4(141)=>DANGLING(2210), 
      OutputImg4(140)=>DANGLING(2211), OutputImg4(139)=>DANGLING(2212), 
      OutputImg4(138)=>DANGLING(2213), OutputImg4(137)=>DANGLING(2214), 
      OutputImg4(136)=>DANGLING(2215), OutputImg4(135)=>DANGLING(2216), 
      OutputImg4(134)=>DANGLING(2217), OutputImg4(133)=>DANGLING(2218), 
      OutputImg4(132)=>DANGLING(2219), OutputImg4(131)=>DANGLING(2220), 
      OutputImg4(130)=>DANGLING(2221), OutputImg4(129)=>DANGLING(2222), 
      OutputImg4(128)=>DANGLING(2223), OutputImg4(127)=>DANGLING(2224), 
      OutputImg4(126)=>DANGLING(2225), OutputImg4(125)=>DANGLING(2226), 
      OutputImg4(124)=>DANGLING(2227), OutputImg4(123)=>DANGLING(2228), 
      OutputImg4(122)=>DANGLING(2229), OutputImg4(121)=>DANGLING(2230), 
      OutputImg4(120)=>DANGLING(2231), OutputImg4(119)=>DANGLING(2232), 
      OutputImg4(118)=>DANGLING(2233), OutputImg4(117)=>DANGLING(2234), 
      OutputImg4(116)=>DANGLING(2235), OutputImg4(115)=>DANGLING(2236), 
      OutputImg4(114)=>DANGLING(2237), OutputImg4(113)=>DANGLING(2238), 
      OutputImg4(112)=>DANGLING(2239), OutputImg4(111)=>DANGLING(2240), 
      OutputImg4(110)=>DANGLING(2241), OutputImg4(109)=>DANGLING(2242), 
      OutputImg4(108)=>DANGLING(2243), OutputImg4(107)=>DANGLING(2244), 
      OutputImg4(106)=>DANGLING(2245), OutputImg4(105)=>DANGLING(2246), 
      OutputImg4(104)=>DANGLING(2247), OutputImg4(103)=>DANGLING(2248), 
      OutputImg4(102)=>DANGLING(2249), OutputImg4(101)=>DANGLING(2250), 
      OutputImg4(100)=>DANGLING(2251), OutputImg4(99)=>DANGLING(2252), 
      OutputImg4(98)=>DANGLING(2253), OutputImg4(97)=>DANGLING(2254), 
      OutputImg4(96)=>DANGLING(2255), OutputImg4(95)=>DANGLING(2256), 
      OutputImg4(94)=>DANGLING(2257), OutputImg4(93)=>DANGLING(2258), 
      OutputImg4(92)=>DANGLING(2259), OutputImg4(91)=>DANGLING(2260), 
      OutputImg4(90)=>DANGLING(2261), OutputImg4(89)=>DANGLING(2262), 
      OutputImg4(88)=>DANGLING(2263), OutputImg4(87)=>DANGLING(2264), 
      OutputImg4(86)=>DANGLING(2265), OutputImg4(85)=>DANGLING(2266), 
      OutputImg4(84)=>DANGLING(2267), OutputImg4(83)=>DANGLING(2268), 
      OutputImg4(82)=>DANGLING(2269), OutputImg4(81)=>DANGLING(2270), 
      OutputImg4(80)=>DANGLING(2271), OutputImg4(79)=>OutputImg4_79, 
      OutputImg4(78)=>OutputImg4_78, OutputImg4(77)=>OutputImg4_77, 
      OutputImg4(76)=>OutputImg4_76, OutputImg4(75)=>OutputImg4_75, 
      OutputImg4(74)=>OutputImg4_74, OutputImg4(73)=>OutputImg4_73, 
      OutputImg4(72)=>OutputImg4_72, OutputImg4(71)=>OutputImg4_71, 
      OutputImg4(70)=>OutputImg4_70, OutputImg4(69)=>OutputImg4_69, 
      OutputImg4(68)=>OutputImg4_68, OutputImg4(67)=>OutputImg4_67, 
      OutputImg4(66)=>OutputImg4_66, OutputImg4(65)=>OutputImg4_65, 
      OutputImg4(64)=>OutputImg4_64, OutputImg4(63)=>OutputImg4_63, 
      OutputImg4(62)=>OutputImg4_62, OutputImg4(61)=>OutputImg4_61, 
      OutputImg4(60)=>OutputImg4_60, OutputImg4(59)=>OutputImg4_59, 
      OutputImg4(58)=>OutputImg4_58, OutputImg4(57)=>OutputImg4_57, 
      OutputImg4(56)=>OutputImg4_56, OutputImg4(55)=>OutputImg4_55, 
      OutputImg4(54)=>OutputImg4_54, OutputImg4(53)=>OutputImg4_53, 
      OutputImg4(52)=>OutputImg4_52, OutputImg4(51)=>OutputImg4_51, 
      OutputImg4(50)=>OutputImg4_50, OutputImg4(49)=>OutputImg4_49, 
      OutputImg4(48)=>OutputImg4_48, OutputImg4(47)=>OutputImg4_47, 
      OutputImg4(46)=>OutputImg4_46, OutputImg4(45)=>OutputImg4_45, 
      OutputImg4(44)=>OutputImg4_44, OutputImg4(43)=>OutputImg4_43, 
      OutputImg4(42)=>OutputImg4_42, OutputImg4(41)=>OutputImg4_41, 
      OutputImg4(40)=>OutputImg4_40, OutputImg4(39)=>OutputImg4_39, 
      OutputImg4(38)=>OutputImg4_38, OutputImg4(37)=>OutputImg4_37, 
      OutputImg4(36)=>OutputImg4_36, OutputImg4(35)=>OutputImg4_35, 
      OutputImg4(34)=>OutputImg4_34, OutputImg4(33)=>OutputImg4_33, 
      OutputImg4(32)=>OutputImg4_32, OutputImg4(31)=>OutputImg4_31, 
      OutputImg4(30)=>OutputImg4_30, OutputImg4(29)=>OutputImg4_29, 
      OutputImg4(28)=>OutputImg4_28, OutputImg4(27)=>OutputImg4_27, 
      OutputImg4(26)=>OutputImg4_26, OutputImg4(25)=>OutputImg4_25, 
      OutputImg4(24)=>OutputImg4_24, OutputImg4(23)=>OutputImg4_23, 
      OutputImg4(22)=>OutputImg4_22, OutputImg4(21)=>OutputImg4_21, 
      OutputImg4(20)=>OutputImg4_20, OutputImg4(19)=>OutputImg4_19, 
      OutputImg4(18)=>OutputImg4_18, OutputImg4(17)=>OutputImg4_17, 
      OutputImg4(16)=>OutputImg4_16, OutputImg4(15)=>OutputImg4_15, 
      OutputImg4(14)=>OutputImg4_14, OutputImg4(13)=>OutputImg4_13, 
      OutputImg4(12)=>OutputImg4_12, OutputImg4(11)=>OutputImg4_11, 
      OutputImg4(10)=>OutputImg4_10, OutputImg4(9)=>OutputImg4_9, 
      OutputImg4(8)=>OutputImg4_8, OutputImg4(7)=>OutputImg4_7, 
      OutputImg4(6)=>OutputImg4_6, OutputImg4(5)=>OutputImg4_5, 
      OutputImg4(4)=>OutputImg4_4, OutputImg4(3)=>OutputImg4_3, 
      OutputImg4(2)=>OutputImg4_2, OutputImg4(1)=>OutputImg4_1, 
      OutputImg4(0)=>OutputImg4_0, OutputImg5(447)=>DANGLING(2272), 
      OutputImg5(446)=>DANGLING(2273), OutputImg5(445)=>DANGLING(2274), 
      OutputImg5(444)=>DANGLING(2275), OutputImg5(443)=>DANGLING(2276), 
      OutputImg5(442)=>DANGLING(2277), OutputImg5(441)=>DANGLING(2278), 
      OutputImg5(440)=>DANGLING(2279), OutputImg5(439)=>DANGLING(2280), 
      OutputImg5(438)=>DANGLING(2281), OutputImg5(437)=>DANGLING(2282), 
      OutputImg5(436)=>DANGLING(2283), OutputImg5(435)=>DANGLING(2284), 
      OutputImg5(434)=>DANGLING(2285), OutputImg5(433)=>DANGLING(2286), 
      OutputImg5(432)=>DANGLING(2287), OutputImg5(431)=>DANGLING(2288), 
      OutputImg5(430)=>DANGLING(2289), OutputImg5(429)=>DANGLING(2290), 
      OutputImg5(428)=>DANGLING(2291), OutputImg5(427)=>DANGLING(2292), 
      OutputImg5(426)=>DANGLING(2293), OutputImg5(425)=>DANGLING(2294), 
      OutputImg5(424)=>DANGLING(2295), OutputImg5(423)=>DANGLING(2296), 
      OutputImg5(422)=>DANGLING(2297), OutputImg5(421)=>DANGLING(2298), 
      OutputImg5(420)=>DANGLING(2299), OutputImg5(419)=>DANGLING(2300), 
      OutputImg5(418)=>DANGLING(2301), OutputImg5(417)=>DANGLING(2302), 
      OutputImg5(416)=>DANGLING(2303), OutputImg5(415)=>DANGLING(2304), 
      OutputImg5(414)=>DANGLING(2305), OutputImg5(413)=>DANGLING(2306), 
      OutputImg5(412)=>DANGLING(2307), OutputImg5(411)=>DANGLING(2308), 
      OutputImg5(410)=>DANGLING(2309), OutputImg5(409)=>DANGLING(2310), 
      OutputImg5(408)=>DANGLING(2311), OutputImg5(407)=>DANGLING(2312), 
      OutputImg5(406)=>DANGLING(2313), OutputImg5(405)=>DANGLING(2314), 
      OutputImg5(404)=>DANGLING(2315), OutputImg5(403)=>DANGLING(2316), 
      OutputImg5(402)=>DANGLING(2317), OutputImg5(401)=>DANGLING(2318), 
      OutputImg5(400)=>DANGLING(2319), OutputImg5(399)=>DANGLING(2320), 
      OutputImg5(398)=>DANGLING(2321), OutputImg5(397)=>DANGLING(2322), 
      OutputImg5(396)=>DANGLING(2323), OutputImg5(395)=>DANGLING(2324), 
      OutputImg5(394)=>DANGLING(2325), OutputImg5(393)=>DANGLING(2326), 
      OutputImg5(392)=>DANGLING(2327), OutputImg5(391)=>DANGLING(2328), 
      OutputImg5(390)=>DANGLING(2329), OutputImg5(389)=>DANGLING(2330), 
      OutputImg5(388)=>DANGLING(2331), OutputImg5(387)=>DANGLING(2332), 
      OutputImg5(386)=>DANGLING(2333), OutputImg5(385)=>DANGLING(2334), 
      OutputImg5(384)=>DANGLING(2335), OutputImg5(383)=>DANGLING(2336), 
      OutputImg5(382)=>DANGLING(2337), OutputImg5(381)=>DANGLING(2338), 
      OutputImg5(380)=>DANGLING(2339), OutputImg5(379)=>DANGLING(2340), 
      OutputImg5(378)=>DANGLING(2341), OutputImg5(377)=>DANGLING(2342), 
      OutputImg5(376)=>DANGLING(2343), OutputImg5(375)=>DANGLING(2344), 
      OutputImg5(374)=>DANGLING(2345), OutputImg5(373)=>DANGLING(2346), 
      OutputImg5(372)=>DANGLING(2347), OutputImg5(371)=>DANGLING(2348), 
      OutputImg5(370)=>DANGLING(2349), OutputImg5(369)=>DANGLING(2350), 
      OutputImg5(368)=>DANGLING(2351), OutputImg5(367)=>DANGLING(2352), 
      OutputImg5(366)=>DANGLING(2353), OutputImg5(365)=>DANGLING(2354), 
      OutputImg5(364)=>DANGLING(2355), OutputImg5(363)=>DANGLING(2356), 
      OutputImg5(362)=>DANGLING(2357), OutputImg5(361)=>DANGLING(2358), 
      OutputImg5(360)=>DANGLING(2359), OutputImg5(359)=>DANGLING(2360), 
      OutputImg5(358)=>DANGLING(2361), OutputImg5(357)=>DANGLING(2362), 
      OutputImg5(356)=>DANGLING(2363), OutputImg5(355)=>DANGLING(2364), 
      OutputImg5(354)=>DANGLING(2365), OutputImg5(353)=>DANGLING(2366), 
      OutputImg5(352)=>DANGLING(2367), OutputImg5(351)=>DANGLING(2368), 
      OutputImg5(350)=>DANGLING(2369), OutputImg5(349)=>DANGLING(2370), 
      OutputImg5(348)=>DANGLING(2371), OutputImg5(347)=>DANGLING(2372), 
      OutputImg5(346)=>DANGLING(2373), OutputImg5(345)=>DANGLING(2374), 
      OutputImg5(344)=>DANGLING(2375), OutputImg5(343)=>DANGLING(2376), 
      OutputImg5(342)=>DANGLING(2377), OutputImg5(341)=>DANGLING(2378), 
      OutputImg5(340)=>DANGLING(2379), OutputImg5(339)=>DANGLING(2380), 
      OutputImg5(338)=>DANGLING(2381), OutputImg5(337)=>DANGLING(2382), 
      OutputImg5(336)=>DANGLING(2383), OutputImg5(335)=>DANGLING(2384), 
      OutputImg5(334)=>DANGLING(2385), OutputImg5(333)=>DANGLING(2386), 
      OutputImg5(332)=>DANGLING(2387), OutputImg5(331)=>DANGLING(2388), 
      OutputImg5(330)=>DANGLING(2389), OutputImg5(329)=>DANGLING(2390), 
      OutputImg5(328)=>DANGLING(2391), OutputImg5(327)=>DANGLING(2392), 
      OutputImg5(326)=>DANGLING(2393), OutputImg5(325)=>DANGLING(2394), 
      OutputImg5(324)=>DANGLING(2395), OutputImg5(323)=>DANGLING(2396), 
      OutputImg5(322)=>DANGLING(2397), OutputImg5(321)=>DANGLING(2398), 
      OutputImg5(320)=>DANGLING(2399), OutputImg5(319)=>DANGLING(2400), 
      OutputImg5(318)=>DANGLING(2401), OutputImg5(317)=>DANGLING(2402), 
      OutputImg5(316)=>DANGLING(2403), OutputImg5(315)=>DANGLING(2404), 
      OutputImg5(314)=>DANGLING(2405), OutputImg5(313)=>DANGLING(2406), 
      OutputImg5(312)=>DANGLING(2407), OutputImg5(311)=>DANGLING(2408), 
      OutputImg5(310)=>DANGLING(2409), OutputImg5(309)=>DANGLING(2410), 
      OutputImg5(308)=>DANGLING(2411), OutputImg5(307)=>DANGLING(2412), 
      OutputImg5(306)=>DANGLING(2413), OutputImg5(305)=>DANGLING(2414), 
      OutputImg5(304)=>DANGLING(2415), OutputImg5(303)=>DANGLING(2416), 
      OutputImg5(302)=>DANGLING(2417), OutputImg5(301)=>DANGLING(2418), 
      OutputImg5(300)=>DANGLING(2419), OutputImg5(299)=>DANGLING(2420), 
      OutputImg5(298)=>DANGLING(2421), OutputImg5(297)=>DANGLING(2422), 
      OutputImg5(296)=>DANGLING(2423), OutputImg5(295)=>DANGLING(2424), 
      OutputImg5(294)=>DANGLING(2425), OutputImg5(293)=>DANGLING(2426), 
      OutputImg5(292)=>DANGLING(2427), OutputImg5(291)=>DANGLING(2428), 
      OutputImg5(290)=>DANGLING(2429), OutputImg5(289)=>DANGLING(2430), 
      OutputImg5(288)=>DANGLING(2431), OutputImg5(287)=>DANGLING(2432), 
      OutputImg5(286)=>DANGLING(2433), OutputImg5(285)=>DANGLING(2434), 
      OutputImg5(284)=>DANGLING(2435), OutputImg5(283)=>DANGLING(2436), 
      OutputImg5(282)=>DANGLING(2437), OutputImg5(281)=>DANGLING(2438), 
      OutputImg5(280)=>DANGLING(2439), OutputImg5(279)=>DANGLING(2440), 
      OutputImg5(278)=>DANGLING(2441), OutputImg5(277)=>DANGLING(2442), 
      OutputImg5(276)=>DANGLING(2443), OutputImg5(275)=>DANGLING(2444), 
      OutputImg5(274)=>DANGLING(2445), OutputImg5(273)=>DANGLING(2446), 
      OutputImg5(272)=>DANGLING(2447), OutputImg5(271)=>DANGLING(2448), 
      OutputImg5(270)=>DANGLING(2449), OutputImg5(269)=>DANGLING(2450), 
      OutputImg5(268)=>DANGLING(2451), OutputImg5(267)=>DANGLING(2452), 
      OutputImg5(266)=>DANGLING(2453), OutputImg5(265)=>DANGLING(2454), 
      OutputImg5(264)=>DANGLING(2455), OutputImg5(263)=>DANGLING(2456), 
      OutputImg5(262)=>DANGLING(2457), OutputImg5(261)=>DANGLING(2458), 
      OutputImg5(260)=>DANGLING(2459), OutputImg5(259)=>DANGLING(2460), 
      OutputImg5(258)=>DANGLING(2461), OutputImg5(257)=>DANGLING(2462), 
      OutputImg5(256)=>DANGLING(2463), OutputImg5(255)=>DANGLING(2464), 
      OutputImg5(254)=>DANGLING(2465), OutputImg5(253)=>DANGLING(2466), 
      OutputImg5(252)=>DANGLING(2467), OutputImg5(251)=>DANGLING(2468), 
      OutputImg5(250)=>DANGLING(2469), OutputImg5(249)=>DANGLING(2470), 
      OutputImg5(248)=>DANGLING(2471), OutputImg5(247)=>DANGLING(2472), 
      OutputImg5(246)=>DANGLING(2473), OutputImg5(245)=>DANGLING(2474), 
      OutputImg5(244)=>DANGLING(2475), OutputImg5(243)=>DANGLING(2476), 
      OutputImg5(242)=>DANGLING(2477), OutputImg5(241)=>DANGLING(2478), 
      OutputImg5(240)=>DANGLING(2479), OutputImg5(239)=>DANGLING(2480), 
      OutputImg5(238)=>DANGLING(2481), OutputImg5(237)=>DANGLING(2482), 
      OutputImg5(236)=>DANGLING(2483), OutputImg5(235)=>DANGLING(2484), 
      OutputImg5(234)=>DANGLING(2485), OutputImg5(233)=>DANGLING(2486), 
      OutputImg5(232)=>DANGLING(2487), OutputImg5(231)=>DANGLING(2488), 
      OutputImg5(230)=>DANGLING(2489), OutputImg5(229)=>DANGLING(2490), 
      OutputImg5(228)=>DANGLING(2491), OutputImg5(227)=>DANGLING(2492), 
      OutputImg5(226)=>DANGLING(2493), OutputImg5(225)=>DANGLING(2494), 
      OutputImg5(224)=>DANGLING(2495), OutputImg5(223)=>DANGLING(2496), 
      OutputImg5(222)=>DANGLING(2497), OutputImg5(221)=>DANGLING(2498), 
      OutputImg5(220)=>DANGLING(2499), OutputImg5(219)=>DANGLING(2500), 
      OutputImg5(218)=>DANGLING(2501), OutputImg5(217)=>DANGLING(2502), 
      OutputImg5(216)=>DANGLING(2503), OutputImg5(215)=>DANGLING(2504), 
      OutputImg5(214)=>DANGLING(2505), OutputImg5(213)=>DANGLING(2506), 
      OutputImg5(212)=>DANGLING(2507), OutputImg5(211)=>DANGLING(2508), 
      OutputImg5(210)=>DANGLING(2509), OutputImg5(209)=>DANGLING(2510), 
      OutputImg5(208)=>DANGLING(2511), OutputImg5(207)=>DANGLING(2512), 
      OutputImg5(206)=>DANGLING(2513), OutputImg5(205)=>DANGLING(2514), 
      OutputImg5(204)=>DANGLING(2515), OutputImg5(203)=>DANGLING(2516), 
      OutputImg5(202)=>DANGLING(2517), OutputImg5(201)=>DANGLING(2518), 
      OutputImg5(200)=>DANGLING(2519), OutputImg5(199)=>DANGLING(2520), 
      OutputImg5(198)=>DANGLING(2521), OutputImg5(197)=>DANGLING(2522), 
      OutputImg5(196)=>DANGLING(2523), OutputImg5(195)=>DANGLING(2524), 
      OutputImg5(194)=>DANGLING(2525), OutputImg5(193)=>DANGLING(2526), 
      OutputImg5(192)=>DANGLING(2527), OutputImg5(191)=>DANGLING(2528), 
      OutputImg5(190)=>DANGLING(2529), OutputImg5(189)=>DANGLING(2530), 
      OutputImg5(188)=>DANGLING(2531), OutputImg5(187)=>DANGLING(2532), 
      OutputImg5(186)=>DANGLING(2533), OutputImg5(185)=>DANGLING(2534), 
      OutputImg5(184)=>DANGLING(2535), OutputImg5(183)=>DANGLING(2536), 
      OutputImg5(182)=>DANGLING(2537), OutputImg5(181)=>DANGLING(2538), 
      OutputImg5(180)=>DANGLING(2539), OutputImg5(179)=>DANGLING(2540), 
      OutputImg5(178)=>DANGLING(2541), OutputImg5(177)=>DANGLING(2542), 
      OutputImg5(176)=>DANGLING(2543), OutputImg5(175)=>DANGLING(2544), 
      OutputImg5(174)=>DANGLING(2545), OutputImg5(173)=>DANGLING(2546), 
      OutputImg5(172)=>DANGLING(2547), OutputImg5(171)=>DANGLING(2548), 
      OutputImg5(170)=>DANGLING(2549), OutputImg5(169)=>DANGLING(2550), 
      OutputImg5(168)=>DANGLING(2551), OutputImg5(167)=>DANGLING(2552), 
      OutputImg5(166)=>DANGLING(2553), OutputImg5(165)=>DANGLING(2554), 
      OutputImg5(164)=>DANGLING(2555), OutputImg5(163)=>DANGLING(2556), 
      OutputImg5(162)=>DANGLING(2557), OutputImg5(161)=>DANGLING(2558), 
      OutputImg5(160)=>DANGLING(2559), OutputImg5(159)=>DANGLING(2560), 
      OutputImg5(158)=>DANGLING(2561), OutputImg5(157)=>DANGLING(2562), 
      OutputImg5(156)=>DANGLING(2563), OutputImg5(155)=>DANGLING(2564), 
      OutputImg5(154)=>DANGLING(2565), OutputImg5(153)=>DANGLING(2566), 
      OutputImg5(152)=>DANGLING(2567), OutputImg5(151)=>DANGLING(2568), 
      OutputImg5(150)=>DANGLING(2569), OutputImg5(149)=>DANGLING(2570), 
      OutputImg5(148)=>DANGLING(2571), OutputImg5(147)=>DANGLING(2572), 
      OutputImg5(146)=>DANGLING(2573), OutputImg5(145)=>DANGLING(2574), 
      OutputImg5(144)=>DANGLING(2575), OutputImg5(143)=>DANGLING(2576), 
      OutputImg5(142)=>DANGLING(2577), OutputImg5(141)=>DANGLING(2578), 
      OutputImg5(140)=>DANGLING(2579), OutputImg5(139)=>DANGLING(2580), 
      OutputImg5(138)=>DANGLING(2581), OutputImg5(137)=>DANGLING(2582), 
      OutputImg5(136)=>DANGLING(2583), OutputImg5(135)=>DANGLING(2584), 
      OutputImg5(134)=>DANGLING(2585), OutputImg5(133)=>DANGLING(2586), 
      OutputImg5(132)=>DANGLING(2587), OutputImg5(131)=>DANGLING(2588), 
      OutputImg5(130)=>DANGLING(2589), OutputImg5(129)=>DANGLING(2590), 
      OutputImg5(128)=>DANGLING(2591), OutputImg5(127)=>DANGLING(2592), 
      OutputImg5(126)=>DANGLING(2593), OutputImg5(125)=>DANGLING(2594), 
      OutputImg5(124)=>DANGLING(2595), OutputImg5(123)=>DANGLING(2596), 
      OutputImg5(122)=>DANGLING(2597), OutputImg5(121)=>DANGLING(2598), 
      OutputImg5(120)=>DANGLING(2599), OutputImg5(119)=>DANGLING(2600), 
      OutputImg5(118)=>DANGLING(2601), OutputImg5(117)=>DANGLING(2602), 
      OutputImg5(116)=>DANGLING(2603), OutputImg5(115)=>DANGLING(2604), 
      OutputImg5(114)=>DANGLING(2605), OutputImg5(113)=>DANGLING(2606), 
      OutputImg5(112)=>DANGLING(2607), OutputImg5(111)=>DANGLING(2608), 
      OutputImg5(110)=>DANGLING(2609), OutputImg5(109)=>DANGLING(2610), 
      OutputImg5(108)=>DANGLING(2611), OutputImg5(107)=>DANGLING(2612), 
      OutputImg5(106)=>DANGLING(2613), OutputImg5(105)=>DANGLING(2614), 
      OutputImg5(104)=>DANGLING(2615), OutputImg5(103)=>DANGLING(2616), 
      OutputImg5(102)=>DANGLING(2617), OutputImg5(101)=>DANGLING(2618), 
      OutputImg5(100)=>DANGLING(2619), OutputImg5(99)=>DANGLING(2620), 
      OutputImg5(98)=>DANGLING(2621), OutputImg5(97)=>DANGLING(2622), 
      OutputImg5(96)=>DANGLING(2623), OutputImg5(95)=>DANGLING(2624), 
      OutputImg5(94)=>DANGLING(2625), OutputImg5(93)=>DANGLING(2626), 
      OutputImg5(92)=>DANGLING(2627), OutputImg5(91)=>DANGLING(2628), 
      OutputImg5(90)=>DANGLING(2629), OutputImg5(89)=>DANGLING(2630), 
      OutputImg5(88)=>DANGLING(2631), OutputImg5(87)=>DANGLING(2632), 
      OutputImg5(86)=>DANGLING(2633), OutputImg5(85)=>DANGLING(2634), 
      OutputImg5(84)=>DANGLING(2635), OutputImg5(83)=>DANGLING(2636), 
      OutputImg5(82)=>DANGLING(2637), OutputImg5(81)=>DANGLING(2638), 
      OutputImg5(80)=>DANGLING(2639), OutputImg5(79)=>DANGLING(2640), 
      OutputImg5(78)=>DANGLING(2641), OutputImg5(77)=>DANGLING(2642), 
      OutputImg5(76)=>DANGLING(2643), OutputImg5(75)=>DANGLING(2644), 
      OutputImg5(74)=>DANGLING(2645), OutputImg5(73)=>DANGLING(2646), 
      OutputImg5(72)=>DANGLING(2647), OutputImg5(71)=>DANGLING(2648), 
      OutputImg5(70)=>DANGLING(2649), OutputImg5(69)=>DANGLING(2650), 
      OutputImg5(68)=>DANGLING(2651), OutputImg5(67)=>DANGLING(2652), 
      OutputImg5(66)=>DANGLING(2653), OutputImg5(65)=>DANGLING(2654), 
      OutputImg5(64)=>DANGLING(2655), OutputImg5(63)=>DANGLING(2656), 
      OutputImg5(62)=>DANGLING(2657), OutputImg5(61)=>DANGLING(2658), 
      OutputImg5(60)=>DANGLING(2659), OutputImg5(59)=>DANGLING(2660), 
      OutputImg5(58)=>DANGLING(2661), OutputImg5(57)=>DANGLING(2662), 
      OutputImg5(56)=>DANGLING(2663), OutputImg5(55)=>DANGLING(2664), 
      OutputImg5(54)=>DANGLING(2665), OutputImg5(53)=>DANGLING(2666), 
      OutputImg5(52)=>DANGLING(2667), OutputImg5(51)=>DANGLING(2668), 
      OutputImg5(50)=>DANGLING(2669), OutputImg5(49)=>DANGLING(2670), 
      OutputImg5(48)=>DANGLING(2671), OutputImg5(47)=>DANGLING(2672), 
      OutputImg5(46)=>DANGLING(2673), OutputImg5(45)=>DANGLING(2674), 
      OutputImg5(44)=>DANGLING(2675), OutputImg5(43)=>DANGLING(2676), 
      OutputImg5(42)=>DANGLING(2677), OutputImg5(41)=>DANGLING(2678), 
      OutputImg5(40)=>DANGLING(2679), OutputImg5(39)=>DANGLING(2680), 
      OutputImg5(38)=>DANGLING(2681), OutputImg5(37)=>DANGLING(2682), 
      OutputImg5(36)=>DANGLING(2683), OutputImg5(35)=>DANGLING(2684), 
      OutputImg5(34)=>DANGLING(2685), OutputImg5(33)=>DANGLING(2686), 
      OutputImg5(32)=>DANGLING(2687), OutputImg5(31)=>DANGLING(2688), 
      OutputImg5(30)=>DANGLING(2689), OutputImg5(29)=>DANGLING(2690), 
      OutputImg5(28)=>DANGLING(2691), OutputImg5(27)=>DANGLING(2692), 
      OutputImg5(26)=>DANGLING(2693), OutputImg5(25)=>DANGLING(2694), 
      OutputImg5(24)=>DANGLING(2695), OutputImg5(23)=>DANGLING(2696), 
      OutputImg5(22)=>DANGLING(2697), OutputImg5(21)=>DANGLING(2698), 
      OutputImg5(20)=>DANGLING(2699), OutputImg5(19)=>DANGLING(2700), 
      OutputImg5(18)=>DANGLING(2701), OutputImg5(17)=>DANGLING(2702), 
      OutputImg5(16)=>DANGLING(2703), OutputImg5(15)=>DANGLING(2704), 
      OutputImg5(14)=>DANGLING(2705), OutputImg5(13)=>DANGLING(2706), 
      OutputImg5(12)=>DANGLING(2707), OutputImg5(11)=>DANGLING(2708), 
      OutputImg5(10)=>DANGLING(2709), OutputImg5(9)=>DANGLING(2710), 
      OutputImg5(8)=>DANGLING(2711), OutputImg5(7)=>DANGLING(2712), 
      OutputImg5(6)=>DANGLING(2713), OutputImg5(5)=>DANGLING(2714), 
      OutputImg5(4)=>DANGLING(2715), OutputImg5(3)=>DANGLING(2716), 
      OutputImg5(2)=>DANGLING(2717), OutputImg5(1)=>DANGLING(2718), 
      OutputImg5(0)=>DANGLING(2719), ImgCounterOuput(2)=>ImgCounterOuput_2, 
      ImgCounterOuput(1)=>ImgCounterOuput_1, ImgCounterOuput(0)=>
      ImgCounterOuput_0, ImgAddToDma(12)=>AddressI_12, ImgAddToDma(11)=>
      AddressI_11, ImgAddToDma(10)=>AddressI_10, ImgAddToDma(9)=>AddressI_9, 
      ImgAddToDma(8)=>AddressI_8, ImgAddToDma(7)=>AddressI_7, ImgAddToDma(6)
      =>AddressI_6, ImgAddToDma(5)=>AddressI_5, ImgAddToDma(4)=>AddressI_4, 
      ImgAddToDma(3)=>AddressI_3, ImgAddToDma(2)=>AddressI_2, ImgAddToDma(1)
      =>AddressI_1, ImgAddToDma(0)=>AddressI_0, UpdatedAddress(12)=>
      ImgAddRegIN_12, UpdatedAddress(11)=>ImgAddRegIN_11, UpdatedAddress(10)
      =>ImgAddRegIN_10, UpdatedAddress(9)=>ImgAddRegIN_9, UpdatedAddress(8)
      =>ImgAddRegIN_8, UpdatedAddress(7)=>ImgAddRegIN_7, UpdatedAddress(6)=>
      ImgAddRegIN_6, UpdatedAddress(5)=>ImgAddRegIN_5, UpdatedAddress(4)=>
      ImgAddRegIN_4, UpdatedAddress(3)=>ImgAddRegIN_3, UpdatedAddress(2)=>
      ImgAddRegIN_2, UpdatedAddress(1)=>ImgAddRegIN_1, UpdatedAddress(0)=>
      ImgAddRegIN_0, ImgIndic(0)=>IndicatorI_0, ImgEn(5)=>DANGLING(2720), 
      ImgEn(4)=>DANGLING(2721), ImgEn(3)=>DANGLING(2722), ImgEn(2)=>DANGLING
      (2723), ImgEn(1)=>DANGLING(2724), ImgEn(0)=>DANGLING(2725), dontTrust
      =>DontRstIndicator);
   Sconv : Convolution port map ( current_state(14)=>zero_11, 
      current_state(13)=>zero_11, current_state(12)=>zero_11, 
      current_state(11)=>zero_11, current_state(10)=>zero_11, 
      current_state(9)=>zero_11, current_state(8)=>zero_11, current_state(7)
      =>nx9962, current_state(6)=>zero_11, current_state(5)=>zero_11, 
      current_state(4)=>zero_11, current_state(3)=>zero_11, current_state(2)
      =>zero_11, current_state(1)=>zero_11, current_state(0)=>zero_11, CLK=>
      nx10424, RST=>rst, QImgStat=>Q, ACK=>DANGLING(2726), LayerInfo(15)=>
      LayerInfoOut_15, LayerInfo(14)=>nx10500, LayerInfo(13)=>zero_11, 
      LayerInfo(12)=>zero_11, LayerInfo(11)=>zero_11, LayerInfo(10)=>zero_11, 
      LayerInfo(9)=>zero_11, LayerInfo(8)=>zero_11, LayerInfo(7)=>zero_11, 
      LayerInfo(6)=>zero_11, LayerInfo(5)=>zero_11, LayerInfo(4)=>zero_11, 
      LayerInfo(3)=>zero_11, LayerInfo(2)=>zero_11, LayerInfo(1)=>zero_11, 
      LayerInfo(0)=>zero_11, ImgAddress(12)=>zero_11, ImgAddress(11)=>
      zero_11, ImgAddress(10)=>zero_11, ImgAddress(9)=>zero_11, 
      ImgAddress(8)=>zero_11, ImgAddress(7)=>zero_11, ImgAddress(6)=>zero_11, 
      ImgAddress(5)=>zero_11, ImgAddress(4)=>zero_11, ImgAddress(3)=>zero_11, 
      ImgAddress(2)=>zero_11, ImgAddress(1)=>zero_11, ImgAddress(0)=>zero_11, 
      OutputImg0(79)=>OutputImg0_79, OutputImg0(78)=>OutputImg0_78, 
      OutputImg0(77)=>OutputImg0_77, OutputImg0(76)=>OutputImg0_76, 
      OutputImg0(75)=>OutputImg0_75, OutputImg0(74)=>OutputImg0_74, 
      OutputImg0(73)=>OutputImg0_73, OutputImg0(72)=>OutputImg0_72, 
      OutputImg0(71)=>OutputImg0_71, OutputImg0(70)=>OutputImg0_70, 
      OutputImg0(69)=>OutputImg0_69, OutputImg0(68)=>OutputImg0_68, 
      OutputImg0(67)=>OutputImg0_67, OutputImg0(66)=>OutputImg0_66, 
      OutputImg0(65)=>OutputImg0_65, OutputImg0(64)=>OutputImg0_64, 
      OutputImg0(63)=>OutputImg0_63, OutputImg0(62)=>OutputImg0_62, 
      OutputImg0(61)=>OutputImg0_61, OutputImg0(60)=>OutputImg0_60, 
      OutputImg0(59)=>OutputImg0_59, OutputImg0(58)=>OutputImg0_58, 
      OutputImg0(57)=>OutputImg0_57, OutputImg0(56)=>OutputImg0_56, 
      OutputImg0(55)=>OutputImg0_55, OutputImg0(54)=>OutputImg0_54, 
      OutputImg0(53)=>OutputImg0_53, OutputImg0(52)=>OutputImg0_52, 
      OutputImg0(51)=>OutputImg0_51, OutputImg0(50)=>OutputImg0_50, 
      OutputImg0(49)=>OutputImg0_49, OutputImg0(48)=>OutputImg0_48, 
      OutputImg0(47)=>OutputImg0_47, OutputImg0(46)=>OutputImg0_46, 
      OutputImg0(45)=>OutputImg0_45, OutputImg0(44)=>OutputImg0_44, 
      OutputImg0(43)=>OutputImg0_43, OutputImg0(42)=>OutputImg0_42, 
      OutputImg0(41)=>OutputImg0_41, OutputImg0(40)=>OutputImg0_40, 
      OutputImg0(39)=>OutputImg0_39, OutputImg0(38)=>OutputImg0_38, 
      OutputImg0(37)=>OutputImg0_37, OutputImg0(36)=>OutputImg0_36, 
      OutputImg0(35)=>OutputImg0_35, OutputImg0(34)=>OutputImg0_34, 
      OutputImg0(33)=>OutputImg0_33, OutputImg0(32)=>OutputImg0_32, 
      OutputImg0(31)=>OutputImg0_31, OutputImg0(30)=>OutputImg0_30, 
      OutputImg0(29)=>OutputImg0_29, OutputImg0(28)=>OutputImg0_28, 
      OutputImg0(27)=>OutputImg0_27, OutputImg0(26)=>OutputImg0_26, 
      OutputImg0(25)=>OutputImg0_25, OutputImg0(24)=>OutputImg0_24, 
      OutputImg0(23)=>OutputImg0_23, OutputImg0(22)=>OutputImg0_22, 
      OutputImg0(21)=>OutputImg0_21, OutputImg0(20)=>OutputImg0_20, 
      OutputImg0(19)=>OutputImg0_19, OutputImg0(18)=>OutputImg0_18, 
      OutputImg0(17)=>OutputImg0_17, OutputImg0(16)=>OutputImg0_16, 
      OutputImg0(15)=>OutputImg0_15, OutputImg0(14)=>OutputImg0_14, 
      OutputImg0(13)=>OutputImg0_13, OutputImg0(12)=>OutputImg0_12, 
      OutputImg0(11)=>OutputImg0_11, OutputImg0(10)=>OutputImg0_10, 
      OutputImg0(9)=>OutputImg0_9, OutputImg0(8)=>OutputImg0_8, 
      OutputImg0(7)=>OutputImg0_7, OutputImg0(6)=>OutputImg0_6, 
      OutputImg0(5)=>OutputImg0_5, OutputImg0(4)=>OutputImg0_4, 
      OutputImg0(3)=>OutputImg0_3, OutputImg0(2)=>OutputImg0_2, 
      OutputImg0(1)=>OutputImg0_1, OutputImg0(0)=>OutputImg0_0, 
      OutputImg1(79)=>OutputImg1_79, OutputImg1(78)=>OutputImg1_78, 
      OutputImg1(77)=>OutputImg1_77, OutputImg1(76)=>OutputImg1_76, 
      OutputImg1(75)=>OutputImg1_75, OutputImg1(74)=>OutputImg1_74, 
      OutputImg1(73)=>OutputImg1_73, OutputImg1(72)=>OutputImg1_72, 
      OutputImg1(71)=>OutputImg1_71, OutputImg1(70)=>OutputImg1_70, 
      OutputImg1(69)=>OutputImg1_69, OutputImg1(68)=>OutputImg1_68, 
      OutputImg1(67)=>OutputImg1_67, OutputImg1(66)=>OutputImg1_66, 
      OutputImg1(65)=>OutputImg1_65, OutputImg1(64)=>OutputImg1_64, 
      OutputImg1(63)=>OutputImg1_63, OutputImg1(62)=>OutputImg1_62, 
      OutputImg1(61)=>OutputImg1_61, OutputImg1(60)=>OutputImg1_60, 
      OutputImg1(59)=>OutputImg1_59, OutputImg1(58)=>OutputImg1_58, 
      OutputImg1(57)=>OutputImg1_57, OutputImg1(56)=>OutputImg1_56, 
      OutputImg1(55)=>OutputImg1_55, OutputImg1(54)=>OutputImg1_54, 
      OutputImg1(53)=>OutputImg1_53, OutputImg1(52)=>OutputImg1_52, 
      OutputImg1(51)=>OutputImg1_51, OutputImg1(50)=>OutputImg1_50, 
      OutputImg1(49)=>OutputImg1_49, OutputImg1(48)=>OutputImg1_48, 
      OutputImg1(47)=>OutputImg1_47, OutputImg1(46)=>OutputImg1_46, 
      OutputImg1(45)=>OutputImg1_45, OutputImg1(44)=>OutputImg1_44, 
      OutputImg1(43)=>OutputImg1_43, OutputImg1(42)=>OutputImg1_42, 
      OutputImg1(41)=>OutputImg1_41, OutputImg1(40)=>OutputImg1_40, 
      OutputImg1(39)=>OutputImg1_39, OutputImg1(38)=>OutputImg1_38, 
      OutputImg1(37)=>OutputImg1_37, OutputImg1(36)=>OutputImg1_36, 
      OutputImg1(35)=>OutputImg1_35, OutputImg1(34)=>OutputImg1_34, 
      OutputImg1(33)=>OutputImg1_33, OutputImg1(32)=>OutputImg1_32, 
      OutputImg1(31)=>OutputImg1_31, OutputImg1(30)=>OutputImg1_30, 
      OutputImg1(29)=>OutputImg1_29, OutputImg1(28)=>OutputImg1_28, 
      OutputImg1(27)=>OutputImg1_27, OutputImg1(26)=>OutputImg1_26, 
      OutputImg1(25)=>OutputImg1_25, OutputImg1(24)=>OutputImg1_24, 
      OutputImg1(23)=>OutputImg1_23, OutputImg1(22)=>OutputImg1_22, 
      OutputImg1(21)=>OutputImg1_21, OutputImg1(20)=>OutputImg1_20, 
      OutputImg1(19)=>OutputImg1_19, OutputImg1(18)=>OutputImg1_18, 
      OutputImg1(17)=>OutputImg1_17, OutputImg1(16)=>OutputImg1_16, 
      OutputImg1(15)=>OutputImg1_15, OutputImg1(14)=>OutputImg1_14, 
      OutputImg1(13)=>OutputImg1_13, OutputImg1(12)=>OutputImg1_12, 
      OutputImg1(11)=>OutputImg1_11, OutputImg1(10)=>OutputImg1_10, 
      OutputImg1(9)=>OutputImg1_9, OutputImg1(8)=>OutputImg1_8, 
      OutputImg1(7)=>OutputImg1_7, OutputImg1(6)=>OutputImg1_6, 
      OutputImg1(5)=>OutputImg1_5, OutputImg1(4)=>OutputImg1_4, 
      OutputImg1(3)=>OutputImg1_3, OutputImg1(2)=>OutputImg1_2, 
      OutputImg1(1)=>OutputImg1_1, OutputImg1(0)=>OutputImg1_0, 
      OutputImg2(79)=>OutputImg2_79, OutputImg2(78)=>OutputImg2_78, 
      OutputImg2(77)=>OutputImg2_77, OutputImg2(76)=>OutputImg2_76, 
      OutputImg2(75)=>OutputImg2_75, OutputImg2(74)=>OutputImg2_74, 
      OutputImg2(73)=>OutputImg2_73, OutputImg2(72)=>OutputImg2_72, 
      OutputImg2(71)=>OutputImg2_71, OutputImg2(70)=>OutputImg2_70, 
      OutputImg2(69)=>OutputImg2_69, OutputImg2(68)=>OutputImg2_68, 
      OutputImg2(67)=>OutputImg2_67, OutputImg2(66)=>OutputImg2_66, 
      OutputImg2(65)=>OutputImg2_65, OutputImg2(64)=>OutputImg2_64, 
      OutputImg2(63)=>OutputImg2_63, OutputImg2(62)=>OutputImg2_62, 
      OutputImg2(61)=>OutputImg2_61, OutputImg2(60)=>OutputImg2_60, 
      OutputImg2(59)=>OutputImg2_59, OutputImg2(58)=>OutputImg2_58, 
      OutputImg2(57)=>OutputImg2_57, OutputImg2(56)=>OutputImg2_56, 
      OutputImg2(55)=>OutputImg2_55, OutputImg2(54)=>OutputImg2_54, 
      OutputImg2(53)=>OutputImg2_53, OutputImg2(52)=>OutputImg2_52, 
      OutputImg2(51)=>OutputImg2_51, OutputImg2(50)=>OutputImg2_50, 
      OutputImg2(49)=>OutputImg2_49, OutputImg2(48)=>OutputImg2_48, 
      OutputImg2(47)=>OutputImg2_47, OutputImg2(46)=>OutputImg2_46, 
      OutputImg2(45)=>OutputImg2_45, OutputImg2(44)=>OutputImg2_44, 
      OutputImg2(43)=>OutputImg2_43, OutputImg2(42)=>OutputImg2_42, 
      OutputImg2(41)=>OutputImg2_41, OutputImg2(40)=>OutputImg2_40, 
      OutputImg2(39)=>OutputImg2_39, OutputImg2(38)=>OutputImg2_38, 
      OutputImg2(37)=>OutputImg2_37, OutputImg2(36)=>OutputImg2_36, 
      OutputImg2(35)=>OutputImg2_35, OutputImg2(34)=>OutputImg2_34, 
      OutputImg2(33)=>OutputImg2_33, OutputImg2(32)=>OutputImg2_32, 
      OutputImg2(31)=>OutputImg2_31, OutputImg2(30)=>OutputImg2_30, 
      OutputImg2(29)=>OutputImg2_29, OutputImg2(28)=>OutputImg2_28, 
      OutputImg2(27)=>OutputImg2_27, OutputImg2(26)=>OutputImg2_26, 
      OutputImg2(25)=>OutputImg2_25, OutputImg2(24)=>OutputImg2_24, 
      OutputImg2(23)=>OutputImg2_23, OutputImg2(22)=>OutputImg2_22, 
      OutputImg2(21)=>OutputImg2_21, OutputImg2(20)=>OutputImg2_20, 
      OutputImg2(19)=>OutputImg2_19, OutputImg2(18)=>OutputImg2_18, 
      OutputImg2(17)=>OutputImg2_17, OutputImg2(16)=>OutputImg2_16, 
      OutputImg2(15)=>OutputImg2_15, OutputImg2(14)=>OutputImg2_14, 
      OutputImg2(13)=>OutputImg2_13, OutputImg2(12)=>OutputImg2_12, 
      OutputImg2(11)=>OutputImg2_11, OutputImg2(10)=>OutputImg2_10, 
      OutputImg2(9)=>OutputImg2_9, OutputImg2(8)=>OutputImg2_8, 
      OutputImg2(7)=>OutputImg2_7, OutputImg2(6)=>OutputImg2_6, 
      OutputImg2(5)=>OutputImg2_5, OutputImg2(4)=>OutputImg2_4, 
      OutputImg2(3)=>OutputImg2_3, OutputImg2(2)=>OutputImg2_2, 
      OutputImg2(1)=>OutputImg2_1, OutputImg2(0)=>OutputImg2_0, 
      OutputImg3(79)=>OutputImg3_79, OutputImg3(78)=>OutputImg3_78, 
      OutputImg3(77)=>OutputImg3_77, OutputImg3(76)=>OutputImg3_76, 
      OutputImg3(75)=>OutputImg3_75, OutputImg3(74)=>OutputImg3_74, 
      OutputImg3(73)=>OutputImg3_73, OutputImg3(72)=>OutputImg3_72, 
      OutputImg3(71)=>OutputImg3_71, OutputImg3(70)=>OutputImg3_70, 
      OutputImg3(69)=>OutputImg3_69, OutputImg3(68)=>OutputImg3_68, 
      OutputImg3(67)=>OutputImg3_67, OutputImg3(66)=>OutputImg3_66, 
      OutputImg3(65)=>OutputImg3_65, OutputImg3(64)=>OutputImg3_64, 
      OutputImg3(63)=>OutputImg3_63, OutputImg3(62)=>OutputImg3_62, 
      OutputImg3(61)=>OutputImg3_61, OutputImg3(60)=>OutputImg3_60, 
      OutputImg3(59)=>OutputImg3_59, OutputImg3(58)=>OutputImg3_58, 
      OutputImg3(57)=>OutputImg3_57, OutputImg3(56)=>OutputImg3_56, 
      OutputImg3(55)=>OutputImg3_55, OutputImg3(54)=>OutputImg3_54, 
      OutputImg3(53)=>OutputImg3_53, OutputImg3(52)=>OutputImg3_52, 
      OutputImg3(51)=>OutputImg3_51, OutputImg3(50)=>OutputImg3_50, 
      OutputImg3(49)=>OutputImg3_49, OutputImg3(48)=>OutputImg3_48, 
      OutputImg3(47)=>OutputImg3_47, OutputImg3(46)=>OutputImg3_46, 
      OutputImg3(45)=>OutputImg3_45, OutputImg3(44)=>OutputImg3_44, 
      OutputImg3(43)=>OutputImg3_43, OutputImg3(42)=>OutputImg3_42, 
      OutputImg3(41)=>OutputImg3_41, OutputImg3(40)=>OutputImg3_40, 
      OutputImg3(39)=>OutputImg3_39, OutputImg3(38)=>OutputImg3_38, 
      OutputImg3(37)=>OutputImg3_37, OutputImg3(36)=>OutputImg3_36, 
      OutputImg3(35)=>OutputImg3_35, OutputImg3(34)=>OutputImg3_34, 
      OutputImg3(33)=>OutputImg3_33, OutputImg3(32)=>OutputImg3_32, 
      OutputImg3(31)=>OutputImg3_31, OutputImg3(30)=>OutputImg3_30, 
      OutputImg3(29)=>OutputImg3_29, OutputImg3(28)=>OutputImg3_28, 
      OutputImg3(27)=>OutputImg3_27, OutputImg3(26)=>OutputImg3_26, 
      OutputImg3(25)=>OutputImg3_25, OutputImg3(24)=>OutputImg3_24, 
      OutputImg3(23)=>OutputImg3_23, OutputImg3(22)=>OutputImg3_22, 
      OutputImg3(21)=>OutputImg3_21, OutputImg3(20)=>OutputImg3_20, 
      OutputImg3(19)=>OutputImg3_19, OutputImg3(18)=>OutputImg3_18, 
      OutputImg3(17)=>OutputImg3_17, OutputImg3(16)=>OutputImg3_16, 
      OutputImg3(15)=>OutputImg3_15, OutputImg3(14)=>OutputImg3_14, 
      OutputImg3(13)=>OutputImg3_13, OutputImg3(12)=>OutputImg3_12, 
      OutputImg3(11)=>OutputImg3_11, OutputImg3(10)=>OutputImg3_10, 
      OutputImg3(9)=>OutputImg3_9, OutputImg3(8)=>OutputImg3_8, 
      OutputImg3(7)=>OutputImg3_7, OutputImg3(6)=>OutputImg3_6, 
      OutputImg3(5)=>OutputImg3_5, OutputImg3(4)=>OutputImg3_4, 
      OutputImg3(3)=>OutputImg3_3, OutputImg3(2)=>OutputImg3_2, 
      OutputImg3(1)=>OutputImg3_1, OutputImg3(0)=>OutputImg3_0, 
      OutputImg4(79)=>OutputImg4_79, OutputImg4(78)=>OutputImg4_78, 
      OutputImg4(77)=>OutputImg4_77, OutputImg4(76)=>OutputImg4_76, 
      OutputImg4(75)=>OutputImg4_75, OutputImg4(74)=>OutputImg4_74, 
      OutputImg4(73)=>OutputImg4_73, OutputImg4(72)=>OutputImg4_72, 
      OutputImg4(71)=>OutputImg4_71, OutputImg4(70)=>OutputImg4_70, 
      OutputImg4(69)=>OutputImg4_69, OutputImg4(68)=>OutputImg4_68, 
      OutputImg4(67)=>OutputImg4_67, OutputImg4(66)=>OutputImg4_66, 
      OutputImg4(65)=>OutputImg4_65, OutputImg4(64)=>OutputImg4_64, 
      OutputImg4(63)=>OutputImg4_63, OutputImg4(62)=>OutputImg4_62, 
      OutputImg4(61)=>OutputImg4_61, OutputImg4(60)=>OutputImg4_60, 
      OutputImg4(59)=>OutputImg4_59, OutputImg4(58)=>OutputImg4_58, 
      OutputImg4(57)=>OutputImg4_57, OutputImg4(56)=>OutputImg4_56, 
      OutputImg4(55)=>OutputImg4_55, OutputImg4(54)=>OutputImg4_54, 
      OutputImg4(53)=>OutputImg4_53, OutputImg4(52)=>OutputImg4_52, 
      OutputImg4(51)=>OutputImg4_51, OutputImg4(50)=>OutputImg4_50, 
      OutputImg4(49)=>OutputImg4_49, OutputImg4(48)=>OutputImg4_48, 
      OutputImg4(47)=>OutputImg4_47, OutputImg4(46)=>OutputImg4_46, 
      OutputImg4(45)=>OutputImg4_45, OutputImg4(44)=>OutputImg4_44, 
      OutputImg4(43)=>OutputImg4_43, OutputImg4(42)=>OutputImg4_42, 
      OutputImg4(41)=>OutputImg4_41, OutputImg4(40)=>OutputImg4_40, 
      OutputImg4(39)=>OutputImg4_39, OutputImg4(38)=>OutputImg4_38, 
      OutputImg4(37)=>OutputImg4_37, OutputImg4(36)=>OutputImg4_36, 
      OutputImg4(35)=>OutputImg4_35, OutputImg4(34)=>OutputImg4_34, 
      OutputImg4(33)=>OutputImg4_33, OutputImg4(32)=>OutputImg4_32, 
      OutputImg4(31)=>OutputImg4_31, OutputImg4(30)=>OutputImg4_30, 
      OutputImg4(29)=>OutputImg4_29, OutputImg4(28)=>OutputImg4_28, 
      OutputImg4(27)=>OutputImg4_27, OutputImg4(26)=>OutputImg4_26, 
      OutputImg4(25)=>OutputImg4_25, OutputImg4(24)=>OutputImg4_24, 
      OutputImg4(23)=>OutputImg4_23, OutputImg4(22)=>OutputImg4_22, 
      OutputImg4(21)=>OutputImg4_21, OutputImg4(20)=>OutputImg4_20, 
      OutputImg4(19)=>OutputImg4_19, OutputImg4(18)=>OutputImg4_18, 
      OutputImg4(17)=>OutputImg4_17, OutputImg4(16)=>OutputImg4_16, 
      OutputImg4(15)=>OutputImg4_15, OutputImg4(14)=>OutputImg4_14, 
      OutputImg4(13)=>OutputImg4_13, OutputImg4(12)=>OutputImg4_12, 
      OutputImg4(11)=>OutputImg4_11, OutputImg4(10)=>OutputImg4_10, 
      OutputImg4(9)=>OutputImg4_9, OutputImg4(8)=>OutputImg4_8, 
      OutputImg4(7)=>OutputImg4_7, OutputImg4(6)=>OutputImg4_6, 
      OutputImg4(5)=>OutputImg4_5, OutputImg4(4)=>OutputImg4_4, 
      OutputImg4(3)=>OutputImg4_3, OutputImg4(2)=>OutputImg4_2, 
      OutputImg4(1)=>OutputImg4_1, OutputImg4(0)=>OutputImg4_0, 
      outFilter0(399)=>Filter1_399, outFilter0(398)=>Filter1_398, 
      outFilter0(397)=>Filter1_397, outFilter0(396)=>Filter1_396, 
      outFilter0(395)=>Filter1_395, outFilter0(394)=>Filter1_394, 
      outFilter0(393)=>Filter1_393, outFilter0(392)=>Filter1_392, 
      outFilter0(391)=>Filter1_391, outFilter0(390)=>Filter1_390, 
      outFilter0(389)=>Filter1_389, outFilter0(388)=>Filter1_388, 
      outFilter0(387)=>Filter1_387, outFilter0(386)=>Filter1_386, 
      outFilter0(385)=>Filter1_385, outFilter0(384)=>Filter1_384, 
      outFilter0(383)=>Filter1_383, outFilter0(382)=>Filter1_382, 
      outFilter0(381)=>Filter1_381, outFilter0(380)=>Filter1_380, 
      outFilter0(379)=>Filter1_379, outFilter0(378)=>Filter1_378, 
      outFilter0(377)=>Filter1_377, outFilter0(376)=>Filter1_376, 
      outFilter0(375)=>Filter1_375, outFilter0(374)=>Filter1_374, 
      outFilter0(373)=>Filter1_373, outFilter0(372)=>Filter1_372, 
      outFilter0(371)=>Filter1_371, outFilter0(370)=>Filter1_370, 
      outFilter0(369)=>Filter1_369, outFilter0(368)=>Filter1_368, 
      outFilter0(367)=>Filter1_367, outFilter0(366)=>Filter1_366, 
      outFilter0(365)=>Filter1_365, outFilter0(364)=>Filter1_364, 
      outFilter0(363)=>Filter1_363, outFilter0(362)=>Filter1_362, 
      outFilter0(361)=>Filter1_361, outFilter0(360)=>Filter1_360, 
      outFilter0(359)=>Filter1_359, outFilter0(358)=>Filter1_358, 
      outFilter0(357)=>Filter1_357, outFilter0(356)=>Filter1_356, 
      outFilter0(355)=>Filter1_355, outFilter0(354)=>Filter1_354, 
      outFilter0(353)=>Filter1_353, outFilter0(352)=>Filter1_352, 
      outFilter0(351)=>Filter1_351, outFilter0(350)=>Filter1_350, 
      outFilter0(349)=>Filter1_349, outFilter0(348)=>Filter1_348, 
      outFilter0(347)=>Filter1_347, outFilter0(346)=>Filter1_346, 
      outFilter0(345)=>Filter1_345, outFilter0(344)=>Filter1_344, 
      outFilter0(343)=>Filter1_343, outFilter0(342)=>Filter1_342, 
      outFilter0(341)=>Filter1_341, outFilter0(340)=>Filter1_340, 
      outFilter0(339)=>Filter1_339, outFilter0(338)=>Filter1_338, 
      outFilter0(337)=>Filter1_337, outFilter0(336)=>Filter1_336, 
      outFilter0(335)=>Filter1_335, outFilter0(334)=>Filter1_334, 
      outFilter0(333)=>Filter1_333, outFilter0(332)=>Filter1_332, 
      outFilter0(331)=>Filter1_331, outFilter0(330)=>Filter1_330, 
      outFilter0(329)=>Filter1_329, outFilter0(328)=>Filter1_328, 
      outFilter0(327)=>Filter1_327, outFilter0(326)=>Filter1_326, 
      outFilter0(325)=>Filter1_325, outFilter0(324)=>Filter1_324, 
      outFilter0(323)=>Filter1_323, outFilter0(322)=>Filter1_322, 
      outFilter0(321)=>Filter1_321, outFilter0(320)=>Filter1_320, 
      outFilter0(319)=>Filter1_319, outFilter0(318)=>Filter1_318, 
      outFilter0(317)=>Filter1_317, outFilter0(316)=>Filter1_316, 
      outFilter0(315)=>Filter1_315, outFilter0(314)=>Filter1_314, 
      outFilter0(313)=>Filter1_313, outFilter0(312)=>Filter1_312, 
      outFilter0(311)=>Filter1_311, outFilter0(310)=>Filter1_310, 
      outFilter0(309)=>Filter1_309, outFilter0(308)=>Filter1_308, 
      outFilter0(307)=>Filter1_307, outFilter0(306)=>Filter1_306, 
      outFilter0(305)=>Filter1_305, outFilter0(304)=>Filter1_304, 
      outFilter0(303)=>Filter1_303, outFilter0(302)=>Filter1_302, 
      outFilter0(301)=>Filter1_301, outFilter0(300)=>Filter1_300, 
      outFilter0(299)=>Filter1_299, outFilter0(298)=>Filter1_298, 
      outFilter0(297)=>Filter1_297, outFilter0(296)=>Filter1_296, 
      outFilter0(295)=>Filter1_295, outFilter0(294)=>Filter1_294, 
      outFilter0(293)=>Filter1_293, outFilter0(292)=>Filter1_292, 
      outFilter0(291)=>Filter1_291, outFilter0(290)=>Filter1_290, 
      outFilter0(289)=>Filter1_289, outFilter0(288)=>Filter1_288, 
      outFilter0(287)=>Filter1_287, outFilter0(286)=>Filter1_286, 
      outFilter0(285)=>Filter1_285, outFilter0(284)=>Filter1_284, 
      outFilter0(283)=>Filter1_283, outFilter0(282)=>Filter1_282, 
      outFilter0(281)=>Filter1_281, outFilter0(280)=>Filter1_280, 
      outFilter0(279)=>Filter1_279, outFilter0(278)=>Filter1_278, 
      outFilter0(277)=>Filter1_277, outFilter0(276)=>Filter1_276, 
      outFilter0(275)=>Filter1_275, outFilter0(274)=>Filter1_274, 
      outFilter0(273)=>Filter1_273, outFilter0(272)=>Filter1_272, 
      outFilter0(271)=>Filter1_271, outFilter0(270)=>Filter1_270, 
      outFilter0(269)=>Filter1_269, outFilter0(268)=>Filter1_268, 
      outFilter0(267)=>Filter1_267, outFilter0(266)=>Filter1_266, 
      outFilter0(265)=>Filter1_265, outFilter0(264)=>Filter1_264, 
      outFilter0(263)=>Filter1_263, outFilter0(262)=>Filter1_262, 
      outFilter0(261)=>Filter1_261, outFilter0(260)=>Filter1_260, 
      outFilter0(259)=>Filter1_259, outFilter0(258)=>Filter1_258, 
      outFilter0(257)=>Filter1_257, outFilter0(256)=>Filter1_256, 
      outFilter0(255)=>Filter1_255, outFilter0(254)=>Filter1_254, 
      outFilter0(253)=>Filter1_253, outFilter0(252)=>Filter1_252, 
      outFilter0(251)=>Filter1_251, outFilter0(250)=>Filter1_250, 
      outFilter0(249)=>Filter1_249, outFilter0(248)=>Filter1_248, 
      outFilter0(247)=>Filter1_247, outFilter0(246)=>Filter1_246, 
      outFilter0(245)=>Filter1_245, outFilter0(244)=>Filter1_244, 
      outFilter0(243)=>Filter1_243, outFilter0(242)=>Filter1_242, 
      outFilter0(241)=>Filter1_241, outFilter0(240)=>Filter1_240, 
      outFilter0(239)=>Filter1_239, outFilter0(238)=>Filter1_238, 
      outFilter0(237)=>Filter1_237, outFilter0(236)=>Filter1_236, 
      outFilter0(235)=>Filter1_235, outFilter0(234)=>Filter1_234, 
      outFilter0(233)=>Filter1_233, outFilter0(232)=>Filter1_232, 
      outFilter0(231)=>Filter1_231, outFilter0(230)=>Filter1_230, 
      outFilter0(229)=>Filter1_229, outFilter0(228)=>Filter1_228, 
      outFilter0(227)=>Filter1_227, outFilter0(226)=>Filter1_226, 
      outFilter0(225)=>Filter1_225, outFilter0(224)=>Filter1_224, 
      outFilter0(223)=>Filter1_223, outFilter0(222)=>Filter1_222, 
      outFilter0(221)=>Filter1_221, outFilter0(220)=>Filter1_220, 
      outFilter0(219)=>Filter1_219, outFilter0(218)=>Filter1_218, 
      outFilter0(217)=>Filter1_217, outFilter0(216)=>Filter1_216, 
      outFilter0(215)=>Filter1_215, outFilter0(214)=>Filter1_214, 
      outFilter0(213)=>Filter1_213, outFilter0(212)=>Filter1_212, 
      outFilter0(211)=>Filter1_211, outFilter0(210)=>Filter1_210, 
      outFilter0(209)=>Filter1_209, outFilter0(208)=>Filter1_208, 
      outFilter0(207)=>Filter1_207, outFilter0(206)=>Filter1_206, 
      outFilter0(205)=>Filter1_205, outFilter0(204)=>Filter1_204, 
      outFilter0(203)=>Filter1_203, outFilter0(202)=>Filter1_202, 
      outFilter0(201)=>Filter1_201, outFilter0(200)=>Filter1_200, 
      outFilter0(199)=>Filter1_199, outFilter0(198)=>Filter1_198, 
      outFilter0(197)=>Filter1_197, outFilter0(196)=>Filter1_196, 
      outFilter0(195)=>Filter1_195, outFilter0(194)=>Filter1_194, 
      outFilter0(193)=>Filter1_193, outFilter0(192)=>Filter1_192, 
      outFilter0(191)=>Filter1_191, outFilter0(190)=>Filter1_190, 
      outFilter0(189)=>Filter1_189, outFilter0(188)=>Filter1_188, 
      outFilter0(187)=>Filter1_187, outFilter0(186)=>Filter1_186, 
      outFilter0(185)=>Filter1_185, outFilter0(184)=>Filter1_184, 
      outFilter0(183)=>Filter1_183, outFilter0(182)=>Filter1_182, 
      outFilter0(181)=>Filter1_181, outFilter0(180)=>Filter1_180, 
      outFilter0(179)=>Filter1_179, outFilter0(178)=>Filter1_178, 
      outFilter0(177)=>Filter1_177, outFilter0(176)=>Filter1_176, 
      outFilter0(175)=>Filter1_175, outFilter0(174)=>Filter1_174, 
      outFilter0(173)=>Filter1_173, outFilter0(172)=>Filter1_172, 
      outFilter0(171)=>Filter1_171, outFilter0(170)=>Filter1_170, 
      outFilter0(169)=>Filter1_169, outFilter0(168)=>Filter1_168, 
      outFilter0(167)=>Filter1_167, outFilter0(166)=>Filter1_166, 
      outFilter0(165)=>Filter1_165, outFilter0(164)=>Filter1_164, 
      outFilter0(163)=>Filter1_163, outFilter0(162)=>Filter1_162, 
      outFilter0(161)=>Filter1_161, outFilter0(160)=>Filter1_160, 
      outFilter0(159)=>Filter1_159, outFilter0(158)=>Filter1_158, 
      outFilter0(157)=>Filter1_157, outFilter0(156)=>Filter1_156, 
      outFilter0(155)=>Filter1_155, outFilter0(154)=>Filter1_154, 
      outFilter0(153)=>Filter1_153, outFilter0(152)=>Filter1_152, 
      outFilter0(151)=>Filter1_151, outFilter0(150)=>Filter1_150, 
      outFilter0(149)=>Filter1_149, outFilter0(148)=>Filter1_148, 
      outFilter0(147)=>Filter1_147, outFilter0(146)=>Filter1_146, 
      outFilter0(145)=>Filter1_145, outFilter0(144)=>Filter1_144, 
      outFilter0(143)=>Filter1_143, outFilter0(142)=>Filter1_142, 
      outFilter0(141)=>Filter1_141, outFilter0(140)=>Filter1_140, 
      outFilter0(139)=>Filter1_139, outFilter0(138)=>Filter1_138, 
      outFilter0(137)=>Filter1_137, outFilter0(136)=>Filter1_136, 
      outFilter0(135)=>Filter1_135, outFilter0(134)=>Filter1_134, 
      outFilter0(133)=>Filter1_133, outFilter0(132)=>Filter1_132, 
      outFilter0(131)=>Filter1_131, outFilter0(130)=>Filter1_130, 
      outFilter0(129)=>Filter1_129, outFilter0(128)=>Filter1_128, 
      outFilter0(127)=>Filter1_127, outFilter0(126)=>Filter1_126, 
      outFilter0(125)=>Filter1_125, outFilter0(124)=>Filter1_124, 
      outFilter0(123)=>Filter1_123, outFilter0(122)=>Filter1_122, 
      outFilter0(121)=>Filter1_121, outFilter0(120)=>Filter1_120, 
      outFilter0(119)=>Filter1_119, outFilter0(118)=>Filter1_118, 
      outFilter0(117)=>Filter1_117, outFilter0(116)=>Filter1_116, 
      outFilter0(115)=>Filter1_115, outFilter0(114)=>Filter1_114, 
      outFilter0(113)=>Filter1_113, outFilter0(112)=>Filter1_112, 
      outFilter0(111)=>Filter1_111, outFilter0(110)=>Filter1_110, 
      outFilter0(109)=>Filter1_109, outFilter0(108)=>Filter1_108, 
      outFilter0(107)=>Filter1_107, outFilter0(106)=>Filter1_106, 
      outFilter0(105)=>Filter1_105, outFilter0(104)=>Filter1_104, 
      outFilter0(103)=>Filter1_103, outFilter0(102)=>Filter1_102, 
      outFilter0(101)=>Filter1_101, outFilter0(100)=>Filter1_100, 
      outFilter0(99)=>Filter1_99, outFilter0(98)=>Filter1_98, outFilter0(97)
      =>Filter1_97, outFilter0(96)=>Filter1_96, outFilter0(95)=>Filter1_95, 
      outFilter0(94)=>Filter1_94, outFilter0(93)=>Filter1_93, outFilter0(92)
      =>Filter1_92, outFilter0(91)=>Filter1_91, outFilter0(90)=>Filter1_90, 
      outFilter0(89)=>Filter1_89, outFilter0(88)=>Filter1_88, outFilter0(87)
      =>Filter1_87, outFilter0(86)=>Filter1_86, outFilter0(85)=>Filter1_85, 
      outFilter0(84)=>Filter1_84, outFilter0(83)=>Filter1_83, outFilter0(82)
      =>Filter1_82, outFilter0(81)=>Filter1_81, outFilter0(80)=>Filter1_80, 
      outFilter0(79)=>Filter1_79, outFilter0(78)=>Filter1_78, outFilter0(77)
      =>Filter1_77, outFilter0(76)=>Filter1_76, outFilter0(75)=>Filter1_75, 
      outFilter0(74)=>Filter1_74, outFilter0(73)=>Filter1_73, outFilter0(72)
      =>Filter1_72, outFilter0(71)=>Filter1_71, outFilter0(70)=>Filter1_70, 
      outFilter0(69)=>Filter1_69, outFilter0(68)=>Filter1_68, outFilter0(67)
      =>Filter1_67, outFilter0(66)=>Filter1_66, outFilter0(65)=>Filter1_65, 
      outFilter0(64)=>Filter1_64, outFilter0(63)=>Filter1_63, outFilter0(62)
      =>Filter1_62, outFilter0(61)=>Filter1_61, outFilter0(60)=>Filter1_60, 
      outFilter0(59)=>Filter1_59, outFilter0(58)=>Filter1_58, outFilter0(57)
      =>Filter1_57, outFilter0(56)=>Filter1_56, outFilter0(55)=>Filter1_55, 
      outFilter0(54)=>Filter1_54, outFilter0(53)=>Filter1_53, outFilter0(52)
      =>Filter1_52, outFilter0(51)=>Filter1_51, outFilter0(50)=>Filter1_50, 
      outFilter0(49)=>Filter1_49, outFilter0(48)=>Filter1_48, outFilter0(47)
      =>Filter1_47, outFilter0(46)=>Filter1_46, outFilter0(45)=>Filter1_45, 
      outFilter0(44)=>Filter1_44, outFilter0(43)=>Filter1_43, outFilter0(42)
      =>Filter1_42, outFilter0(41)=>Filter1_41, outFilter0(40)=>Filter1_40, 
      outFilter0(39)=>Filter1_39, outFilter0(38)=>Filter1_38, outFilter0(37)
      =>Filter1_37, outFilter0(36)=>Filter1_36, outFilter0(35)=>Filter1_35, 
      outFilter0(34)=>Filter1_34, outFilter0(33)=>Filter1_33, outFilter0(32)
      =>Filter1_32, outFilter0(31)=>Filter1_31, outFilter0(30)=>Filter1_30, 
      outFilter0(29)=>Filter1_29, outFilter0(28)=>Filter1_28, outFilter0(27)
      =>Filter1_27, outFilter0(26)=>Filter1_26, outFilter0(25)=>Filter1_25, 
      outFilter0(24)=>Filter1_24, outFilter0(23)=>Filter1_23, outFilter0(22)
      =>Filter1_22, outFilter0(21)=>Filter1_21, outFilter0(20)=>Filter1_20, 
      outFilter0(19)=>Filter1_19, outFilter0(18)=>Filter1_18, outFilter0(17)
      =>Filter1_17, outFilter0(16)=>Filter1_16, outFilter0(15)=>Filter1_15, 
      outFilter0(14)=>Filter1_14, outFilter0(13)=>Filter1_13, outFilter0(12)
      =>Filter1_12, outFilter0(11)=>Filter1_11, outFilter0(10)=>Filter1_10, 
      outFilter0(9)=>Filter1_9, outFilter0(8)=>Filter1_8, outFilter0(7)=>
      Filter1_7, outFilter0(6)=>Filter1_6, outFilter0(5)=>Filter1_5, 
      outFilter0(4)=>Filter1_4, outFilter0(3)=>Filter1_3, outFilter0(2)=>
      Filter1_2, outFilter0(1)=>Filter1_1, outFilter0(0)=>Filter1_0, 
      outFilter1(399)=>Filter2_399, outFilter1(398)=>Filter2_398, 
      outFilter1(397)=>Filter2_397, outFilter1(396)=>Filter2_396, 
      outFilter1(395)=>Filter2_395, outFilter1(394)=>Filter2_394, 
      outFilter1(393)=>Filter2_393, outFilter1(392)=>Filter2_392, 
      outFilter1(391)=>Filter2_391, outFilter1(390)=>Filter2_390, 
      outFilter1(389)=>Filter2_389, outFilter1(388)=>Filter2_388, 
      outFilter1(387)=>Filter2_387, outFilter1(386)=>Filter2_386, 
      outFilter1(385)=>Filter2_385, outFilter1(384)=>Filter2_384, 
      outFilter1(383)=>Filter2_383, outFilter1(382)=>Filter2_382, 
      outFilter1(381)=>Filter2_381, outFilter1(380)=>Filter2_380, 
      outFilter1(379)=>Filter2_379, outFilter1(378)=>Filter2_378, 
      outFilter1(377)=>Filter2_377, outFilter1(376)=>Filter2_376, 
      outFilter1(375)=>Filter2_375, outFilter1(374)=>Filter2_374, 
      outFilter1(373)=>Filter2_373, outFilter1(372)=>Filter2_372, 
      outFilter1(371)=>Filter2_371, outFilter1(370)=>Filter2_370, 
      outFilter1(369)=>Filter2_369, outFilter1(368)=>Filter2_368, 
      outFilter1(367)=>Filter2_367, outFilter1(366)=>Filter2_366, 
      outFilter1(365)=>Filter2_365, outFilter1(364)=>Filter2_364, 
      outFilter1(363)=>Filter2_363, outFilter1(362)=>Filter2_362, 
      outFilter1(361)=>Filter2_361, outFilter1(360)=>Filter2_360, 
      outFilter1(359)=>Filter2_359, outFilter1(358)=>Filter2_358, 
      outFilter1(357)=>Filter2_357, outFilter1(356)=>Filter2_356, 
      outFilter1(355)=>Filter2_355, outFilter1(354)=>Filter2_354, 
      outFilter1(353)=>Filter2_353, outFilter1(352)=>Filter2_352, 
      outFilter1(351)=>Filter2_351, outFilter1(350)=>Filter2_350, 
      outFilter1(349)=>Filter2_349, outFilter1(348)=>Filter2_348, 
      outFilter1(347)=>Filter2_347, outFilter1(346)=>Filter2_346, 
      outFilter1(345)=>Filter2_345, outFilter1(344)=>Filter2_344, 
      outFilter1(343)=>Filter2_343, outFilter1(342)=>Filter2_342, 
      outFilter1(341)=>Filter2_341, outFilter1(340)=>Filter2_340, 
      outFilter1(339)=>Filter2_339, outFilter1(338)=>Filter2_338, 
      outFilter1(337)=>Filter2_337, outFilter1(336)=>Filter2_336, 
      outFilter1(335)=>Filter2_335, outFilter1(334)=>Filter2_334, 
      outFilter1(333)=>Filter2_333, outFilter1(332)=>Filter2_332, 
      outFilter1(331)=>Filter2_331, outFilter1(330)=>Filter2_330, 
      outFilter1(329)=>Filter2_329, outFilter1(328)=>Filter2_328, 
      outFilter1(327)=>Filter2_327, outFilter1(326)=>Filter2_326, 
      outFilter1(325)=>Filter2_325, outFilter1(324)=>Filter2_324, 
      outFilter1(323)=>Filter2_323, outFilter1(322)=>Filter2_322, 
      outFilter1(321)=>Filter2_321, outFilter1(320)=>Filter2_320, 
      outFilter1(319)=>Filter2_319, outFilter1(318)=>Filter2_318, 
      outFilter1(317)=>Filter2_317, outFilter1(316)=>Filter2_316, 
      outFilter1(315)=>Filter2_315, outFilter1(314)=>Filter2_314, 
      outFilter1(313)=>Filter2_313, outFilter1(312)=>Filter2_312, 
      outFilter1(311)=>Filter2_311, outFilter1(310)=>Filter2_310, 
      outFilter1(309)=>Filter2_309, outFilter1(308)=>Filter2_308, 
      outFilter1(307)=>Filter2_307, outFilter1(306)=>Filter2_306, 
      outFilter1(305)=>Filter2_305, outFilter1(304)=>Filter2_304, 
      outFilter1(303)=>Filter2_303, outFilter1(302)=>Filter2_302, 
      outFilter1(301)=>Filter2_301, outFilter1(300)=>Filter2_300, 
      outFilter1(299)=>Filter2_299, outFilter1(298)=>Filter2_298, 
      outFilter1(297)=>Filter2_297, outFilter1(296)=>Filter2_296, 
      outFilter1(295)=>Filter2_295, outFilter1(294)=>Filter2_294, 
      outFilter1(293)=>Filter2_293, outFilter1(292)=>Filter2_292, 
      outFilter1(291)=>Filter2_291, outFilter1(290)=>Filter2_290, 
      outFilter1(289)=>Filter2_289, outFilter1(288)=>Filter2_288, 
      outFilter1(287)=>Filter2_287, outFilter1(286)=>Filter2_286, 
      outFilter1(285)=>Filter2_285, outFilter1(284)=>Filter2_284, 
      outFilter1(283)=>Filter2_283, outFilter1(282)=>Filter2_282, 
      outFilter1(281)=>Filter2_281, outFilter1(280)=>Filter2_280, 
      outFilter1(279)=>Filter2_279, outFilter1(278)=>Filter2_278, 
      outFilter1(277)=>Filter2_277, outFilter1(276)=>Filter2_276, 
      outFilter1(275)=>Filter2_275, outFilter1(274)=>Filter2_274, 
      outFilter1(273)=>Filter2_273, outFilter1(272)=>Filter2_272, 
      outFilter1(271)=>Filter2_271, outFilter1(270)=>Filter2_270, 
      outFilter1(269)=>Filter2_269, outFilter1(268)=>Filter2_268, 
      outFilter1(267)=>Filter2_267, outFilter1(266)=>Filter2_266, 
      outFilter1(265)=>Filter2_265, outFilter1(264)=>Filter2_264, 
      outFilter1(263)=>Filter2_263, outFilter1(262)=>Filter2_262, 
      outFilter1(261)=>Filter2_261, outFilter1(260)=>Filter2_260, 
      outFilter1(259)=>Filter2_259, outFilter1(258)=>Filter2_258, 
      outFilter1(257)=>Filter2_257, outFilter1(256)=>Filter2_256, 
      outFilter1(255)=>Filter2_255, outFilter1(254)=>Filter2_254, 
      outFilter1(253)=>Filter2_253, outFilter1(252)=>Filter2_252, 
      outFilter1(251)=>Filter2_251, outFilter1(250)=>Filter2_250, 
      outFilter1(249)=>Filter2_249, outFilter1(248)=>Filter2_248, 
      outFilter1(247)=>Filter2_247, outFilter1(246)=>Filter2_246, 
      outFilter1(245)=>Filter2_245, outFilter1(244)=>Filter2_244, 
      outFilter1(243)=>Filter2_243, outFilter1(242)=>Filter2_242, 
      outFilter1(241)=>Filter2_241, outFilter1(240)=>Filter2_240, 
      outFilter1(239)=>Filter2_239, outFilter1(238)=>Filter2_238, 
      outFilter1(237)=>Filter2_237, outFilter1(236)=>Filter2_236, 
      outFilter1(235)=>Filter2_235, outFilter1(234)=>Filter2_234, 
      outFilter1(233)=>Filter2_233, outFilter1(232)=>Filter2_232, 
      outFilter1(231)=>Filter2_231, outFilter1(230)=>Filter2_230, 
      outFilter1(229)=>Filter2_229, outFilter1(228)=>Filter2_228, 
      outFilter1(227)=>Filter2_227, outFilter1(226)=>Filter2_226, 
      outFilter1(225)=>Filter2_225, outFilter1(224)=>Filter2_224, 
      outFilter1(223)=>Filter2_223, outFilter1(222)=>Filter2_222, 
      outFilter1(221)=>Filter2_221, outFilter1(220)=>Filter2_220, 
      outFilter1(219)=>Filter2_219, outFilter1(218)=>Filter2_218, 
      outFilter1(217)=>Filter2_217, outFilter1(216)=>Filter2_216, 
      outFilter1(215)=>Filter2_215, outFilter1(214)=>Filter2_214, 
      outFilter1(213)=>Filter2_213, outFilter1(212)=>Filter2_212, 
      outFilter1(211)=>Filter2_211, outFilter1(210)=>Filter2_210, 
      outFilter1(209)=>Filter2_209, outFilter1(208)=>Filter2_208, 
      outFilter1(207)=>Filter2_207, outFilter1(206)=>Filter2_206, 
      outFilter1(205)=>Filter2_205, outFilter1(204)=>Filter2_204, 
      outFilter1(203)=>Filter2_203, outFilter1(202)=>Filter2_202, 
      outFilter1(201)=>Filter2_201, outFilter1(200)=>Filter2_200, 
      outFilter1(199)=>Filter2_199, outFilter1(198)=>Filter2_198, 
      outFilter1(197)=>Filter2_197, outFilter1(196)=>Filter2_196, 
      outFilter1(195)=>Filter2_195, outFilter1(194)=>Filter2_194, 
      outFilter1(193)=>Filter2_193, outFilter1(192)=>Filter2_192, 
      outFilter1(191)=>Filter2_191, outFilter1(190)=>Filter2_190, 
      outFilter1(189)=>Filter2_189, outFilter1(188)=>Filter2_188, 
      outFilter1(187)=>Filter2_187, outFilter1(186)=>Filter2_186, 
      outFilter1(185)=>Filter2_185, outFilter1(184)=>Filter2_184, 
      outFilter1(183)=>Filter2_183, outFilter1(182)=>Filter2_182, 
      outFilter1(181)=>Filter2_181, outFilter1(180)=>Filter2_180, 
      outFilter1(179)=>Filter2_179, outFilter1(178)=>Filter2_178, 
      outFilter1(177)=>Filter2_177, outFilter1(176)=>Filter2_176, 
      outFilter1(175)=>Filter2_175, outFilter1(174)=>Filter2_174, 
      outFilter1(173)=>Filter2_173, outFilter1(172)=>Filter2_172, 
      outFilter1(171)=>Filter2_171, outFilter1(170)=>Filter2_170, 
      outFilter1(169)=>Filter2_169, outFilter1(168)=>Filter2_168, 
      outFilter1(167)=>Filter2_167, outFilter1(166)=>Filter2_166, 
      outFilter1(165)=>Filter2_165, outFilter1(164)=>Filter2_164, 
      outFilter1(163)=>Filter2_163, outFilter1(162)=>Filter2_162, 
      outFilter1(161)=>Filter2_161, outFilter1(160)=>Filter2_160, 
      outFilter1(159)=>Filter2_159, outFilter1(158)=>Filter2_158, 
      outFilter1(157)=>Filter2_157, outFilter1(156)=>Filter2_156, 
      outFilter1(155)=>Filter2_155, outFilter1(154)=>Filter2_154, 
      outFilter1(153)=>Filter2_153, outFilter1(152)=>Filter2_152, 
      outFilter1(151)=>Filter2_151, outFilter1(150)=>Filter2_150, 
      outFilter1(149)=>Filter2_149, outFilter1(148)=>Filter2_148, 
      outFilter1(147)=>Filter2_147, outFilter1(146)=>Filter2_146, 
      outFilter1(145)=>Filter2_145, outFilter1(144)=>Filter2_144, 
      outFilter1(143)=>Filter2_143, outFilter1(142)=>Filter2_142, 
      outFilter1(141)=>Filter2_141, outFilter1(140)=>Filter2_140, 
      outFilter1(139)=>Filter2_139, outFilter1(138)=>Filter2_138, 
      outFilter1(137)=>Filter2_137, outFilter1(136)=>Filter2_136, 
      outFilter1(135)=>Filter2_135, outFilter1(134)=>Filter2_134, 
      outFilter1(133)=>Filter2_133, outFilter1(132)=>Filter2_132, 
      outFilter1(131)=>Filter2_131, outFilter1(130)=>Filter2_130, 
      outFilter1(129)=>Filter2_129, outFilter1(128)=>Filter2_128, 
      outFilter1(127)=>Filter2_127, outFilter1(126)=>Filter2_126, 
      outFilter1(125)=>Filter2_125, outFilter1(124)=>Filter2_124, 
      outFilter1(123)=>Filter2_123, outFilter1(122)=>Filter2_122, 
      outFilter1(121)=>Filter2_121, outFilter1(120)=>Filter2_120, 
      outFilter1(119)=>Filter2_119, outFilter1(118)=>Filter2_118, 
      outFilter1(117)=>Filter2_117, outFilter1(116)=>Filter2_116, 
      outFilter1(115)=>Filter2_115, outFilter1(114)=>Filter2_114, 
      outFilter1(113)=>Filter2_113, outFilter1(112)=>Filter2_112, 
      outFilter1(111)=>Filter2_111, outFilter1(110)=>Filter2_110, 
      outFilter1(109)=>Filter2_109, outFilter1(108)=>Filter2_108, 
      outFilter1(107)=>Filter2_107, outFilter1(106)=>Filter2_106, 
      outFilter1(105)=>Filter2_105, outFilter1(104)=>Filter2_104, 
      outFilter1(103)=>Filter2_103, outFilter1(102)=>Filter2_102, 
      outFilter1(101)=>Filter2_101, outFilter1(100)=>Filter2_100, 
      outFilter1(99)=>Filter2_99, outFilter1(98)=>Filter2_98, outFilter1(97)
      =>Filter2_97, outFilter1(96)=>Filter2_96, outFilter1(95)=>Filter2_95, 
      outFilter1(94)=>Filter2_94, outFilter1(93)=>Filter2_93, outFilter1(92)
      =>Filter2_92, outFilter1(91)=>Filter2_91, outFilter1(90)=>Filter2_90, 
      outFilter1(89)=>Filter2_89, outFilter1(88)=>Filter2_88, outFilter1(87)
      =>Filter2_87, outFilter1(86)=>Filter2_86, outFilter1(85)=>Filter2_85, 
      outFilter1(84)=>Filter2_84, outFilter1(83)=>Filter2_83, outFilter1(82)
      =>Filter2_82, outFilter1(81)=>Filter2_81, outFilter1(80)=>Filter2_80, 
      outFilter1(79)=>Filter2_79, outFilter1(78)=>Filter2_78, outFilter1(77)
      =>Filter2_77, outFilter1(76)=>Filter2_76, outFilter1(75)=>Filter2_75, 
      outFilter1(74)=>Filter2_74, outFilter1(73)=>Filter2_73, outFilter1(72)
      =>Filter2_72, outFilter1(71)=>Filter2_71, outFilter1(70)=>Filter2_70, 
      outFilter1(69)=>Filter2_69, outFilter1(68)=>Filter2_68, outFilter1(67)
      =>Filter2_67, outFilter1(66)=>Filter2_66, outFilter1(65)=>Filter2_65, 
      outFilter1(64)=>Filter2_64, outFilter1(63)=>Filter2_63, outFilter1(62)
      =>Filter2_62, outFilter1(61)=>Filter2_61, outFilter1(60)=>Filter2_60, 
      outFilter1(59)=>Filter2_59, outFilter1(58)=>Filter2_58, outFilter1(57)
      =>Filter2_57, outFilter1(56)=>Filter2_56, outFilter1(55)=>Filter2_55, 
      outFilter1(54)=>Filter2_54, outFilter1(53)=>Filter2_53, outFilter1(52)
      =>Filter2_52, outFilter1(51)=>Filter2_51, outFilter1(50)=>Filter2_50, 
      outFilter1(49)=>Filter2_49, outFilter1(48)=>Filter2_48, outFilter1(47)
      =>Filter2_47, outFilter1(46)=>Filter2_46, outFilter1(45)=>Filter2_45, 
      outFilter1(44)=>Filter2_44, outFilter1(43)=>Filter2_43, outFilter1(42)
      =>Filter2_42, outFilter1(41)=>Filter2_41, outFilter1(40)=>Filter2_40, 
      outFilter1(39)=>Filter2_39, outFilter1(38)=>Filter2_38, outFilter1(37)
      =>Filter2_37, outFilter1(36)=>Filter2_36, outFilter1(35)=>Filter2_35, 
      outFilter1(34)=>Filter2_34, outFilter1(33)=>Filter2_33, outFilter1(32)
      =>Filter2_32, outFilter1(31)=>Filter2_31, outFilter1(30)=>Filter2_30, 
      outFilter1(29)=>Filter2_29, outFilter1(28)=>Filter2_28, outFilter1(27)
      =>Filter2_27, outFilter1(26)=>Filter2_26, outFilter1(25)=>Filter2_25, 
      outFilter1(24)=>Filter2_24, outFilter1(23)=>Filter2_23, outFilter1(22)
      =>Filter2_22, outFilter1(21)=>Filter2_21, outFilter1(20)=>Filter2_20, 
      outFilter1(19)=>Filter2_19, outFilter1(18)=>Filter2_18, outFilter1(17)
      =>Filter2_17, outFilter1(16)=>Filter2_16, outFilter1(15)=>Filter2_15, 
      outFilter1(14)=>Filter2_14, outFilter1(13)=>Filter2_13, outFilter1(12)
      =>Filter2_12, outFilter1(11)=>Filter2_11, outFilter1(10)=>Filter2_10, 
      outFilter1(9)=>Filter2_9, outFilter1(8)=>Filter2_8, outFilter1(7)=>
      Filter2_7, outFilter1(6)=>Filter2_6, outFilter1(5)=>Filter2_5, 
      outFilter1(4)=>Filter2_4, outFilter1(3)=>Filter2_3, outFilter1(2)=>
      Filter2_2, outFilter1(1)=>Filter2_1, outFilter1(0)=>Filter2_0, 
      ConvOuput(15)=>ConvOuput_15, ConvOuput(14)=>ConvOuput_14, 
      ConvOuput(13)=>ConvOuput_13, ConvOuput(12)=>ConvOuput_12, 
      ConvOuput(11)=>ConvOuput_11, ConvOuput(10)=>ConvOuput_10, ConvOuput(9)
      =>ConvOuput_9, ConvOuput(8)=>ConvOuput_8, ConvOuput(7)=>ConvOuput_7, 
      ConvOuput(6)=>ConvOuput_6, ConvOuput(5)=>ConvOuput_5, ConvOuput(4)=>
      ConvOuput_4, ConvOuput(3)=>ConvOuput_3, ConvOuput(2)=>ConvOuput_2, 
      ConvOuput(1)=>ConvOuput_1, ConvOuput(0)=>ConvOuput_0);
   Ssave : saveState port map ( DMAOutput(15)=>nx10314, DMAOutput(14)=>
      nx10318, DMAOutput(13)=>nx10322, DMAOutput(12)=>nx10326, DMAOutput(11)
      =>nx10330, DMAOutput(10)=>nx10334, DMAOutput(9)=>nx10338, DMAOutput(8)
      =>nx10342, DMAOutput(7)=>nx10346, DMAOutput(6)=>nx10350, DMAOutput(5)
      =>nx10354, DMAOutput(4)=>nx10358, DMAOutput(3)=>nx10362, DMAOutput(2)
      =>nx10366, DMAOutput(1)=>nx10370, DMAOutput(0)=>nx10374, 
      RegisterOutput(15)=>nx10396, RegisterOutput(14)=>ConvOuput_14, 
      RegisterOutput(13)=>ConvOuput_13, RegisterOutput(12)=>ConvOuput_12, 
      RegisterOutput(11)=>ConvOuput_11, RegisterOutput(10)=>ConvOuput_10, 
      RegisterOutput(9)=>ConvOuput_9, RegisterOutput(8)=>ConvOuput_8, 
      RegisterOutput(7)=>ConvOuput_7, RegisterOutput(6)=>ConvOuput_6, 
      RegisterOutput(5)=>ConvOuput_5, RegisterOutput(4)=>ConvOuput_4, 
      RegisterOutput(3)=>ConvOuput_3, RegisterOutput(2)=>ConvOuput_2, 
      RegisterOutput(1)=>ConvOuput_1, RegisterOutput(0)=>ConvOuput_0, 
      bias1(15)=>Bias0_15, bias1(14)=>Bias0_14, bias1(13)=>Bias0_13, 
      bias1(12)=>Bias0_12, bias1(11)=>Bias0_11, bias1(10)=>Bias0_10, 
      bias1(9)=>Bias0_9, bias1(8)=>Bias0_8, bias1(7)=>Bias0_7, bias1(6)=>
      Bias0_6, bias1(5)=>Bias0_5, bias1(4)=>Bias0_4, bias1(3)=>Bias0_3, 
      bias1(2)=>Bias0_2, bias1(1)=>Bias0_1, bias1(0)=>Bias0_0, bias2(15)=>
      Bias1_15, bias2(14)=>Bias1_14, bias2(13)=>Bias1_13, bias2(12)=>
      Bias1_12, bias2(11)=>Bias1_11, bias2(10)=>Bias1_10, bias2(9)=>Bias1_9, 
      bias2(8)=>Bias1_8, bias2(7)=>Bias1_7, bias2(6)=>Bias1_6, bias2(5)=>
      Bias1_5, bias2(4)=>Bias1_4, bias2(3)=>Bias1_3, bias2(2)=>Bias1_2, 
      bias2(1)=>Bias1_1, bias2(0)=>Bias1_0, bias3(15)=>Bias2_15, bias3(14)=>
      Bias2_14, bias3(13)=>Bias2_13, bias3(12)=>Bias2_12, bias3(11)=>
      Bias2_11, bias3(10)=>Bias2_10, bias3(9)=>Bias2_9, bias3(8)=>Bias2_8, 
      bias3(7)=>Bias2_7, bias3(6)=>Bias2_6, bias3(5)=>Bias2_5, bias3(4)=>
      Bias2_4, bias3(3)=>Bias2_3, bias3(2)=>Bias2_2, bias3(1)=>Bias2_1, 
      bias3(0)=>Bias2_0, bias4(15)=>Bias3_15, bias4(14)=>Bias3_14, bias4(13)
      =>Bias3_13, bias4(12)=>Bias3_12, bias4(11)=>Bias3_11, bias4(10)=>
      Bias3_10, bias4(9)=>Bias3_9, bias4(8)=>Bias3_8, bias4(7)=>Bias3_7, 
      bias4(6)=>Bias3_6, bias4(5)=>Bias3_5, bias4(4)=>Bias3_4, bias4(3)=>
      Bias3_3, bias4(2)=>Bias3_2, bias4(1)=>Bias3_1, bias4(0)=>Bias3_0, 
      bias5(15)=>Bias4_15, bias5(14)=>Bias4_14, bias5(13)=>Bias4_13, 
      bias5(12)=>Bias4_12, bias5(11)=>Bias4_11, bias5(10)=>Bias4_10, 
      bias5(9)=>Bias4_9, bias5(8)=>Bias4_8, bias5(7)=>Bias4_7, bias5(6)=>
      Bias4_6, bias5(5)=>Bias4_5, bias5(4)=>Bias4_4, bias5(3)=>Bias4_3, 
      bias5(2)=>Bias4_2, bias5(1)=>Bias4_1, bias5(0)=>Bias4_0, bias6(15)=>
      Bias5_15, bias6(14)=>Bias5_14, bias6(13)=>Bias5_13, bias6(12)=>
      Bias5_12, bias6(11)=>Bias5_11, bias6(10)=>Bias5_10, bias6(9)=>Bias5_9, 
      bias6(8)=>Bias5_8, bias6(7)=>Bias5_7, bias6(6)=>Bias5_6, bias6(5)=>
      Bias5_5, bias6(4)=>Bias5_4, bias6(3)=>Bias5_3, bias6(2)=>Bias5_2, 
      bias6(1)=>Bias5_1, bias6(0)=>Bias5_0, bias7(15)=>Bias6_15, bias7(14)=>
      Bias6_14, bias7(13)=>Bias6_13, bias7(12)=>Bias6_12, bias7(11)=>
      Bias6_11, bias7(10)=>Bias6_10, bias7(9)=>Bias6_9, bias7(8)=>Bias6_8, 
      bias7(7)=>Bias6_7, bias7(6)=>Bias6_6, bias7(5)=>Bias6_5, bias7(4)=>
      Bias6_4, bias7(3)=>Bias6_3, bias7(2)=>Bias6_2, bias7(1)=>Bias6_1, 
      bias7(0)=>Bias6_0, bias8(15)=>Bias7_15, bias8(14)=>Bias7_14, bias8(13)
      =>Bias7_13, bias8(12)=>Bias7_12, bias8(11)=>Bias7_11, bias8(10)=>
      Bias7_10, bias8(9)=>Bias7_9, bias8(8)=>Bias7_8, bias8(7)=>Bias7_7, 
      bias8(6)=>Bias7_6, bias8(5)=>Bias7_5, bias8(4)=>Bias7_4, bias8(3)=>
      Bias7_3, bias8(2)=>Bias7_2, bias8(1)=>Bias7_1, bias8(0)=>Bias7_0, 
      Depth(3)=>nx10406, Depth(2)=>nx10408, Depth(1)=>nx10410, Depth(0)=>
      nx10412, NumberOfFiltersCounter(3)=>nx10398, NumberOfFiltersCounter(2)
      =>nx10400, NumberOfFiltersCounter(1)=>nx10402, 
      NumberOfFiltersCounter(0)=>nx10404, rst=>rst, stateinput(14)=>zero_11, 
      stateinput(13)=>nx9950, stateinput(12)=>nx9954, stateinput(11)=>
      zero_11, stateinput(10)=>current_state_10, stateinput(9)=>nx9958, 
      stateinput(8)=>current_state_8, stateinput(7)=>zero_11, stateinput(6)
      =>zero_11, stateinput(5)=>zero_11, stateinput(4)=>zero_11, 
      stateinput(3)=>zero_11, stateinput(2)=>zero_11, stateinput(1)=>zero_11, 
      stateinput(0)=>zero_11, clk=>nx10424, outputCounterToDma(12)=>
      AddressI_12, outputCounterToDma(11)=>AddressI_11, 
      outputCounterToDma(10)=>AddressI_10, outputCounterToDma(9)=>AddressI_9, 
      outputCounterToDma(8)=>AddressI_8, outputCounterToDma(7)=>AddressI_7, 
      outputCounterToDma(6)=>AddressI_6, outputCounterToDma(5)=>AddressI_5, 
      outputCounterToDma(4)=>AddressI_4, outputCounterToDma(3)=>AddressI_3, 
      outputCounterToDma(2)=>AddressI_2, outputCounterToDma(1)=>AddressI_1, 
      outputCounterToDma(0)=>AddressI_0, RealOutputCounter(12)=>
      RealOutputCounter_12, RealOutputCounter(11)=>RealOutputCounter_11, 
      RealOutputCounter(10)=>RealOutputCounter_10, RealOutputCounter(9)=>
      RealOutputCounter_9, RealOutputCounter(8)=>RealOutputCounter_8, 
      RealOutputCounter(7)=>RealOutputCounter_7, RealOutputCounter(6)=>
      RealOutputCounter_6, RealOutputCounter(5)=>RealOutputCounter_5, 
      RealOutputCounter(4)=>RealOutputCounter_4, RealOutputCounter(3)=>
      RealOutputCounter_3, RealOutputCounter(2)=>RealOutputCounter_2, 
      RealOutputCounter(1)=>RealOutputCounter_1, RealOutputCounter(0)=>
      RealOutputCounter_0, output(15)=>DataIIn_15, output(14)=>DataIIn_14, 
      output(13)=>DataIIn_13, output(12)=>DataIIn_12, output(11)=>DataIIn_11, 
      output(10)=>DataIIn_10, output(9)=>DataIIn_9, output(8)=>DataIIn_8, 
      output(7)=>DataIIn_7, output(6)=>DataIIn_6, output(5)=>DataIIn_5, 
      output(4)=>DataIIn_4, output(3)=>DataIIn_3, output(2)=>DataIIn_2, 
      output(1)=>DataIIn_1, output(0)=>DataIIn_0, ShiftLeftCounterOutput(4)
      =>ShiftLeftCounterOutput_4, ShiftLeftCounterOutput(3)=>
      ShiftLeftCounterOutput_3, ShiftLeftCounterOutput(2)=>
      ShiftLeftCounterOutput_2, ShiftLeftCounterOutput(1)=>
      ShiftLeftCounterOutput_1, ShiftLeftCounterOutput(0)=>
      ShiftLeftCounterOutput_0, ShiftCounterRst=>ShiftCounterRst, 
      AddresCounterLoad(12)=>OutputCounterLoad_12, AddresCounterLoad(11)=>
      OutputCounterLoad_11, AddresCounterLoad(10)=>OutputCounterLoad_10, 
      AddresCounterLoad(9)=>OutputCounterLoad_9, AddresCounterLoad(8)=>
      OutputCounterLoad_8, AddresCounterLoad(7)=>OutputCounterLoad_7, 
      AddresCounterLoad(6)=>OutputCounterLoad_6, AddresCounterLoad(5)=>
      OutputCounterLoad_5, AddresCounterLoad(4)=>OutputCounterLoad_4, 
      AddresCounterLoad(3)=>OutputCounterLoad_3, AddresCounterLoad(2)=>
      OutputCounterLoad_2, AddresCounterLoad(1)=>OutputCounterLoad_1, 
      AddresCounterLoad(0)=>OutputCounterLoad_0, X=>X, Y=>Y);
   Istate : ImageState port map ( current_state(14)=>zero_11, 
      current_state(13)=>nx9950, current_state(12)=>nx9954, 
      current_state(11)=>current_state_11, current_state(10)=>zero_11, 
      current_state(9)=>nx9958, current_state(8)=>zero_11, current_state(7)
      =>zero_11, current_state(6)=>zero_11, current_state(5)=>zero_11, 
      current_state(4)=>zero_11, current_state(3)=>zero_11, current_state(2)
      =>zero_11, current_state(1)=>zero_11, current_state(0)=>zero_11, 
      WSquared(9)=>WidthSquareOut_9, WSquared(8)=>WidthSquareOut_8, 
      WSquared(7)=>WidthSquareOut_7, WSquared(6)=>WidthSquareOut_6, 
      WSquared(5)=>WidthSquareOut_5, WSquared(4)=>WidthSquareOut_4, 
      WSquared(3)=>WidthSquareOut_3, WSquared(2)=>WidthSquareOut_2, 
      WSquared(1)=>WidthSquareOut_1, WSquared(0)=>WidthSquareOut_0, 
      AddresCounterIN(12)=>RealOutputCounter_12, AddresCounterIN(11)=>
      RealOutputCounter_11, AddresCounterIN(10)=>RealOutputCounter_10, 
      AddresCounterIN(9)=>RealOutputCounter_9, AddresCounterIN(8)=>
      RealOutputCounter_8, AddresCounterIN(7)=>RealOutputCounter_7, 
      AddresCounterIN(6)=>RealOutputCounter_6, AddresCounterIN(5)=>
      RealOutputCounter_5, AddresCounterIN(4)=>RealOutputCounter_4, 
      AddresCounterIN(3)=>RealOutputCounter_3, AddresCounterIN(2)=>
      RealOutputCounter_2, AddresCounterIN(1)=>RealOutputCounter_1, 
      AddresCounterIN(0)=>RealOutputCounter_0, AddresCounterLoad(12)=>
      OutputCounterLoad_12, AddresCounterLoad(11)=>OutputCounterLoad_11, 
      AddresCounterLoad(10)=>OutputCounterLoad_10, AddresCounterLoad(9)=>
      OutputCounterLoad_9, AddresCounterLoad(8)=>OutputCounterLoad_8, 
      AddresCounterLoad(7)=>OutputCounterLoad_7, AddresCounterLoad(6)=>
      OutputCounterLoad_6, AddresCounterLoad(5)=>OutputCounterLoad_5, 
      AddresCounterLoad(4)=>OutputCounterLoad_4, AddresCounterLoad(3)=>
      OutputCounterLoad_3, AddresCounterLoad(2)=>OutputCounterLoad_2, 
      AddresCounterLoad(1)=>OutputCounterLoad_1, AddresCounterLoad(0)=>
      OutputCounterLoad_0, NoOfShiftsCounter(4)=>ShiftLeftCounterOutput_4, 
      NoOfShiftsCounter(3)=>ShiftLeftCounterOutput_3, NoOfShiftsCounter(2)=>
      ShiftLeftCounterOutput_2, NoOfShiftsCounter(1)=>
      ShiftLeftCounterOutput_1, NoOfShiftsCounter(0)=>
      ShiftLeftCounterOutput_0, LayerInfoIn(15)=>zero_11, LayerInfoIn(14)=>
      zero_11, LayerInfoIn(13)=>zero_11, LayerInfoIn(12)=>zero_11, 
      LayerInfoIn(11)=>zero_11, LayerInfoIn(10)=>zero_11, LayerInfoIn(9)=>
      zero_11, LayerInfoIn(8)=>nx10378, LayerInfoIn(7)=>nx10382, 
      LayerInfoIn(6)=>nx10386, LayerInfoIn(5)=>nx10388, LayerInfoIn(4)=>
      nx10392, LayerInfoIn(3)=>LayerInfoOut_3, LayerInfoIn(2)=>
      LayerInfoOut_2, LayerInfoIn(1)=>LayerInfoOut_1, LayerInfoIn(0)=>
      LayerInfoOut_0, CLK=>nx10426, RST=>rst, Q=>Q, NumOfFilters(3)=>
      NumOfFilters_3, NumOfFilters(2)=>NumOfFilters_2, NumOfFilters(1)=>
      NumOfFilters_1, NumOfFilters(0)=>NumOfFilters_0, NumOfHeight(4)=>
      NumOfHeight_4, NumOfHeight(3)=>NumOfHeight_3, NumOfHeight(2)=>
      NumOfHeight_2, NumOfHeight(1)=>NumOfHeight_1, NumOfHeight(0)=>
      NumOfHeight_0, X1=>X, Y1=>Y, K1=>K);
   ChState : StateChecks port map ( current_state(14)=>zero_11, 
      current_state(13)=>nx9950, current_state(12)=>nx9956, 
      current_state(11)=>zero_11, current_state(10)=>zero_11, 
      current_state(9)=>zero_11, current_state(8)=>zero_11, current_state(7)
      =>zero_11, current_state(6)=>zero_11, current_state(5)=>zero_11, 
      current_state(4)=>zero_11, current_state(3)=>zero_11, current_state(2)
      =>zero_11, current_state(1)=>zero_11, current_state(0)=>zero_11, 
      noOfLayers(15)=>zero_11, noOfLayers(14)=>zero_11, noOfLayers(13)=>
      zero_11, noOfLayers(12)=>zero_11, noOfLayers(11)=>zero_11, 
      noOfLayers(10)=>zero_11, noOfLayers(9)=>zero_11, noOfLayers(8)=>
      zero_11, noOfLayers(7)=>zero_11, noOfLayers(6)=>zero_11, noOfLayers(5)
      =>zero_11, noOfLayers(4)=>zero_11, noOfLayers(3)=>zero_11, 
      noOfLayers(2)=>zero_11, noOfLayers(1)=>NoOfLayers_1, noOfLayers(0)=>
      NoOfLayers_0, LayerInfo(15)=>zero_11, LayerInfo(14)=>zero_11, 
      LayerInfo(13)=>zero_11, LayerInfo(12)=>LayerInfoOut_12, LayerInfo(11)
      =>LayerInfoOut_11, LayerInfo(10)=>LayerInfoOut_10, LayerInfo(9)=>
      LayerInfoOut_9, LayerInfo(8)=>zero_11, LayerInfo(7)=>zero_11, 
      LayerInfo(6)=>zero_11, LayerInfo(5)=>zero_11, LayerInfo(4)=>zero_11, 
      LayerInfo(3)=>zero_11, LayerInfo(2)=>zero_11, LayerInfo(1)=>zero_11, 
      LayerInfo(0)=>zero_11, CLK=>zero_11, RST=>rst, L=>L, D=>D, 
      CNDoutput(3)=>CNDepthoutput_3, CNDoutput(2)=>CNDepthoutput_2, 
      CNDoutput(1)=>CNDepthoutput_1, CNDoutput(0)=>CNDepthoutput_0, 
      CNLoutput(1)=>DANGLING(2727), CNLoutput(0)=>DANGLING(2728));
   Owidth : outWidthState port map ( currentState(14)=>zero_11, 
      currentState(13)=>nx9950, currentState(12)=>zero_11, currentState(11)
      =>zero_11, currentState(10)=>zero_11, currentState(9)=>zero_11, 
      currentState(8)=>zero_11, currentState(7)=>zero_11, currentState(6)=>
      zero_11, currentState(5)=>zero_11, currentState(4)=>zero_11, 
      currentState(3)=>zero_11, currentState(2)=>zero_11, currentState(1)=>
      zero_11, currentState(0)=>zero_11, infoReg(15)=>zero_11, infoReg(14)=>
      zero_11, infoReg(13)=>zero_11, infoReg(12)=>zero_11, infoReg(11)=>
      zero_11, infoReg(10)=>zero_11, infoReg(9)=>zero_11, infoReg(8)=>
      nx10378, infoReg(7)=>nx10382, infoReg(6)=>nx10386, infoReg(5)=>nx10388, 
      infoReg(4)=>nx10392, infoReg(3)=>zero_11, infoReg(2)=>zero_11, 
      infoReg(1)=>zero_11, infoReg(0)=>zero_11, address(12)=>AddressI_12, 
      address(11)=>AddressI_11, address(10)=>AddressI_10, address(9)=>
      AddressI_9, address(8)=>AddressI_8, address(7)=>AddressI_7, address(6)
      =>AddressI_6, address(5)=>AddressI_5, address(4)=>AddressI_4, 
      address(3)=>AddressI_3, address(2)=>AddressI_2, address(1)=>AddressI_1, 
      address(0)=>AddressI_0, outWidth(15)=>DataIIn_15, outWidth(14)=>
      DataIIn_14, outWidth(13)=>DataIIn_13, outWidth(12)=>DataIIn_12, 
      outWidth(11)=>DataIIn_11, outWidth(10)=>DataIIn_10, outWidth(9)=>
      DataIIn_9, outWidth(8)=>DataIIn_8, outWidth(7)=>DataIIn_7, outWidth(6)
      =>DataIIn_6, outWidth(5)=>DataIIn_5, outWidth(4)=>DataIIn_4, 
      outWidth(3)=>DataIIn_3, outWidth(2)=>DataIIn_2, outWidth(1)=>DataIIn_1, 
      outWidth(0)=>DataIIn_0);
   ix9649 : fake_vcc port map ( Y=>PWR);
   ix9647 : fake_gnd port map ( Y=>zero_11);
   ix399 : or02 port map ( Y=>ramSelector, A0=>current_state_8, A1=>nx9950);
   reg_current_state_8 : dffr port map ( Q=>current_state_8, QB=>OPEN, D=>
      next_state_8, CLK=>nx10430, R=>rst);
   lat_next_state_8 : latch port map ( Q=>next_state_8, D=>nx9962, CLK=>
      nx10434);
   reg_current_state_7 : dffr port map ( Q=>OPEN, QB=>nx9870, D=>
      next_state_7, CLK=>nx10428, R=>rst);
   lat_next_state_7 : latch port map ( Q=>next_state_7, D=>nx154, CLK=>
      nx10434);
   ix155 : nand02 port map ( Y=>nx154, A0=>nx9760, A1=>nx9814);
   ix9761 : aoi22 port map ( Y=>nx9760, A0=>K, A1=>current_state_11, B0=>X, 
      B1=>nx9960);
   reg_current_state_11 : dffr port map ( Q=>current_state_11, QB=>OPEN, D=>
      next_state_11, CLK=>nx10426, R=>rst);
   lat_next_state_11 : latch port map ( Q=>next_state_11, D=>nx256, CLK=>
      nx10432);
   ix257 : nor03_2x port map ( Y=>nx256, A0=>nx9765, A1=>Y, A2=>nx9768);
   ix9766 : nand04 port map ( Y=>nx9765, A0=>ShiftLeftCounterOutput_2, A1=>
      ShiftLeftCounterOutput_4, A2=>ShiftLeftCounterOutput_3, A3=>nx18);
   ix19 : nor02_2x port map ( Y=>nx18, A0=>ShiftLeftCounterOutput_1, A1=>
      ShiftLeftCounterOutput_0);
   lat_next_state_10 : latch port map ( Q=>next_state_10, D=>nx240, CLK=>
      nx10432);
   reg_current_state_9 : dffr port map ( Q=>current_state_9, QB=>OPEN, D=>
      next_state_9, CLK=>nx10426, R=>rst);
   lat_next_state_9 : latch port map ( Q=>next_state_9, D=>nx224, CLK=>
      nx10432);
   ix225 : and02 port map ( Y=>nx224, A0=>next_state_dup_124, A1=>
      current_state_8);
   reg_next_state_dup_124 : dff port map ( Q=>next_state_dup_124, QB=>OPEN, 
      D=>nx9738, CLK=>nx10028);
   ix9739 : or02 port map ( Y=>nx9738, A0=>next_state_dup_124, A1=>WriteI);
   ix217 : nand02 port map ( Y=>WriteI, A0=>nx9780, A1=>nx9792);
   ix9781 : oai21 port map ( Y=>nx9780, A0=>nx210, A1=>SaveAckLatch, B0=>
      current_state_8);
   ix211 : nor04 port map ( Y=>nx210, A0=>nx10406, A1=>nx10408, A2=>nx10410, 
      A3=>nx10412);
   ix9064 : dffr port map ( Q=>nx9063, QB=>OPEN, D=>PWR, CLK=>nx10436, R=>
      nx180);
   ix9786 : nand02 port map ( Y=>NOT_nx0, A0=>start, A1=>cl);
   ix181 : nand02 port map ( Y=>nx180, A0=>current_state_8, A1=>nx10026);
   lat_next_state_13 : latch port map ( Q=>next_state_13, D=>nx9711, CLK=>
      nx10432);
   ix289 : aoi21 port map ( Y=>nx9711, A0=>L, A1=>D, B0=>nx9796);
   reg_current_state_12 : dffr port map ( Q=>OPEN, QB=>nx9796, D=>
      next_state_12, CLK=>nx10426, R=>rst);
   lat_next_state_12 : latch port map ( Q=>next_state_12, D=>nx270, CLK=>
      nx10432);
   ix271 : nor02ii port map ( Y=>nx270, A0=>K, A1=>current_state_11);
   reg_current_state_14 : dffr port map ( Q=>done_EXMPLR, QB=>OPEN, D=>
      next_state_14, CLK=>nx10420, R=>rst);
   lat_next_state_14 : latch port map ( Q=>next_state_14, D=>nx300, CLK=>
      nx10432);
   reg_next_state_dup_134 : dff port map ( Q=>next_state_dup_134, QB=>OPEN, 
      D=>NOT_L, CLK=>nx10028);
   ix9806 : inv01 port map ( Y=>NOT_L, A=>L);
   reg_current_state_13 : dffr port map ( Q=>OPEN, QB=>nx9792, D=>
      next_state_13, CLK=>nx10418, R=>rst);
   reg_current_state_10 : dffr port map ( Q=>current_state_10, QB=>nx9768, D
      =>next_state_10, CLK=>nx10426, R=>rst);
   ix9815 : aoi32 port map ( Y=>nx9814, A0=>nx20, A1=>Y, A2=>
      current_state_10, B0=>next_state_dup_96, B1=>nx142);
   reg_next_state_dup_96 : dff port map ( Q=>next_state_dup_96, QB=>OPEN, D
      =>nx9718, CLK=>nx10028);
   ix9719 : or02 port map ( Y=>nx9718, A0=>next_state_dup_96, A1=>nx48);
   ix49 : aoi21 port map ( Y=>nx48, A0=>nx9822, A1=>nx9826, B0=>
      ImgCounterOuput_0);
   ix9823 : nand03 port map ( Y=>nx9822, A0=>nx10500, A1=>ImgCounterOuput_2, 
      A2=>nx9824);
   ix9825 : inv01 port map ( Y=>nx9824, A=>ImgCounterOuput_1);
   ix9827 : or03 port map ( Y=>nx9826, A0=>nx10502, A1=>ImgCounterOuput_2, 
      A2=>nx9824);
   reg_current_state_3 : dffr port map ( Q=>current_state_3, QB=>OPEN, D=>
      next_state_3, CLK=>nx10428, R=>rst);
   lat_next_state_3 : latch port map ( Q=>next_state_3, D=>nx130, CLK=>
      nx10434);
   ix131 : nand02 port map ( Y=>nx130, A0=>nx9833, A1=>nx9835);
   ix9834 : nand04 port map ( Y=>nx9833, A0=>nx9954, A1=>L, A2=>D, A3=>
      LayerInfoOut_15);
   reg_current_state_2 : dffr port map ( Q=>current_state_2, QB=>nx9835, D=>
      next_state_2, CLK=>nx10428, R=>rst);
   lat_next_state_2 : latch port map ( Q=>next_state_2, D=>nx112, CLK=>
      nx10434);
   reg_next_state_dup_26 : dff port map ( Q=>next_state_dup_26, QB=>OPEN, D
      =>nx9728, CLK=>nx10436);
   ix9729 : mux21_ni port map ( Y=>nx9728, A0=>next_state_dup_26, A1=>
      nx10304, S0=>nx10308);
   reg_current_state_1 : dffr port map ( Q=>OPEN, QB=>nx9849, D=>
      next_state_1, CLK=>nx10428, R=>rst);
   lat_next_state_1 : latch port map ( Q=>next_state_1, D=>nx100, CLK=>
      nx10432);
   ix101 : ao21 port map ( Y=>nx100, A0=>next_state_dup_147, A1=>nx9950, B0
      =>current_state_0);
   reg_next_state_dup_147 : dff port map ( Q=>next_state_dup_147, QB=>OPEN, 
      D=>L, CLK=>nx10028);
   reg_current_state_0 : dffs_ni port map ( Q=>current_state_0, QB=>OPEN, D
      =>zero_11, CLK=>nx10426, S=>rst);
   reg_current_state_6 : dffr port map ( Q=>current_state_6, QB=>OPEN, D=>
      next_state_6, CLK=>nx10428, R=>rst);
   lat_next_state_6 : latch port map ( Q=>next_state_6, D=>nx66, CLK=>
      nx10434);
   ix67 : nand02 port map ( Y=>nx66, A0=>nx9854, A1=>nx9858);
   ix9855 : nand04 port map ( Y=>nx9854, A0=>nx9954, A1=>L, A2=>D, A3=>
      nx9856);
   ix9857 : inv01 port map ( Y=>nx9856, A=>LayerInfoOut_15);
   reg_current_state_5 : dffr port map ( Q=>current_state_5, QB=>nx9858, D=>
      next_state_5, CLK=>nx10428, R=>rst);
   lat_next_state_5 : latch port map ( Q=>next_state_5, D=>nx9966, CLK=>
      nx10434);
   reg_current_state_4 : dffr port map ( Q=>current_state_4, QB=>OPEN, D=>
      next_state_4, CLK=>nx10428, R=>rst);
   lat_next_state_4 : latch port map ( Q=>next_state_4, D=>nx322, CLK=>
      nx10434);
   reg_next_state_dup_24 : dff port map ( Q=>next_state_dup_24, QB=>nx9866, 
      D=>nx9748, CLK=>nx10436);
   ix401 : or02 port map ( Y=>ImgAddRST, A0=>nx9952, A1=>rst);
   ix403 : or02 port map ( Y=>TriChnagerToaddEN, A0=>current_state_6, A1=>
      current_state_10);
   ix455 : oai21 port map ( Y=>AddressChangerEN, A0=>nx9875, A1=>nx9883, B0
      =>nx9893);
   ix9876 : nand04 port map ( Y=>nx9875, A0=>DontRstIndicator, A1=>nx9960, 
      A2=>nx418, A3=>nx9881);
   ix419 : or02 port map ( Y=>nx418, A0=>nx416, A1=>lastFilter);
   ix417 : nor04 port map ( Y=>nx416, A0=>nx9879, A1=>LayerInfoOut_3, A2=>
      LayerInfoOut_2, A3=>LayerInfoOut_1);
   ix9880 : inv01 port map ( Y=>nx9879, A=>LayerInfoOut_0);
   ix9882 : xnor2 port map ( Y=>nx9881, A0=>ShiftLeftCounterOutput_4, A1=>
      nx10378);
   ix9884 : nand04 port map ( Y=>nx9883, A0=>nx9885, A1=>nx9887, A2=>nx9889, 
      A3=>nx9891);
   ix9886 : xnor2 port map ( Y=>nx9885, A0=>ShiftLeftCounterOutput_0, A1=>
      nx10392);
   ix9888 : xnor2 port map ( Y=>nx9887, A0=>ShiftLeftCounterOutput_1, A1=>
      nx10388);
   ix9890 : xnor2 port map ( Y=>nx9889, A0=>ShiftLeftCounterOutput_2, A1=>
      nx10386);
   ix9892 : xnor2 port map ( Y=>nx9891, A0=>ShiftLeftCounterOutput_3, A1=>
      nx10382);
   ix9894 : nand02 port map ( Y=>nx9893, A0=>nx10310, A1=>nx9966);
   ix461 : or03 port map ( Y=>ShiftCounterRst, A0=>nx456, A1=>
      current_state_11, A2=>rst);
   ix469 : and02 port map ( Y=>ImgAddRegEN, A0=>nx10028, A1=>nx466);
   ix467 : nand04 port map ( Y=>nx466, A0=>nx9899, A1=>nx9903, A2=>nx9905, 
      A3=>nx9849);
   ix9900 : aoi21 port map ( Y=>nx9899, A0=>nx9901, A1=>nx9964, B0=>
      current_state_2);
   ix9902 : inv01 port map ( Y=>nx9901, A=>IndicatorI_0);
   ix9904 : nor02_2x port map ( Y=>nx9903, A0=>current_state_3, A1=>
      current_state_6);
   ix517 : aoi21 port map ( Y=>FilterAddressEN, A0=>nx9908, A1=>nx9913, B0=>
      LayerInfoOut_15);
   ix9909 : aoi21 port map ( Y=>nx9908, A0=>lastFilter, A1=>current_state_6, 
      B0=>TriStateCounterEN);
   ix507 : inv01 port map ( Y=>TriStateCounterEN, A=>nx9911);
   ix9912 : oai21 port map ( Y=>nx9911, A0=>current_state_0, A1=>nx9972, B0
      =>nx10310);
   ix9914 : aoi32 port map ( Y=>nx9913, A0=>nx494, A1=>current_state_10, A2
      =>nx418, B0=>nx10310, B1=>nx350);
   ix495 : oai21 port map ( Y=>nx494, A0=>DontRstIndicator, A1=>nx9916, B0=>
      lastDepthOut);
   ix9917 : nor03_2x port map ( Y=>nx9916, A0=>nx482, A1=>nx480, A2=>nx478);
   ix483 : xor2 port map ( Y=>nx482, A0=>NumOfHeight_3, A1=>nx10382);
   ix481 : xor2 port map ( Y=>nx480, A0=>NumOfHeight_2, A1=>nx10386);
   ix479 : nand03 port map ( Y=>nx478, A0=>nx9921, A1=>nx9923, A2=>nx9925);
   ix9922 : xnor2 port map ( Y=>nx9921, A0=>NumOfHeight_0, A1=>nx10394);
   ix9924 : xnor2 port map ( Y=>nx9923, A0=>NumOfHeight_4, A1=>nx10378);
   ix9926 : xnor2 port map ( Y=>nx9925, A0=>NumOfHeight_1, A1=>nx10390);
   ix351 : oai21 port map ( Y=>nx350, A0=>IndicatorF_0, A1=>nx9870, B0=>
      nx9905);
   ix9930 : inv01 port map ( Y=>SwitchBar_0, A=>SwitchMEM_0);
   ix397 : nand04 port map ( Y=>ReadI, A0=>nx9932, A1=>nx9934, A2=>nx9899, 
      A3=>nx9903);
   ix9933 : nor03_2x port map ( Y=>nx9932, A0=>nx9966, A1=>current_state_5, 
      A2=>nx9972);
   ix9935 : nand03 port map ( Y=>nx9934, A0=>nx382, A1=>current_state_8, A2
      =>nx9941);
   ix383 : mux21 port map ( Y=>nx382, A0=>nx9937, A1=>nx9939, S0=>nx10406);
   ix9938 : nor03_2x port map ( Y=>nx9937, A0=>nx10410, A1=>nx10408, A2=>
      nx10412);
   ix9940 : and03 port map ( Y=>nx9939, A0=>nx10410, A1=>nx10408, A2=>
      nx10412);
   ix355 : or03 port map ( Y=>ReadF, A0=>current_state_0, A1=>nx9972, A2=>
      nx350);
   tri_dmaStartSignal : tri01 port map ( Y=>dmaStartSignal, A=>PWR, E=>
      zero_11);
   ix143 : inv01 port map ( Y=>nx142, A=>nx9903);
   ix21 : inv01 port map ( Y=>nx20, A=>nx9765);
   ix1 : inv01 port map ( Y=>CLK, A=>NOT_nx0);
   ix9949 : inv01 port map ( Y=>nx9950, A=>nx9792);
   ix9951 : inv01 port map ( Y=>nx9952, A=>nx9792);
   ix9953 : inv01 port map ( Y=>nx9954, A=>nx9796);
   ix9955 : inv01 port map ( Y=>nx9956, A=>nx9796);
   ix9957 : buf02 port map ( Y=>nx9958, A=>current_state_9);
   ix9959 : buf02 port map ( Y=>nx9960, A=>current_state_9);
   ix9961 : inv01 port map ( Y=>nx9962, A=>nx9870);
   ix9963 : inv01 port map ( Y=>nx9964, A=>nx9870);
   ix9965 : buf02 port map ( Y=>nx9966, A=>current_state_4);
   ix9967 : buf02 port map ( Y=>nx9968, A=>current_state_4);
   ix9969 : inv02 port map ( Y=>nx9970, A=>nx9849);
   ix9971 : inv02 port map ( Y=>nx9972, A=>nx9849);
   ix9973 : buf02 port map ( Y=>nx9974, A=>FilterAddressOut_12);
   ix9975 : buf02 port map ( Y=>nx9976, A=>FilterAddressOut_12);
   ix9977 : buf02 port map ( Y=>nx9978, A=>FilterAddressOut_11);
   ix9979 : buf02 port map ( Y=>nx9980, A=>FilterAddressOut_11);
   ix9981 : buf02 port map ( Y=>nx9982, A=>FilterAddressOut_10);
   ix9983 : buf02 port map ( Y=>nx9984, A=>FilterAddressOut_10);
   ix9985 : buf02 port map ( Y=>nx9986, A=>FilterAddressOut_9);
   ix9987 : buf02 port map ( Y=>nx9988, A=>FilterAddressOut_9);
   ix9989 : buf02 port map ( Y=>nx9990, A=>FilterAddressOut_8);
   ix9991 : buf02 port map ( Y=>nx9992, A=>FilterAddressOut_8);
   ix9993 : buf02 port map ( Y=>nx9994, A=>FilterAddressOut_7);
   ix9995 : buf02 port map ( Y=>nx9996, A=>FilterAddressOut_7);
   ix9997 : buf02 port map ( Y=>nx9998, A=>FilterAddressOut_6);
   ix9999 : buf02 port map ( Y=>nx10000, A=>FilterAddressOut_6);
   ix10001 : buf02 port map ( Y=>nx10002, A=>FilterAddressOut_5);
   ix10003 : buf02 port map ( Y=>nx10004, A=>FilterAddressOut_5);
   ix10005 : buf02 port map ( Y=>nx10006, A=>FilterAddressOut_4);
   ix10007 : buf02 port map ( Y=>nx10008, A=>FilterAddressOut_4);
   ix10009 : buf02 port map ( Y=>nx10010, A=>FilterAddressOut_3);
   ix10011 : buf02 port map ( Y=>nx10012, A=>FilterAddressOut_3);
   ix10013 : buf02 port map ( Y=>nx10014, A=>FilterAddressOut_2);
   ix10015 : buf02 port map ( Y=>nx10016, A=>FilterAddressOut_2);
   ix10017 : buf02 port map ( Y=>nx10018, A=>FilterAddressOut_1);
   ix10019 : buf02 port map ( Y=>nx10020, A=>FilterAddressOut_1);
   ix10021 : buf02 port map ( Y=>nx10022, A=>FilterAddressOut_0);
   ix10023 : buf02 port map ( Y=>nx10024, A=>FilterAddressOut_0);
   ix10025 : buf02 port map ( Y=>nx10026, A=>ImgAddACKTriIN_0);
   ix10027 : buf02 port map ( Y=>nx10028, A=>ImgAddACKTriIN_0);
   ix10031 : inv02 port map ( Y=>nx10032, A=>nx10490);
   ix10033 : inv02 port map ( Y=>nx10034, A=>nx10490);
   ix10035 : inv02 port map ( Y=>nx10036, A=>nx10490);
   ix10037 : inv02 port map ( Y=>nx10038, A=>nx10490);
   ix10039 : inv02 port map ( Y=>nx10040, A=>nx10490);
   ix10041 : inv02 port map ( Y=>nx10042, A=>nx10490);
   ix10043 : inv02 port map ( Y=>nx10044, A=>nx10490);
   ix10045 : inv02 port map ( Y=>nx10046, A=>nx10442);
   ix10047 : inv02 port map ( Y=>nx10048, A=>nx10442);
   ix10049 : inv02 port map ( Y=>nx10050, A=>nx10442);
   ix10051 : inv02 port map ( Y=>nx10052, A=>nx10442);
   ix10053 : inv02 port map ( Y=>nx10054, A=>nx10442);
   ix10055 : inv02 port map ( Y=>nx10056, A=>nx10442);
   ix10057 : inv02 port map ( Y=>nx10058, A=>nx10442);
   ix10059 : inv02 port map ( Y=>nx10060, A=>nx10444);
   ix10061 : inv02 port map ( Y=>nx10062, A=>nx10444);
   ix10063 : inv02 port map ( Y=>nx10064, A=>nx10444);
   ix10065 : inv02 port map ( Y=>nx10066, A=>nx10444);
   ix10067 : inv02 port map ( Y=>nx10068, A=>nx10444);
   ix10069 : inv02 port map ( Y=>nx10070, A=>nx10444);
   ix10071 : inv02 port map ( Y=>nx10072, A=>nx10444);
   ix10073 : inv02 port map ( Y=>nx10074, A=>nx10446);
   ix10075 : inv02 port map ( Y=>nx10076, A=>nx10446);
   ix10077 : inv02 port map ( Y=>nx10078, A=>nx10446);
   ix10079 : inv02 port map ( Y=>nx10080, A=>nx10446);
   ix10081 : inv02 port map ( Y=>nx10082, A=>nx10446);
   ix10083 : inv02 port map ( Y=>nx10084, A=>nx10446);
   ix10085 : inv02 port map ( Y=>nx10086, A=>nx10446);
   ix10087 : inv02 port map ( Y=>nx10088, A=>nx10448);
   ix10089 : inv02 port map ( Y=>nx10090, A=>nx10448);
   ix10091 : inv02 port map ( Y=>nx10092, A=>nx10448);
   ix10093 : inv02 port map ( Y=>nx10094, A=>nx10448);
   ix10095 : inv02 port map ( Y=>nx10096, A=>nx10448);
   ix10097 : inv02 port map ( Y=>nx10098, A=>nx10448);
   ix10099 : inv02 port map ( Y=>nx10100, A=>nx10448);
   ix10101 : inv02 port map ( Y=>nx10102, A=>nx10450);
   ix10103 : inv02 port map ( Y=>nx10104, A=>nx10450);
   ix10105 : inv02 port map ( Y=>nx10106, A=>nx10450);
   ix10107 : inv02 port map ( Y=>nx10108, A=>nx10450);
   ix10109 : inv02 port map ( Y=>nx10110, A=>nx10450);
   ix10111 : inv02 port map ( Y=>nx10112, A=>nx10450);
   ix10113 : inv02 port map ( Y=>nx10114, A=>nx10450);
   ix10115 : inv02 port map ( Y=>nx10116, A=>nx10452);
   ix10117 : inv02 port map ( Y=>nx10118, A=>nx10452);
   ix10119 : inv02 port map ( Y=>nx10120, A=>nx10452);
   ix10121 : inv02 port map ( Y=>nx10122, A=>nx10452);
   ix10123 : inv02 port map ( Y=>nx10124, A=>nx10452);
   ix10125 : inv02 port map ( Y=>nx10126, A=>nx10452);
   ix10127 : inv02 port map ( Y=>nx10128, A=>nx10452);
   ix10129 : inv02 port map ( Y=>nx10130, A=>nx10454);
   ix10131 : inv02 port map ( Y=>nx10132, A=>nx10454);
   ix10133 : inv02 port map ( Y=>nx10134, A=>nx10454);
   ix10135 : inv02 port map ( Y=>nx10136, A=>nx10454);
   ix10137 : inv02 port map ( Y=>nx10138, A=>nx10454);
   ix10139 : inv02 port map ( Y=>nx10140, A=>nx10454);
   ix10141 : inv02 port map ( Y=>nx10142, A=>nx10454);
   ix10143 : inv02 port map ( Y=>nx10144, A=>nx10456);
   ix10145 : inv02 port map ( Y=>nx10146, A=>nx10456);
   ix10147 : inv02 port map ( Y=>nx10148, A=>nx10456);
   ix10149 : inv02 port map ( Y=>nx10150, A=>nx10456);
   ix10151 : inv02 port map ( Y=>nx10152, A=>nx10456);
   ix10153 : inv02 port map ( Y=>nx10154, A=>nx10456);
   ix10155 : inv02 port map ( Y=>nx10156, A=>nx10456);
   ix10157 : inv02 port map ( Y=>nx10158, A=>nx10458);
   ix10159 : inv02 port map ( Y=>nx10160, A=>nx10458);
   ix10161 : inv02 port map ( Y=>nx10162, A=>nx10458);
   ix10163 : inv02 port map ( Y=>nx10164, A=>nx10458);
   ix10165 : inv02 port map ( Y=>nx10166, A=>nx10458);
   ix10167 : inv02 port map ( Y=>nx10168, A=>nx10458);
   ix10169 : inv02 port map ( Y=>nx10170, A=>nx10458);
   ix10171 : inv02 port map ( Y=>nx10172, A=>nx10460);
   ix10173 : inv02 port map ( Y=>nx10174, A=>nx10460);
   ix10175 : inv02 port map ( Y=>nx10176, A=>nx10460);
   ix10177 : inv02 port map ( Y=>nx10178, A=>nx10460);
   ix10179 : inv02 port map ( Y=>nx10180, A=>nx10460);
   ix10181 : inv02 port map ( Y=>nx10182, A=>nx10460);
   ix10183 : inv02 port map ( Y=>nx10184, A=>nx10460);
   ix10185 : inv02 port map ( Y=>nx10186, A=>nx10462);
   ix10187 : inv02 port map ( Y=>nx10188, A=>nx10462);
   ix10189 : inv02 port map ( Y=>nx10190, A=>nx10462);
   ix10191 : inv02 port map ( Y=>nx10192, A=>nx10462);
   ix10193 : inv02 port map ( Y=>nx10194, A=>nx10462);
   ix10195 : inv02 port map ( Y=>nx10196, A=>nx10462);
   ix10197 : inv02 port map ( Y=>nx10198, A=>nx10462);
   ix10199 : inv02 port map ( Y=>nx10200, A=>nx10464);
   ix10201 : inv02 port map ( Y=>nx10202, A=>nx10464);
   ix10203 : inv02 port map ( Y=>nx10204, A=>nx10464);
   ix10205 : inv02 port map ( Y=>nx10206, A=>nx10464);
   ix10207 : inv02 port map ( Y=>nx10208, A=>nx10464);
   ix10209 : inv02 port map ( Y=>nx10210, A=>nx10464);
   ix10211 : inv02 port map ( Y=>nx10212, A=>nx10464);
   ix10213 : inv02 port map ( Y=>nx10214, A=>nx10466);
   ix10215 : inv02 port map ( Y=>nx10216, A=>nx10466);
   ix10217 : inv02 port map ( Y=>nx10218, A=>nx10466);
   ix10219 : inv02 port map ( Y=>nx10220, A=>nx10466);
   ix10221 : inv02 port map ( Y=>nx10222, A=>nx10466);
   ix10223 : inv02 port map ( Y=>nx10224, A=>nx10466);
   ix10225 : inv02 port map ( Y=>nx10226, A=>nx10466);
   ix10227 : inv02 port map ( Y=>nx10228, A=>nx10468);
   ix10229 : inv02 port map ( Y=>nx10230, A=>nx10468);
   ix10231 : inv02 port map ( Y=>nx10232, A=>nx10468);
   ix10233 : inv02 port map ( Y=>nx10234, A=>nx10468);
   ix10235 : inv02 port map ( Y=>nx10236, A=>nx10468);
   ix10237 : inv02 port map ( Y=>nx10238, A=>nx10468);
   ix10239 : inv02 port map ( Y=>nx10240, A=>nx10468);
   ix10241 : inv02 port map ( Y=>nx10242, A=>nx10470);
   ix10243 : inv02 port map ( Y=>nx10244, A=>nx10470);
   ix10245 : inv02 port map ( Y=>nx10246, A=>nx10470);
   ix10247 : inv02 port map ( Y=>nx10248, A=>nx10470);
   ix10249 : inv02 port map ( Y=>nx10250, A=>nx10470);
   ix10251 : inv02 port map ( Y=>nx10252, A=>nx10470);
   ix10253 : inv02 port map ( Y=>nx10254, A=>nx10470);
   ix10255 : inv02 port map ( Y=>nx10256, A=>nx10472);
   ix10257 : inv02 port map ( Y=>nx10258, A=>nx10472);
   ix10259 : inv02 port map ( Y=>nx10260, A=>nx10472);
   ix10261 : inv02 port map ( Y=>nx10262, A=>nx10472);
   ix10263 : inv02 port map ( Y=>nx10264, A=>nx10472);
   ix10265 : inv02 port map ( Y=>nx10266, A=>nx10472);
   ix10267 : inv02 port map ( Y=>nx10268, A=>nx10472);
   ix10269 : inv02 port map ( Y=>nx10270, A=>nx10474);
   ix10271 : inv02 port map ( Y=>nx10272, A=>nx10474);
   ix10273 : inv02 port map ( Y=>nx10274, A=>nx10474);
   ix10275 : inv02 port map ( Y=>nx10276, A=>nx10474);
   ix10277 : inv02 port map ( Y=>nx10278, A=>nx10474);
   ix10279 : inv02 port map ( Y=>nx10280, A=>nx10474);
   ix10281 : inv02 port map ( Y=>nx10282, A=>nx10474);
   ix10283 : inv02 port map ( Y=>nx10284, A=>nx10476);
   ix10285 : inv02 port map ( Y=>nx10286, A=>nx10476);
   ix10287 : inv02 port map ( Y=>nx10288, A=>nx10476);
   ix10289 : inv02 port map ( Y=>nx10290, A=>nx10476);
   ix10291 : inv02 port map ( Y=>nx10292, A=>nx10476);
   ix10293 : inv02 port map ( Y=>nx10294, A=>nx10476);
   ix10295 : inv02 port map ( Y=>nx10296, A=>nx10476);
   ix10297 : inv02 port map ( Y=>nx10298, A=>nx10478);
   ix10299 : inv02 port map ( Y=>nx10300, A=>nx10478);
   ix10301 : inv02 port map ( Y=>nx10302, A=>nx10478);
   ix10303 : inv02 port map ( Y=>nx10304, A=>nx10478);
   ix10305 : inv02 port map ( Y=>nx10306, A=>nx10478);
   ix10307 : buf02 port map ( Y=>nx10308, A=>ACKF);
   ix10309 : buf02 port map ( Y=>nx10310, A=>ACKF);
   ix10311 : buf02 port map ( Y=>nx10312, A=>DataIOut_15);
   ix10313 : buf02 port map ( Y=>nx10314, A=>DataIOut_15);
   ix10315 : buf02 port map ( Y=>nx10316, A=>DataIOut_14);
   ix10317 : buf02 port map ( Y=>nx10318, A=>DataIOut_14);
   ix10319 : buf02 port map ( Y=>nx10320, A=>DataIOut_13);
   ix10321 : buf02 port map ( Y=>nx10322, A=>DataIOut_13);
   ix10323 : buf02 port map ( Y=>nx10324, A=>DataIOut_12);
   ix10325 : buf02 port map ( Y=>nx10326, A=>DataIOut_12);
   ix10327 : buf02 port map ( Y=>nx10328, A=>DataIOut_11);
   ix10329 : buf02 port map ( Y=>nx10330, A=>DataIOut_11);
   ix10331 : buf02 port map ( Y=>nx10332, A=>DataIOut_10);
   ix10333 : buf02 port map ( Y=>nx10334, A=>DataIOut_10);
   ix10335 : buf02 port map ( Y=>nx10336, A=>DataIOut_9);
   ix10337 : buf02 port map ( Y=>nx10338, A=>DataIOut_9);
   ix10339 : buf02 port map ( Y=>nx10340, A=>DataIOut_8);
   ix10341 : buf02 port map ( Y=>nx10342, A=>DataIOut_8);
   ix10343 : buf02 port map ( Y=>nx10344, A=>DataIOut_7);
   ix10345 : buf02 port map ( Y=>nx10346, A=>DataIOut_7);
   ix10347 : buf02 port map ( Y=>nx10348, A=>DataIOut_6);
   ix10349 : buf02 port map ( Y=>nx10350, A=>DataIOut_6);
   ix10351 : buf02 port map ( Y=>nx10352, A=>DataIOut_5);
   ix10353 : buf02 port map ( Y=>nx10354, A=>DataIOut_5);
   ix10355 : buf02 port map ( Y=>nx10356, A=>DataIOut_4);
   ix10357 : buf02 port map ( Y=>nx10358, A=>DataIOut_4);
   ix10359 : buf02 port map ( Y=>nx10360, A=>DataIOut_3);
   ix10361 : buf02 port map ( Y=>nx10362, A=>DataIOut_3);
   ix10363 : buf02 port map ( Y=>nx10364, A=>DataIOut_2);
   ix10365 : buf02 port map ( Y=>nx10366, A=>DataIOut_2);
   ix10367 : buf02 port map ( Y=>nx10368, A=>DataIOut_1);
   ix10369 : buf02 port map ( Y=>nx10370, A=>DataIOut_1);
   ix10371 : buf02 port map ( Y=>nx10372, A=>DataIOut_0);
   ix10373 : buf02 port map ( Y=>nx10374, A=>DataIOut_0);
   ix10375 : buf02 port map ( Y=>nx10376, A=>LayerInfoOut_8);
   ix10377 : buf02 port map ( Y=>nx10378, A=>LayerInfoOut_8);
   ix10379 : buf02 port map ( Y=>nx10380, A=>LayerInfoOut_7);
   ix10381 : buf02 port map ( Y=>nx10382, A=>LayerInfoOut_7);
   ix10383 : buf02 port map ( Y=>nx10384, A=>LayerInfoOut_6);
   ix10385 : buf02 port map ( Y=>nx10386, A=>LayerInfoOut_6);
   ix10387 : buf02 port map ( Y=>nx10388, A=>LayerInfoOut_5);
   ix10389 : buf02 port map ( Y=>nx10390, A=>LayerInfoOut_5);
   ix10391 : buf02 port map ( Y=>nx10392, A=>LayerInfoOut_4);
   ix10393 : buf02 port map ( Y=>nx10394, A=>LayerInfoOut_4);
   ix10395 : buf02 port map ( Y=>nx10396, A=>ConvOuput_15);
   ix10397 : buf02 port map ( Y=>nx10398, A=>NumOfFilters_3);
   ix10399 : buf02 port map ( Y=>nx10400, A=>NumOfFilters_2);
   ix10401 : buf02 port map ( Y=>nx10402, A=>NumOfFilters_1);
   ix10403 : buf02 port map ( Y=>nx10404, A=>NumOfFilters_0);
   ix10405 : buf02 port map ( Y=>nx10406, A=>CNDepthoutput_3);
   ix10407 : buf02 port map ( Y=>nx10408, A=>CNDepthoutput_2);
   ix10409 : buf02 port map ( Y=>nx10410, A=>CNDepthoutput_1);
   ix10411 : buf02 port map ( Y=>nx10412, A=>CNDepthoutput_0);
   ix10413 : inv02 port map ( Y=>nx10414, A=>nx10436);
   ix10415 : inv02 port map ( Y=>nx10416, A=>nx10436);
   ix10417 : inv02 port map ( Y=>nx10418, A=>nx10436);
   ix10419 : inv02 port map ( Y=>nx10420, A=>nx10436);
   ix10421 : inv02 port map ( Y=>nx10422, A=>nx10438);
   ix10423 : inv02 port map ( Y=>nx10424, A=>nx10438);
   ix10425 : inv02 port map ( Y=>nx10426, A=>nx10438);
   ix10427 : inv02 port map ( Y=>nx10428, A=>nx10438);
   ix10429 : inv02 port map ( Y=>nx10430, A=>nx10438);
   ix10431 : inv02 port map ( Y=>nx10432, A=>done_EXMPLR);
   ix10433 : inv02 port map ( Y=>nx10434, A=>done_EXMPLR);
   ix10435 : inv02 port map ( Y=>nx10436, A=>CLK);
   ix10437 : inv02 port map ( Y=>nx10438, A=>CLK);
   ix10439 : inv02 port map ( Y=>nx10440, A=>DataFOut_399);
   ix10441 : inv02 port map ( Y=>nx10442, A=>nx10484);
   ix10443 : inv02 port map ( Y=>nx10444, A=>nx10484);
   ix10445 : inv02 port map ( Y=>nx10446, A=>nx10484);
   ix10447 : inv02 port map ( Y=>nx10448, A=>nx10484);
   ix10449 : inv02 port map ( Y=>nx10450, A=>nx10484);
   ix10451 : inv02 port map ( Y=>nx10452, A=>nx10484);
   ix10453 : inv02 port map ( Y=>nx10454, A=>nx10484);
   ix10455 : inv02 port map ( Y=>nx10456, A=>nx10486);
   ix10457 : inv02 port map ( Y=>nx10458, A=>nx10486);
   ix10459 : inv02 port map ( Y=>nx10460, A=>nx10486);
   ix10461 : inv02 port map ( Y=>nx10462, A=>nx10486);
   ix10463 : inv02 port map ( Y=>nx10464, A=>nx10486);
   ix10465 : inv02 port map ( Y=>nx10466, A=>nx10486);
   ix10467 : inv02 port map ( Y=>nx10468, A=>nx10486);
   ix10469 : inv02 port map ( Y=>nx10470, A=>nx10488);
   ix10471 : inv02 port map ( Y=>nx10472, A=>nx10488);
   ix10473 : inv02 port map ( Y=>nx10474, A=>nx10488);
   ix10475 : inv02 port map ( Y=>nx10476, A=>nx10488);
   ix10477 : inv02 port map ( Y=>nx10478, A=>nx10488);
   ix10483 : inv02 port map ( Y=>nx10484, A=>nx10440);
   ix10485 : inv02 port map ( Y=>nx10486, A=>nx10440);
   ix10487 : inv02 port map ( Y=>nx10488, A=>nx10440);
   ix10489 : inv02 port map ( Y=>nx10490, A=>DataFOut_399);
   ix241 : oai22 port map ( Y=>nx240, A0=>X, A1=>nx10496, B0=>nx9768, B1=>
      nx20);
   ix10495 : inv01 port map ( Y=>nx10496, A=>nx9960);
   ix187 : nand03 port map ( Y=>nx186, A0=>nx9870, A1=>nx10498, A2=>nx180);
   ix10497 : inv01 port map ( Y=>nx10498, A=>nx9958);
   ix301 : nor02ii port map ( Y=>nx300, A0=>nx9792, A1=>next_state_dup_134);
   ix113 : nor02ii port map ( Y=>nx112, A0=>nx9849, A1=>next_state_dup_26);
   ix323 : nor02_2x port map ( Y=>nx322, A0=>nx9866, A1=>nx9849);
   ix9749 : mux21_ni port map ( Y=>nx9748, A0=>next_state_dup_24, A1=>
      nx10478, S0=>nx10308);
   ix457 : nor02_2x port map ( Y=>nx456, A0=>nx9765, A1=>nx9870);
   ix9906 : nor02ii port map ( Y=>nx9905, A0=>nx9966, A1=>nx9858);
   ix519 : nor02ii port map ( Y=>SwitchClk, A0=>nx9792, A1=>nx10028);
   lat_SaveAckLatch_u1 : latchr port map ( QB=>nx5, D=>nx9063, CLK=>nx186, R
      =>zero_11);
   lat_SaveAckLatch_u2 : inv01 port map ( Y=>SaveAckLatch, A=>nx5);
   lat_SaveAckLatch_u3 : buf02 port map ( Y=>nx9941, A=>nx5);
   ix10499 : buf02 port map ( Y=>nx10500, A=>LayerInfoOut_14);
   ix10501 : buf02 port map ( Y=>nx10502, A=>LayerInfoOut_14);
   ix10503 : inv02 port map ( Y=>nx10504, A=>nx10438);
end vlsi ;


