library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity ReadInfoState is
  port (
    CLK,state:in std_logic;
    noOfLayersReg,filterAddressReg
  ) ;
end ReadInfoState;
architecture archReadInfoState of ent is

    signal 

begin

end archReadInfoState ; -- arch