//
// Verilog description for cell Main, 
// Sat May 11 17:20:02 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module Main ( rst, cl, start, dmaStartSignal, done ) ;

    input rst ;
    input cl ;
    input start ;
    inout dmaStartSignal ;
    output done ;

    wire current_state_11, current_state_10, current_state_9, current_state_8, 
         current_state_6, current_state_5, current_state_4, current_state_3, 
         current_state_2, current_state_0, FilterAddressIN_12, 
         FilterAddressIN_11, FilterAddressIN_10, FilterAddressIN_9, 
         FilterAddressIN_8, FilterAddressIN_7, FilterAddressIN_6, 
         FilterAddressIN_5, FilterAddressIN_4, FilterAddressIN_3, 
         FilterAddressIN_2, FilterAddressIN_1, FilterAddressIN_0, 
         FilterAddressOut_12, FilterAddressOut_11, FilterAddressOut_10, 
         FilterAddressOut_9, FilterAddressOut_8, FilterAddressOut_7, 
         FilterAddressOut_6, FilterAddressOut_5, FilterAddressOut_4, 
         FilterAddressOut_3, FilterAddressOut_2, FilterAddressOut_1, 
         FilterAddressOut_0, AddressChangerIN_12, AddressChangerIN_11, 
         AddressChangerIN_10, AddressChangerIN_9, AddressChangerIN_8, 
         AddressChangerIN_7, AddressChangerIN_6, AddressChangerIN_5, 
         AddressChangerIN_4, AddressChangerIN_3, AddressChangerIN_2, 
         AddressChangerIN_1, AddressChangerIN_0, AddressChangerOut_12, 
         AddressChangerOut_11, AddressChangerOut_10, AddressChangerOut_9, 
         AddressChangerOut_8, AddressChangerOut_7, AddressChangerOut_6, 
         AddressChangerOut_5, AddressChangerOut_4, AddressChangerOut_3, 
         AddressChangerOut_2, AddressChangerOut_1, AddressChangerOut_0, 
         ImgAddRegIN_12, ImgAddRegIN_11, ImgAddRegIN_10, ImgAddRegIN_9, 
         ImgAddRegIN_8, ImgAddRegIN_7, ImgAddRegIN_6, ImgAddRegIN_5, 
         ImgAddRegIN_4, ImgAddRegIN_3, ImgAddRegIN_2, ImgAddRegIN_1, 
         ImgAddRegIN_0, ImgAddRegOut_12, ImgAddRegOut_11, ImgAddRegOut_10, 
         ImgAddRegOut_9, ImgAddRegOut_8, ImgAddRegOut_7, ImgAddRegOut_6, 
         ImgAddRegOut_5, ImgAddRegOut_4, ImgAddRegOut_3, ImgAddRegOut_2, 
         ImgAddRegOut_1, ImgAddRegOut_0, TriStateCounterOUT_12, 
         TriStateCounterOUT_11, TriStateCounterOUT_10, TriStateCounterOUT_9, 
         TriStateCounterOUT_8, TriStateCounterOUT_7, TriStateCounterOUT_6, 
         TriStateCounterOUT_5, TriStateCounterOUT_4, TriStateCounterOUT_3, 
         TriStateCounterOUT_2, TriStateCounterOUT_1, TriStateCounterOUT_0, 
         ImgAddACKTriIN_0, ReadF, AddressF_12, AddressF_11, AddressF_10, 
         AddressF_9, AddressF_8, AddressF_7, AddressF_6, AddressF_5, AddressF_4, 
         AddressF_3, AddressF_2, AddressF_1, AddressF_0, DataFOut_399, ACKF, 
         WriteI, ReadI, AddressI_12, AddressI_11, AddressI_10, AddressI_9, 
         AddressI_8, AddressI_7, AddressI_6, AddressI_5, AddressI_4, AddressI_3, 
         AddressI_2, AddressI_1, AddressI_0, DataIIn_15, DataIIn_14, DataIIn_13, 
         DataIIn_12, DataIIn_11, DataIIn_10, DataIIn_9, DataIIn_8, DataIIn_7, 
         DataIIn_6, DataIIn_5, DataIIn_4, DataIIn_3, DataIIn_2, DataIIn_1, 
         DataIIn_0, DataIOut_447, DataIOut_446, DataIOut_445, DataIOut_444, 
         DataIOut_443, DataIOut_442, DataIOut_441, DataIOut_440, DataIOut_439, 
         DataIOut_438, DataIOut_437, DataIOut_436, DataIOut_435, DataIOut_434, 
         DataIOut_433, DataIOut_432, DataIOut_431, DataIOut_430, DataIOut_429, 
         DataIOut_428, DataIOut_427, DataIOut_426, DataIOut_425, DataIOut_424, 
         DataIOut_423, DataIOut_422, DataIOut_421, DataIOut_420, DataIOut_419, 
         DataIOut_418, DataIOut_417, DataIOut_416, DataIOut_415, DataIOut_414, 
         DataIOut_413, DataIOut_412, DataIOut_411, DataIOut_410, DataIOut_409, 
         DataIOut_408, DataIOut_407, DataIOut_406, DataIOut_405, DataIOut_404, 
         DataIOut_403, DataIOut_402, DataIOut_401, DataIOut_400, DataIOut_399, 
         DataIOut_398, DataIOut_397, DataIOut_396, DataIOut_395, DataIOut_394, 
         DataIOut_393, DataIOut_392, DataIOut_391, DataIOut_390, DataIOut_389, 
         DataIOut_388, DataIOut_387, DataIOut_386, DataIOut_385, DataIOut_384, 
         DataIOut_383, DataIOut_382, DataIOut_381, DataIOut_380, DataIOut_379, 
         DataIOut_378, DataIOut_377, DataIOut_376, DataIOut_375, DataIOut_374, 
         DataIOut_373, DataIOut_372, DataIOut_371, DataIOut_370, DataIOut_369, 
         DataIOut_368, DataIOut_367, DataIOut_366, DataIOut_365, DataIOut_364, 
         DataIOut_363, DataIOut_362, DataIOut_361, DataIOut_360, DataIOut_359, 
         DataIOut_358, DataIOut_357, DataIOut_356, DataIOut_355, DataIOut_354, 
         DataIOut_353, DataIOut_352, DataIOut_351, DataIOut_350, DataIOut_349, 
         DataIOut_348, DataIOut_347, DataIOut_346, DataIOut_345, DataIOut_344, 
         DataIOut_343, DataIOut_342, DataIOut_341, DataIOut_340, DataIOut_339, 
         DataIOut_338, DataIOut_337, DataIOut_336, DataIOut_335, DataIOut_334, 
         DataIOut_333, DataIOut_332, DataIOut_331, DataIOut_330, DataIOut_329, 
         DataIOut_328, DataIOut_327, DataIOut_326, DataIOut_325, DataIOut_324, 
         DataIOut_323, DataIOut_322, DataIOut_321, DataIOut_320, DataIOut_319, 
         DataIOut_318, DataIOut_317, DataIOut_316, DataIOut_315, DataIOut_314, 
         DataIOut_313, DataIOut_312, DataIOut_311, DataIOut_310, DataIOut_309, 
         DataIOut_308, DataIOut_307, DataIOut_306, DataIOut_305, DataIOut_304, 
         DataIOut_303, DataIOut_302, DataIOut_301, DataIOut_300, DataIOut_299, 
         DataIOut_298, DataIOut_297, DataIOut_296, DataIOut_295, DataIOut_294, 
         DataIOut_293, DataIOut_292, DataIOut_291, DataIOut_290, DataIOut_289, 
         DataIOut_288, DataIOut_287, DataIOut_286, DataIOut_285, DataIOut_284, 
         DataIOut_283, DataIOut_282, DataIOut_281, DataIOut_280, DataIOut_279, 
         DataIOut_278, DataIOut_277, DataIOut_276, DataIOut_275, DataIOut_274, 
         DataIOut_273, DataIOut_272, DataIOut_271, DataIOut_270, DataIOut_269, 
         DataIOut_268, DataIOut_267, DataIOut_266, DataIOut_265, DataIOut_264, 
         DataIOut_263, DataIOut_262, DataIOut_261, DataIOut_260, DataIOut_259, 
         DataIOut_258, DataIOut_257, DataIOut_256, DataIOut_255, DataIOut_254, 
         DataIOut_253, DataIOut_252, DataIOut_251, DataIOut_250, DataIOut_249, 
         DataIOut_248, DataIOut_247, DataIOut_246, DataIOut_245, DataIOut_244, 
         DataIOut_243, DataIOut_242, DataIOut_241, DataIOut_240, DataIOut_239, 
         DataIOut_238, DataIOut_237, DataIOut_236, DataIOut_235, DataIOut_234, 
         DataIOut_233, DataIOut_232, DataIOut_231, DataIOut_230, DataIOut_229, 
         DataIOut_228, DataIOut_227, DataIOut_226, DataIOut_225, DataIOut_224, 
         DataIOut_223, DataIOut_222, DataIOut_221, DataIOut_220, DataIOut_219, 
         DataIOut_218, DataIOut_217, DataIOut_216, DataIOut_215, DataIOut_214, 
         DataIOut_213, DataIOut_212, DataIOut_211, DataIOut_210, DataIOut_209, 
         DataIOut_208, DataIOut_207, DataIOut_206, DataIOut_205, DataIOut_204, 
         DataIOut_203, DataIOut_202, DataIOut_201, DataIOut_200, DataIOut_199, 
         DataIOut_198, DataIOut_197, DataIOut_196, DataIOut_195, DataIOut_194, 
         DataIOut_193, DataIOut_192, DataIOut_191, DataIOut_190, DataIOut_189, 
         DataIOut_188, DataIOut_187, DataIOut_186, DataIOut_185, DataIOut_184, 
         DataIOut_183, DataIOut_182, DataIOut_181, DataIOut_180, DataIOut_179, 
         DataIOut_178, DataIOut_177, DataIOut_176, DataIOut_175, DataIOut_174, 
         DataIOut_173, DataIOut_172, DataIOut_171, DataIOut_170, DataIOut_169, 
         DataIOut_168, DataIOut_167, DataIOut_166, DataIOut_165, DataIOut_164, 
         DataIOut_163, DataIOut_162, DataIOut_161, DataIOut_160, DataIOut_159, 
         DataIOut_158, DataIOut_157, DataIOut_156, DataIOut_155, DataIOut_154, 
         DataIOut_153, DataIOut_152, DataIOut_151, DataIOut_150, DataIOut_149, 
         DataIOut_148, DataIOut_147, DataIOut_146, DataIOut_145, DataIOut_144, 
         DataIOut_143, DataIOut_142, DataIOut_141, DataIOut_140, DataIOut_139, 
         DataIOut_138, DataIOut_137, DataIOut_136, DataIOut_135, DataIOut_134, 
         DataIOut_133, DataIOut_132, DataIOut_131, DataIOut_130, DataIOut_129, 
         DataIOut_128, DataIOut_127, DataIOut_126, DataIOut_125, DataIOut_124, 
         DataIOut_123, DataIOut_122, DataIOut_121, DataIOut_120, DataIOut_119, 
         DataIOut_118, DataIOut_117, DataIOut_116, DataIOut_115, DataIOut_114, 
         DataIOut_113, DataIOut_112, DataIOut_111, DataIOut_110, DataIOut_109, 
         DataIOut_108, DataIOut_107, DataIOut_106, DataIOut_105, DataIOut_104, 
         DataIOut_103, DataIOut_102, DataIOut_101, DataIOut_100, DataIOut_99, 
         DataIOut_98, DataIOut_97, DataIOut_96, DataIOut_95, DataIOut_94, 
         DataIOut_93, DataIOut_92, DataIOut_91, DataIOut_90, DataIOut_89, 
         DataIOut_88, DataIOut_87, DataIOut_86, DataIOut_85, DataIOut_84, 
         DataIOut_83, DataIOut_82, DataIOut_81, DataIOut_80, DataIOut_79, 
         DataIOut_78, DataIOut_77, DataIOut_76, DataIOut_75, DataIOut_74, 
         DataIOut_73, DataIOut_72, DataIOut_71, DataIOut_70, DataIOut_69, 
         DataIOut_68, DataIOut_67, DataIOut_66, DataIOut_65, DataIOut_64, 
         DataIOut_63, DataIOut_62, DataIOut_61, DataIOut_60, DataIOut_59, 
         DataIOut_58, DataIOut_57, DataIOut_56, DataIOut_55, DataIOut_54, 
         DataIOut_53, DataIOut_52, DataIOut_51, DataIOut_50, DataIOut_49, 
         DataIOut_48, DataIOut_47, DataIOut_46, DataIOut_45, DataIOut_44, 
         DataIOut_43, DataIOut_42, DataIOut_41, DataIOut_40, DataIOut_39, 
         DataIOut_38, DataIOut_37, DataIOut_36, DataIOut_35, DataIOut_34, 
         DataIOut_33, DataIOut_32, DataIOut_31, DataIOut_30, DataIOut_29, 
         DataIOut_28, DataIOut_27, DataIOut_26, DataIOut_25, DataIOut_24, 
         DataIOut_23, DataIOut_22, DataIOut_21, DataIOut_20, DataIOut_19, 
         DataIOut_18, DataIOut_17, DataIOut_16, DataIOut_15, DataIOut_14, 
         DataIOut_13, DataIOut_12, DataIOut_11, DataIOut_10, DataIOut_9, 
         DataIOut_8, DataIOut_7, DataIOut_6, DataIOut_5, DataIOut_4, DataIOut_3, 
         DataIOut_2, DataIOut_1, DataIOut_0, NoOfLayers_1, NoOfLayers_0, 
         LayerInfoOut_15, LayerInfoOut_14, LayerInfoOut_12, LayerInfoOut_11, 
         LayerInfoOut_10, LayerInfoOut_9, LayerInfoOut_8, LayerInfoOut_7, 
         LayerInfoOut_6, LayerInfoOut_5, LayerInfoOut_4, LayerInfoOut_3, 
         LayerInfoOut_2, LayerInfoOut_1, LayerInfoOut_0, ImgWidthOut_15, 
         ImgWidthOut_14, ImgWidthOut_13, ImgWidthOut_12, ImgWidthOut_11, 
         ImgWidthOut_10, ImgWidthOut_9, ImgWidthOut_8, ImgWidthOut_7, 
         ImgWidthOut_6, ImgWidthOut_5, ImgWidthOut_4, ImgWidthOut_3, 
         ImgWidthOut_2, ImgWidthOut_1, ImgWidthOut_0, WidthSquareOut_9, 
         WidthSquareOut_8, WidthSquareOut_7, WidthSquareOut_6, WidthSquareOut_5, 
         WidthSquareOut_4, WidthSquareOut_3, WidthSquareOut_2, WidthSquareOut_1, 
         WidthSquareOut_0, Bias0_15, Bias0_14, Bias0_13, Bias0_12, Bias0_11, 
         Bias0_10, Bias0_9, Bias0_8, Bias0_7, Bias0_6, Bias0_5, Bias0_4, Bias0_3, 
         Bias0_2, Bias0_1, Bias0_0, Bias1_15, Bias1_14, Bias1_13, Bias1_12, 
         Bias1_11, Bias1_10, Bias1_9, Bias1_8, Bias1_7, Bias1_6, Bias1_5, 
         Bias1_4, Bias1_3, Bias1_2, Bias1_1, Bias1_0, Bias2_15, Bias2_14, 
         Bias2_13, Bias2_12, Bias2_11, Bias2_10, Bias2_9, Bias2_8, Bias2_7, 
         Bias2_6, Bias2_5, Bias2_4, Bias2_3, Bias2_2, Bias2_1, Bias2_0, Bias3_15, 
         Bias3_14, Bias3_13, Bias3_12, Bias3_11, Bias3_10, Bias3_9, Bias3_8, 
         Bias3_7, Bias3_6, Bias3_5, Bias3_4, Bias3_3, Bias3_2, Bias3_1, Bias3_0, 
         Bias4_15, Bias4_14, Bias4_13, Bias4_12, Bias4_11, Bias4_10, Bias4_9, 
         Bias4_8, Bias4_7, Bias4_6, Bias4_5, Bias4_4, Bias4_3, Bias4_2, Bias4_1, 
         Bias4_0, Bias5_15, Bias5_14, Bias5_13, Bias5_12, Bias5_11, Bias5_10, 
         Bias5_9, Bias5_8, Bias5_7, Bias5_6, Bias5_5, Bias5_4, Bias5_3, Bias5_2, 
         Bias5_1, Bias5_0, Bias6_15, Bias6_14, Bias6_13, Bias6_12, Bias6_11, 
         Bias6_10, Bias6_9, Bias6_8, Bias6_7, Bias6_6, Bias6_5, Bias6_4, Bias6_3, 
         Bias6_2, Bias6_1, Bias6_0, Bias7_15, Bias7_14, Bias7_13, Bias7_12, 
         Bias7_11, Bias7_10, Bias7_9, Bias7_8, Bias7_7, Bias7_6, Bias7_5, 
         Bias7_4, Bias7_3, Bias7_2, Bias7_1, Bias7_0, IndicatorF_0, Filter2_399, 
         Filter2_398, Filter2_397, Filter2_396, Filter2_395, Filter2_394, 
         Filter2_393, Filter2_392, Filter2_391, Filter2_390, Filter2_389, 
         Filter2_388, Filter2_387, Filter2_386, Filter2_385, Filter2_384, 
         Filter2_383, Filter2_382, Filter2_381, Filter2_380, Filter2_379, 
         Filter2_378, Filter2_377, Filter2_376, Filter2_375, Filter2_374, 
         Filter2_373, Filter2_372, Filter2_371, Filter2_370, Filter2_369, 
         Filter2_368, Filter2_367, Filter2_366, Filter2_365, Filter2_364, 
         Filter2_363, Filter2_362, Filter2_361, Filter2_360, Filter2_359, 
         Filter2_358, Filter2_357, Filter2_356, Filter2_355, Filter2_354, 
         Filter2_353, Filter2_352, Filter2_351, Filter2_350, Filter2_349, 
         Filter2_348, Filter2_347, Filter2_346, Filter2_345, Filter2_344, 
         Filter2_343, Filter2_342, Filter2_341, Filter2_340, Filter2_339, 
         Filter2_338, Filter2_337, Filter2_336, Filter2_335, Filter2_334, 
         Filter2_333, Filter2_332, Filter2_331, Filter2_330, Filter2_329, 
         Filter2_328, Filter2_327, Filter2_326, Filter2_325, Filter2_324, 
         Filter2_323, Filter2_322, Filter2_321, Filter2_320, Filter2_319, 
         Filter2_318, Filter2_317, Filter2_316, Filter2_315, Filter2_314, 
         Filter2_313, Filter2_312, Filter2_311, Filter2_310, Filter2_309, 
         Filter2_308, Filter2_307, Filter2_306, Filter2_305, Filter2_304, 
         Filter2_303, Filter2_302, Filter2_301, Filter2_300, Filter2_299, 
         Filter2_298, Filter2_297, Filter2_296, Filter2_295, Filter2_294, 
         Filter2_293, Filter2_292, Filter2_291, Filter2_290, Filter2_289, 
         Filter2_288, Filter2_287, Filter2_286, Filter2_285, Filter2_284, 
         Filter2_283, Filter2_282, Filter2_281, Filter2_280, Filter2_279, 
         Filter2_278, Filter2_277, Filter2_276, Filter2_275, Filter2_274, 
         Filter2_273, Filter2_272, Filter2_271, Filter2_270, Filter2_269, 
         Filter2_268, Filter2_267, Filter2_266, Filter2_265, Filter2_264, 
         Filter2_263, Filter2_262, Filter2_261, Filter2_260, Filter2_259, 
         Filter2_258, Filter2_257, Filter2_256, Filter2_255, Filter2_254, 
         Filter2_253, Filter2_252, Filter2_251, Filter2_250, Filter2_249, 
         Filter2_248, Filter2_247, Filter2_246, Filter2_245, Filter2_244, 
         Filter2_243, Filter2_242, Filter2_241, Filter2_240, Filter2_239, 
         Filter2_238, Filter2_237, Filter2_236, Filter2_235, Filter2_234, 
         Filter2_233, Filter2_232, Filter2_231, Filter2_230, Filter2_229, 
         Filter2_228, Filter2_227, Filter2_226, Filter2_225, Filter2_224, 
         Filter2_223, Filter2_222, Filter2_221, Filter2_220, Filter2_219, 
         Filter2_218, Filter2_217, Filter2_216, Filter2_215, Filter2_214, 
         Filter2_213, Filter2_212, Filter2_211, Filter2_210, Filter2_209, 
         Filter2_208, Filter2_207, Filter2_206, Filter2_205, Filter2_204, 
         Filter2_203, Filter2_202, Filter2_201, Filter2_200, Filter2_199, 
         Filter2_198, Filter2_197, Filter2_196, Filter2_195, Filter2_194, 
         Filter2_193, Filter2_192, Filter2_191, Filter2_190, Filter2_189, 
         Filter2_188, Filter2_187, Filter2_186, Filter2_185, Filter2_184, 
         Filter2_183, Filter2_182, Filter2_181, Filter2_180, Filter2_179, 
         Filter2_178, Filter2_177, Filter2_176, Filter2_175, Filter2_174, 
         Filter2_173, Filter2_172, Filter2_171, Filter2_170, Filter2_169, 
         Filter2_168, Filter2_167, Filter2_166, Filter2_165, Filter2_164, 
         Filter2_163, Filter2_162, Filter2_161, Filter2_160, Filter2_159, 
         Filter2_158, Filter2_157, Filter2_156, Filter2_155, Filter2_154, 
         Filter2_153, Filter2_152, Filter2_151, Filter2_150, Filter2_149, 
         Filter2_148, Filter2_147, Filter2_146, Filter2_145, Filter2_144, 
         Filter2_143, Filter2_142, Filter2_141, Filter2_140, Filter2_139, 
         Filter2_138, Filter2_137, Filter2_136, Filter2_135, Filter2_134, 
         Filter2_133, Filter2_132, Filter2_131, Filter2_130, Filter2_129, 
         Filter2_128, Filter2_127, Filter2_126, Filter2_125, Filter2_124, 
         Filter2_123, Filter2_122, Filter2_121, Filter2_120, Filter2_119, 
         Filter2_118, Filter2_117, Filter2_116, Filter2_115, Filter2_114, 
         Filter2_113, Filter2_112, Filter2_111, Filter2_110, Filter2_109, 
         Filter2_108, Filter2_107, Filter2_106, Filter2_105, Filter2_104, 
         Filter2_103, Filter2_102, Filter2_101, Filter2_100, Filter2_99, 
         Filter2_98, Filter2_97, Filter2_96, Filter2_95, Filter2_94, Filter2_93, 
         Filter2_92, Filter2_91, Filter2_90, Filter2_89, Filter2_88, Filter2_87, 
         Filter2_86, Filter2_85, Filter2_84, Filter2_83, Filter2_82, Filter2_81, 
         Filter2_80, Filter2_79, Filter2_78, Filter2_77, Filter2_76, Filter2_75, 
         Filter2_74, Filter2_73, Filter2_72, Filter2_71, Filter2_70, Filter2_69, 
         Filter2_68, Filter2_67, Filter2_66, Filter2_65, Filter2_64, Filter2_63, 
         Filter2_62, Filter2_61, Filter2_60, Filter2_59, Filter2_58, Filter2_57, 
         Filter2_56, Filter2_55, Filter2_54, Filter2_53, Filter2_52, Filter2_51, 
         Filter2_50, Filter2_49, Filter2_48, Filter2_47, Filter2_46, Filter2_45, 
         Filter2_44, Filter2_43, Filter2_42, Filter2_41, Filter2_40, Filter2_39, 
         Filter2_38, Filter2_37, Filter2_36, Filter2_35, Filter2_34, Filter2_33, 
         Filter2_32, Filter2_31, Filter2_30, Filter2_29, Filter2_28, Filter2_27, 
         Filter2_26, Filter2_25, Filter2_24, Filter2_23, Filter2_22, Filter2_21, 
         Filter2_20, Filter2_19, Filter2_18, Filter2_17, Filter2_16, Filter2_15, 
         Filter2_14, Filter2_13, Filter2_12, Filter2_11, Filter2_10, Filter2_9, 
         Filter2_8, Filter2_7, Filter2_6, Filter2_5, Filter2_4, Filter2_3, 
         Filter2_2, Filter2_1, Filter2_0, Filter1_399, Filter1_398, Filter1_397, 
         Filter1_396, Filter1_395, Filter1_394, Filter1_393, Filter1_392, 
         Filter1_391, Filter1_390, Filter1_389, Filter1_388, Filter1_387, 
         Filter1_386, Filter1_385, Filter1_384, Filter1_383, Filter1_382, 
         Filter1_381, Filter1_380, Filter1_379, Filter1_378, Filter1_377, 
         Filter1_376, Filter1_375, Filter1_374, Filter1_373, Filter1_372, 
         Filter1_371, Filter1_370, Filter1_369, Filter1_368, Filter1_367, 
         Filter1_366, Filter1_365, Filter1_364, Filter1_363, Filter1_362, 
         Filter1_361, Filter1_360, Filter1_359, Filter1_358, Filter1_357, 
         Filter1_356, Filter1_355, Filter1_354, Filter1_353, Filter1_352, 
         Filter1_351, Filter1_350, Filter1_349, Filter1_348, Filter1_347, 
         Filter1_346, Filter1_345, Filter1_344, Filter1_343, Filter1_342, 
         Filter1_341, Filter1_340, Filter1_339, Filter1_338, Filter1_337, 
         Filter1_336, Filter1_335, Filter1_334, Filter1_333, Filter1_332, 
         Filter1_331, Filter1_330, Filter1_329, Filter1_328, Filter1_327, 
         Filter1_326, Filter1_325, Filter1_324, Filter1_323, Filter1_322, 
         Filter1_321, Filter1_320, Filter1_319, Filter1_318, Filter1_317, 
         Filter1_316, Filter1_315, Filter1_314, Filter1_313, Filter1_312, 
         Filter1_311, Filter1_310, Filter1_309, Filter1_308, Filter1_307, 
         Filter1_306, Filter1_305, Filter1_304, Filter1_303, Filter1_302, 
         Filter1_301, Filter1_300, Filter1_299, Filter1_298, Filter1_297, 
         Filter1_296, Filter1_295, Filter1_294, Filter1_293, Filter1_292, 
         Filter1_291, Filter1_290, Filter1_289, Filter1_288, Filter1_287, 
         Filter1_286, Filter1_285, Filter1_284, Filter1_283, Filter1_282, 
         Filter1_281, Filter1_280, Filter1_279, Filter1_278, Filter1_277, 
         Filter1_276, Filter1_275, Filter1_274, Filter1_273, Filter1_272, 
         Filter1_271, Filter1_270, Filter1_269, Filter1_268, Filter1_267, 
         Filter1_266, Filter1_265, Filter1_264, Filter1_263, Filter1_262, 
         Filter1_261, Filter1_260, Filter1_259, Filter1_258, Filter1_257, 
         Filter1_256, Filter1_255, Filter1_254, Filter1_253, Filter1_252, 
         Filter1_251, Filter1_250, Filter1_249, Filter1_248, Filter1_247, 
         Filter1_246, Filter1_245, Filter1_244, Filter1_243, Filter1_242, 
         Filter1_241, Filter1_240, Filter1_239, Filter1_238, Filter1_237, 
         Filter1_236, Filter1_235, Filter1_234, Filter1_233, Filter1_232, 
         Filter1_231, Filter1_230, Filter1_229, Filter1_228, Filter1_227, 
         Filter1_226, Filter1_225, Filter1_224, Filter1_223, Filter1_222, 
         Filter1_221, Filter1_220, Filter1_219, Filter1_218, Filter1_217, 
         Filter1_216, Filter1_215, Filter1_214, Filter1_213, Filter1_212, 
         Filter1_211, Filter1_210, Filter1_209, Filter1_208, Filter1_207, 
         Filter1_206, Filter1_205, Filter1_204, Filter1_203, Filter1_202, 
         Filter1_201, Filter1_200, Filter1_199, Filter1_198, Filter1_197, 
         Filter1_196, Filter1_195, Filter1_194, Filter1_193, Filter1_192, 
         Filter1_191, Filter1_190, Filter1_189, Filter1_188, Filter1_187, 
         Filter1_186, Filter1_185, Filter1_184, Filter1_183, Filter1_182, 
         Filter1_181, Filter1_180, Filter1_179, Filter1_178, Filter1_177, 
         Filter1_176, Filter1_175, Filter1_174, Filter1_173, Filter1_172, 
         Filter1_171, Filter1_170, Filter1_169, Filter1_168, Filter1_167, 
         Filter1_166, Filter1_165, Filter1_164, Filter1_163, Filter1_162, 
         Filter1_161, Filter1_160, Filter1_159, Filter1_158, Filter1_157, 
         Filter1_156, Filter1_155, Filter1_154, Filter1_153, Filter1_152, 
         Filter1_151, Filter1_150, Filter1_149, Filter1_148, Filter1_147, 
         Filter1_146, Filter1_145, Filter1_144, Filter1_143, Filter1_142, 
         Filter1_141, Filter1_140, Filter1_139, Filter1_138, Filter1_137, 
         Filter1_136, Filter1_135, Filter1_134, Filter1_133, Filter1_132, 
         Filter1_131, Filter1_130, Filter1_129, Filter1_128, Filter1_127, 
         Filter1_126, Filter1_125, Filter1_124, Filter1_123, Filter1_122, 
         Filter1_121, Filter1_120, Filter1_119, Filter1_118, Filter1_117, 
         Filter1_116, Filter1_115, Filter1_114, Filter1_113, Filter1_112, 
         Filter1_111, Filter1_110, Filter1_109, Filter1_108, Filter1_107, 
         Filter1_106, Filter1_105, Filter1_104, Filter1_103, Filter1_102, 
         Filter1_101, Filter1_100, Filter1_99, Filter1_98, Filter1_97, 
         Filter1_96, Filter1_95, Filter1_94, Filter1_93, Filter1_92, Filter1_91, 
         Filter1_90, Filter1_89, Filter1_88, Filter1_87, Filter1_86, Filter1_85, 
         Filter1_84, Filter1_83, Filter1_82, Filter1_81, Filter1_80, Filter1_79, 
         Filter1_78, Filter1_77, Filter1_76, Filter1_75, Filter1_74, Filter1_73, 
         Filter1_72, Filter1_71, Filter1_70, Filter1_69, Filter1_68, Filter1_67, 
         Filter1_66, Filter1_65, Filter1_64, Filter1_63, Filter1_62, Filter1_61, 
         Filter1_60, Filter1_59, Filter1_58, Filter1_57, Filter1_56, Filter1_55, 
         Filter1_54, Filter1_53, Filter1_52, Filter1_51, Filter1_50, Filter1_49, 
         Filter1_48, Filter1_47, Filter1_46, Filter1_45, Filter1_44, Filter1_43, 
         Filter1_42, Filter1_41, Filter1_40, Filter1_39, Filter1_38, Filter1_37, 
         Filter1_36, Filter1_35, Filter1_34, Filter1_33, Filter1_32, Filter1_31, 
         Filter1_30, Filter1_29, Filter1_28, Filter1_27, Filter1_26, Filter1_25, 
         Filter1_24, Filter1_23, Filter1_22, Filter1_21, Filter1_20, Filter1_19, 
         Filter1_18, Filter1_17, Filter1_16, Filter1_15, Filter1_14, Filter1_13, 
         Filter1_12, Filter1_11, Filter1_10, Filter1_9, Filter1_8, Filter1_7, 
         Filter1_6, Filter1_5, Filter1_4, Filter1_3, Filter1_2, Filter1_1, 
         Filter1_0, IndicatorI_0, ImgCounterOuput_2, ImgCounterOuput_1, 
         ImgCounterOuput_0, OutputImg0_79, OutputImg0_78, OutputImg0_77, 
         OutputImg0_76, OutputImg0_75, OutputImg0_74, OutputImg0_73, 
         OutputImg0_72, OutputImg0_71, OutputImg0_70, OutputImg0_69, 
         OutputImg0_68, OutputImg0_67, OutputImg0_66, OutputImg0_65, 
         OutputImg0_64, OutputImg0_63, OutputImg0_62, OutputImg0_61, 
         OutputImg0_60, OutputImg0_59, OutputImg0_58, OutputImg0_57, 
         OutputImg0_56, OutputImg0_55, OutputImg0_54, OutputImg0_53, 
         OutputImg0_52, OutputImg0_51, OutputImg0_50, OutputImg0_49, 
         OutputImg0_48, OutputImg0_47, OutputImg0_46, OutputImg0_45, 
         OutputImg0_44, OutputImg0_43, OutputImg0_42, OutputImg0_41, 
         OutputImg0_40, OutputImg0_39, OutputImg0_38, OutputImg0_37, 
         OutputImg0_36, OutputImg0_35, OutputImg0_34, OutputImg0_33, 
         OutputImg0_32, OutputImg0_31, OutputImg0_30, OutputImg0_29, 
         OutputImg0_28, OutputImg0_27, OutputImg0_26, OutputImg0_25, 
         OutputImg0_24, OutputImg0_23, OutputImg0_22, OutputImg0_21, 
         OutputImg0_20, OutputImg0_19, OutputImg0_18, OutputImg0_17, 
         OutputImg0_16, OutputImg0_15, OutputImg0_14, OutputImg0_13, 
         OutputImg0_12, OutputImg0_11, OutputImg0_10, OutputImg0_9, OutputImg0_8, 
         OutputImg0_7, OutputImg0_6, OutputImg0_5, OutputImg0_4, OutputImg0_3, 
         OutputImg0_2, OutputImg0_1, OutputImg0_0, OutputImg1_79, OutputImg1_78, 
         OutputImg1_77, OutputImg1_76, OutputImg1_75, OutputImg1_74, 
         OutputImg1_73, OutputImg1_72, OutputImg1_71, OutputImg1_70, 
         OutputImg1_69, OutputImg1_68, OutputImg1_67, OutputImg1_66, 
         OutputImg1_65, OutputImg1_64, OutputImg1_63, OutputImg1_62, 
         OutputImg1_61, OutputImg1_60, OutputImg1_59, OutputImg1_58, 
         OutputImg1_57, OutputImg1_56, OutputImg1_55, OutputImg1_54, 
         OutputImg1_53, OutputImg1_52, OutputImg1_51, OutputImg1_50, 
         OutputImg1_49, OutputImg1_48, OutputImg1_47, OutputImg1_46, 
         OutputImg1_45, OutputImg1_44, OutputImg1_43, OutputImg1_42, 
         OutputImg1_41, OutputImg1_40, OutputImg1_39, OutputImg1_38, 
         OutputImg1_37, OutputImg1_36, OutputImg1_35, OutputImg1_34, 
         OutputImg1_33, OutputImg1_32, OutputImg1_31, OutputImg1_30, 
         OutputImg1_29, OutputImg1_28, OutputImg1_27, OutputImg1_26, 
         OutputImg1_25, OutputImg1_24, OutputImg1_23, OutputImg1_22, 
         OutputImg1_21, OutputImg1_20, OutputImg1_19, OutputImg1_18, 
         OutputImg1_17, OutputImg1_16, OutputImg1_15, OutputImg1_14, 
         OutputImg1_13, OutputImg1_12, OutputImg1_11, OutputImg1_10, 
         OutputImg1_9, OutputImg1_8, OutputImg1_7, OutputImg1_6, OutputImg1_5, 
         OutputImg1_4, OutputImg1_3, OutputImg1_2, OutputImg1_1, OutputImg1_0, 
         OutputImg2_79, OutputImg2_78, OutputImg2_77, OutputImg2_76, 
         OutputImg2_75, OutputImg2_74, OutputImg2_73, OutputImg2_72, 
         OutputImg2_71, OutputImg2_70, OutputImg2_69, OutputImg2_68, 
         OutputImg2_67, OutputImg2_66, OutputImg2_65, OutputImg2_64, 
         OutputImg2_63, OutputImg2_62, OutputImg2_61, OutputImg2_60, 
         OutputImg2_59, OutputImg2_58, OutputImg2_57, OutputImg2_56, 
         OutputImg2_55, OutputImg2_54, OutputImg2_53, OutputImg2_52, 
         OutputImg2_51, OutputImg2_50, OutputImg2_49, OutputImg2_48, 
         OutputImg2_47, OutputImg2_46, OutputImg2_45, OutputImg2_44, 
         OutputImg2_43, OutputImg2_42, OutputImg2_41, OutputImg2_40, 
         OutputImg2_39, OutputImg2_38, OutputImg2_37, OutputImg2_36, 
         OutputImg2_35, OutputImg2_34, OutputImg2_33, OutputImg2_32, 
         OutputImg2_31, OutputImg2_30, OutputImg2_29, OutputImg2_28, 
         OutputImg2_27, OutputImg2_26, OutputImg2_25, OutputImg2_24, 
         OutputImg2_23, OutputImg2_22, OutputImg2_21, OutputImg2_20, 
         OutputImg2_19, OutputImg2_18, OutputImg2_17, OutputImg2_16, 
         OutputImg2_15, OutputImg2_14, OutputImg2_13, OutputImg2_12, 
         OutputImg2_11, OutputImg2_10, OutputImg2_9, OutputImg2_8, OutputImg2_7, 
         OutputImg2_6, OutputImg2_5, OutputImg2_4, OutputImg2_3, OutputImg2_2, 
         OutputImg2_1, OutputImg2_0, OutputImg3_79, OutputImg3_78, OutputImg3_77, 
         OutputImg3_76, OutputImg3_75, OutputImg3_74, OutputImg3_73, 
         OutputImg3_72, OutputImg3_71, OutputImg3_70, OutputImg3_69, 
         OutputImg3_68, OutputImg3_67, OutputImg3_66, OutputImg3_65, 
         OutputImg3_64, OutputImg3_63, OutputImg3_62, OutputImg3_61, 
         OutputImg3_60, OutputImg3_59, OutputImg3_58, OutputImg3_57, 
         OutputImg3_56, OutputImg3_55, OutputImg3_54, OutputImg3_53, 
         OutputImg3_52, OutputImg3_51, OutputImg3_50, OutputImg3_49, 
         OutputImg3_48, OutputImg3_47, OutputImg3_46, OutputImg3_45, 
         OutputImg3_44, OutputImg3_43, OutputImg3_42, OutputImg3_41, 
         OutputImg3_40, OutputImg3_39, OutputImg3_38, OutputImg3_37, 
         OutputImg3_36, OutputImg3_35, OutputImg3_34, OutputImg3_33, 
         OutputImg3_32, OutputImg3_31, OutputImg3_30, OutputImg3_29, 
         OutputImg3_28, OutputImg3_27, OutputImg3_26, OutputImg3_25, 
         OutputImg3_24, OutputImg3_23, OutputImg3_22, OutputImg3_21, 
         OutputImg3_20, OutputImg3_19, OutputImg3_18, OutputImg3_17, 
         OutputImg3_16, OutputImg3_15, OutputImg3_14, OutputImg3_13, 
         OutputImg3_12, OutputImg3_11, OutputImg3_10, OutputImg3_9, OutputImg3_8, 
         OutputImg3_7, OutputImg3_6, OutputImg3_5, OutputImg3_4, OutputImg3_3, 
         OutputImg3_2, OutputImg3_1, OutputImg3_0, OutputImg4_79, OutputImg4_78, 
         OutputImg4_77, OutputImg4_76, OutputImg4_75, OutputImg4_74, 
         OutputImg4_73, OutputImg4_72, OutputImg4_71, OutputImg4_70, 
         OutputImg4_69, OutputImg4_68, OutputImg4_67, OutputImg4_66, 
         OutputImg4_65, OutputImg4_64, OutputImg4_63, OutputImg4_62, 
         OutputImg4_61, OutputImg4_60, OutputImg4_59, OutputImg4_58, 
         OutputImg4_57, OutputImg4_56, OutputImg4_55, OutputImg4_54, 
         OutputImg4_53, OutputImg4_52, OutputImg4_51, OutputImg4_50, 
         OutputImg4_49, OutputImg4_48, OutputImg4_47, OutputImg4_46, 
         OutputImg4_45, OutputImg4_44, OutputImg4_43, OutputImg4_42, 
         OutputImg4_41, OutputImg4_40, OutputImg4_39, OutputImg4_38, 
         OutputImg4_37, OutputImg4_36, OutputImg4_35, OutputImg4_34, 
         OutputImg4_33, OutputImg4_32, OutputImg4_31, OutputImg4_30, 
         OutputImg4_29, OutputImg4_28, OutputImg4_27, OutputImg4_26, 
         OutputImg4_25, OutputImg4_24, OutputImg4_23, OutputImg4_22, 
         OutputImg4_21, OutputImg4_20, OutputImg4_19, OutputImg4_18, 
         OutputImg4_17, OutputImg4_16, OutputImg4_15, OutputImg4_14, 
         OutputImg4_13, OutputImg4_12, OutputImg4_11, OutputImg4_10, 
         OutputImg4_9, OutputImg4_8, OutputImg4_7, OutputImg4_6, OutputImg4_5, 
         OutputImg4_4, OutputImg4_3, OutputImg4_2, OutputImg4_1, OutputImg4_0, 
         ConvOuput_15, ConvOuput_14, ConvOuput_13, ConvOuput_12, ConvOuput_11, 
         ConvOuput_10, ConvOuput_9, ConvOuput_8, ConvOuput_7, ConvOuput_6, 
         ConvOuput_5, ConvOuput_4, ConvOuput_3, ConvOuput_2, ConvOuput_1, 
         ConvOuput_0, ShiftLeftCounterOutput_4, ShiftLeftCounterOutput_3, 
         ShiftLeftCounterOutput_2, ShiftLeftCounterOutput_1, 
         ShiftLeftCounterOutput_0, RealOutputCounter_12, RealOutputCounter_11, 
         RealOutputCounter_10, RealOutputCounter_9, RealOutputCounter_8, 
         RealOutputCounter_7, RealOutputCounter_6, RealOutputCounter_5, 
         RealOutputCounter_4, RealOutputCounter_3, RealOutputCounter_2, 
         RealOutputCounter_1, RealOutputCounter_0, OutputCounterLoad_12, 
         OutputCounterLoad_11, OutputCounterLoad_10, OutputCounterLoad_9, 
         OutputCounterLoad_8, OutputCounterLoad_7, OutputCounterLoad_6, 
         OutputCounterLoad_5, OutputCounterLoad_4, OutputCounterLoad_3, 
         OutputCounterLoad_2, OutputCounterLoad_1, OutputCounterLoad_0, Q, 
         NumOfFilters_3, NumOfFilters_2, NumOfFilters_1, NumOfFilters_0, 
         NumOfHeight_4, NumOfHeight_3, NumOfHeight_2, NumOfHeight_1, 
         NumOfHeight_0, X, Y, K, L, D, CNDepthoutput_3, CNDepthoutput_2, 
         CNDepthoutput_1, CNDepthoutput_0, SwitchMEM_0, SwitchBar_0, CLK, 
         DontRstIndicator, lastFilter, lastDepthOut, SwitchClk, 
         TriStateCounterEN, FilterAddressEN, ImgAddRegEN, ShiftCounterRst, 
         AddressChangerEN, TriChnagerToaddEN, ImgAddRST, ramSelector, zero_11, 
         PWR, next_state_5, next_state_14, next_state_dup_134, NOT_L, 
         next_state_13, next_state_12, next_state_11, nx18, nx20, next_state_10, 
         next_state_9, next_state_dup_124, next_state_8, next_state_7, 
         next_state_dup_96, nx48, next_state_6, nx9711, nx66, next_state_3, 
         next_state_2, next_state_dup_26, NOT_nx0, next_state_1, 
         next_state_dup_147, nx100, nx112, nx130, nx142, nx154, SaveAckLatch, 
         nx180, nx186, nx9063, nx210, nx224, nx240, nx256, nx270, nx300, 
         next_state_4, next_state_dup_24, nx322, nx350, nx382, nx416, nx418, 
         nx456, nx466, nx478, nx480, nx482, nx494, nx9718, nx9728, nx9738, 
         nx9748, nx9760, nx9765, nx9768, nx9780, nx9792, nx9796, nx9814, nx9822, 
         nx9824, nx9826, nx9833, nx9835, nx9849, nx9854, nx9856, nx9858, nx9866, 
         nx9870, nx9875, nx9879, nx9881, nx9883, nx9885, nx9887, nx9889, nx9891, 
         nx9893, nx9899, nx9901, nx9903, nx9905, nx9908, nx9911, nx9913, nx9916, 
         nx9921, nx9923, nx9925, nx9932, nx9934, nx9937, nx9939, nx9941, nx9950, 
         nx9952, nx9954, nx9956, nx9958, nx9960, nx9962, nx9964, nx9966, nx9968, 
         nx9970, nx9972, nx9974, nx9976, nx9978, nx9980, nx9982, nx9984, nx9986, 
         nx9988, nx9990, nx9992, nx9994, nx9996, nx9998, nx10000, nx10002, 
         nx10004, nx10006, nx10008, nx10010, nx10012, nx10014, nx10016, nx10018, 
         nx10020, nx10022, nx10024, nx10026, nx10028, nx10032, nx10034, nx10036, 
         nx10038, nx10040, nx10042, nx10044, nx10046, nx10048, nx10050, nx10052, 
         nx10054, nx10056, nx10058, nx10060, nx10062, nx10064, nx10066, nx10068, 
         nx10070, nx10072, nx10074, nx10076, nx10078, nx10080, nx10082, nx10084, 
         nx10086, nx10088, nx10090, nx10092, nx10094, nx10096, nx10098, nx10100, 
         nx10102, nx10104, nx10106, nx10108, nx10110, nx10112, nx10114, nx10116, 
         nx10118, nx10120, nx10122, nx10124, nx10126, nx10128, nx10130, nx10132, 
         nx10134, nx10136, nx10138, nx10140, nx10142, nx10144, nx10146, nx10148, 
         nx10150, nx10152, nx10154, nx10156, nx10158, nx10160, nx10162, nx10164, 
         nx10166, nx10168, nx10170, nx10172, nx10174, nx10176, nx10178, nx10180, 
         nx10182, nx10184, nx10186, nx10188, nx10190, nx10192, nx10194, nx10196, 
         nx10198, nx10200, nx10202, nx10204, nx10206, nx10208, nx10210, nx10212, 
         nx10214, nx10216, nx10218, nx10220, nx10222, nx10224, nx10226, nx10228, 
         nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, nx10242, nx10244, 
         nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, nx10260, 
         nx10262, nx10264, nx10266, nx10268, nx10270, nx10272, nx10274, nx10276, 
         nx10278, nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, 
         nx10294, nx10296, nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, 
         nx10310, nx10312, nx10314, nx10316, nx10318, nx10320, nx10322, nx10324, 
         nx10326, nx10328, nx10330, nx10332, nx10334, nx10336, nx10338, nx10340, 
         nx10342, nx10344, nx10346, nx10348, nx10350, nx10352, nx10354, nx10356, 
         nx10358, nx10360, nx10362, nx10364, nx10366, nx10368, nx10370, nx10372, 
         nx10374, nx10376, nx10378, nx10380, nx10382, nx10384, nx10386, nx10388, 
         nx10390, nx10392, nx10394, nx10396, nx10398, nx10400, nx10402, nx10404, 
         nx10406, nx10408, nx10410, nx10412, nx10414, nx10416, nx10418, nx10420, 
         nx10422, nx10424, nx10426, nx10428, nx10430, nx10432, nx10434, nx10436, 
         nx10438, nx10440, nx10442, nx10444, nx10446, nx10448, nx10450, nx10452, 
         nx10454, nx10456, nx10458, nx10460, nx10462, nx10464, nx10466, nx10468, 
         nx10470, nx10472, nx10474, nx10476, nx10478, nx10484, nx10486, nx10488, 
         nx10490, nx10496, nx10498, nx5, nx10500, nx10502, nx10504;
    wire [2746:0] \$dummy ;




    nBitRegister_1 DDF0 (.D ({SwitchBar_0}), .CLK (SwitchClk), .RST (rst), .EN (
                   PWR), .Q ({SwitchMEM_0})) ;
    triStateBuffer_13 TriStateAddchanger (.D ({nx9974,nx9978,nx9982,nx9986,
                      nx9990,nx9994,nx9998,nx10002,nx10006,nx10010,nx10014,
                      nx10018,nx10022}), .EN (nx9958), .F ({AddressChangerIN_12,
                      AddressChangerIN_11,AddressChangerIN_10,AddressChangerIN_9
                      ,AddressChangerIN_8,AddressChangerIN_7,AddressChangerIN_6,
                      AddressChangerIN_5,AddressChangerIN_4,AddressChangerIN_3,
                      AddressChangerIN_2,AddressChangerIN_1,AddressChangerIN_0})
                      ) ;
    triStateBuffer_13 TriStateAddgfd (.D ({AddressChangerOut_12,
                      AddressChangerOut_11,AddressChangerOut_10,
                      AddressChangerOut_9,AddressChangerOut_8,
                      AddressChangerOut_7,AddressChangerOut_6,
                      AddressChangerOut_5,AddressChangerOut_4,
                      AddressChangerOut_3,AddressChangerOut_2,
                      AddressChangerOut_1,AddressChangerOut_0}), .EN (
                      TriChnagerToaddEN), .F ({FilterAddressIN_12,
                      FilterAddressIN_11,FilterAddressIN_10,FilterAddressIN_9,
                      FilterAddressIN_8,FilterAddressIN_7,FilterAddressIN_6,
                      FilterAddressIN_5,FilterAddressIN_4,FilterAddressIN_3,
                      FilterAddressIN_2,FilterAddressIN_1,FilterAddressIN_0})) ;
    nBitRegister_13 addChanger (.D ({AddressChangerIN_12,AddressChangerIN_11,
                    AddressChangerIN_10,AddressChangerIN_9,AddressChangerIN_8,
                    AddressChangerIN_7,AddressChangerIN_6,AddressChangerIN_5,
                    AddressChangerIN_4,AddressChangerIN_3,AddressChangerIN_2,
                    AddressChangerIN_1,AddressChangerIN_0}), .CLK (nx10414), .RST (
                    rst), .EN (AddressChangerEN), .Q ({AddressChangerOut_12,
                    AddressChangerOut_11,AddressChangerOut_10,
                    AddressChangerOut_9,AddressChangerOut_8,AddressChangerOut_7,
                    AddressChangerOut_6,AddressChangerOut_5,AddressChangerOut_4,
                    AddressChangerOut_3,AddressChangerOut_2,AddressChangerOut_1,
                    AddressChangerOut_0})) ;
    RAM_25 FilterMem (.reset (rst), .CLK (nx10414), .W (zero_11), .R (ReadF), .address (
           {AddressF_12,AddressF_11,AddressF_10,AddressF_9,AddressF_8,AddressF_7
           ,AddressF_6,AddressF_5,AddressF_4,AddressF_3,AddressF_2,AddressF_1,
           AddressF_0}), .dataIn ({zero_11,zero_11,zero_11,zero_11,zero_11,
           zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
           zero_11,zero_11,zero_11}), .dataOut ({DataFOut_399,\$dummy [0],
           \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
           \$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],
           \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],\$dummy [15],
           \$dummy [16],\$dummy [17],\$dummy [18],\$dummy [19],\$dummy [20],
           \$dummy [21],\$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],
           \$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],\$dummy [30],
           \$dummy [31],\$dummy [32],\$dummy [33],\$dummy [34],\$dummy [35],
           \$dummy [36],\$dummy [37],\$dummy [38],\$dummy [39],\$dummy [40],
           \$dummy [41],\$dummy [42],\$dummy [43],\$dummy [44],\$dummy [45],
           \$dummy [46],\$dummy [47],\$dummy [48],\$dummy [49],\$dummy [50],
           \$dummy [51],\$dummy [52],\$dummy [53],\$dummy [54],\$dummy [55],
           \$dummy [56],\$dummy [57],\$dummy [58],\$dummy [59],\$dummy [60],
           \$dummy [61],\$dummy [62],\$dummy [63],\$dummy [64],\$dummy [65],
           \$dummy [66],\$dummy [67],\$dummy [68],\$dummy [69],\$dummy [70],
           \$dummy [71],\$dummy [72],\$dummy [73],\$dummy [74],\$dummy [75],
           \$dummy [76],\$dummy [77],\$dummy [78],\$dummy [79],\$dummy [80],
           \$dummy [81],\$dummy [82],\$dummy [83],\$dummy [84],\$dummy [85],
           \$dummy [86],\$dummy [87],\$dummy [88],\$dummy [89],\$dummy [90],
           \$dummy [91],\$dummy [92],\$dummy [93],\$dummy [94],\$dummy [95],
           \$dummy [96],\$dummy [97],\$dummy [98],\$dummy [99],\$dummy [100],
           \$dummy [101],\$dummy [102],\$dummy [103],\$dummy [104],\$dummy [105]
           ,\$dummy [106],\$dummy [107],\$dummy [108],\$dummy [109],
           \$dummy [110],\$dummy [111],\$dummy [112],\$dummy [113],\$dummy [114]
           ,\$dummy [115],\$dummy [116],\$dummy [117],\$dummy [118],
           \$dummy [119],\$dummy [120],\$dummy [121],\$dummy [122],\$dummy [123]
           ,\$dummy [124],\$dummy [125],\$dummy [126],\$dummy [127],
           \$dummy [128],\$dummy [129],\$dummy [130],\$dummy [131],\$dummy [132]
           ,\$dummy [133],\$dummy [134],\$dummy [135],\$dummy [136],
           \$dummy [137],\$dummy [138],\$dummy [139],\$dummy [140],\$dummy [141]
           ,\$dummy [142],\$dummy [143],\$dummy [144],\$dummy [145],
           \$dummy [146],\$dummy [147],\$dummy [148],\$dummy [149],\$dummy [150]
           ,\$dummy [151],\$dummy [152],\$dummy [153],\$dummy [154],
           \$dummy [155],\$dummy [156],\$dummy [157],\$dummy [158],\$dummy [159]
           ,\$dummy [160],\$dummy [161],\$dummy [162],\$dummy [163],
           \$dummy [164],\$dummy [165],\$dummy [166],\$dummy [167],\$dummy [168]
           ,\$dummy [169],\$dummy [170],\$dummy [171],\$dummy [172],
           \$dummy [173],\$dummy [174],\$dummy [175],\$dummy [176],\$dummy [177]
           ,\$dummy [178],\$dummy [179],\$dummy [180],\$dummy [181],
           \$dummy [182],\$dummy [183],\$dummy [184],\$dummy [185],\$dummy [186]
           ,\$dummy [187],\$dummy [188],\$dummy [189],\$dummy [190],
           \$dummy [191],\$dummy [192],\$dummy [193],\$dummy [194],\$dummy [195]
           ,\$dummy [196],\$dummy [197],\$dummy [198],\$dummy [199],
           \$dummy [200],\$dummy [201],\$dummy [202],\$dummy [203],\$dummy [204]
           ,\$dummy [205],\$dummy [206],\$dummy [207],\$dummy [208],
           \$dummy [209],\$dummy [210],\$dummy [211],\$dummy [212],\$dummy [213]
           ,\$dummy [214],\$dummy [215],\$dummy [216],\$dummy [217],
           \$dummy [218],\$dummy [219],\$dummy [220],\$dummy [221],\$dummy [222]
           ,\$dummy [223],\$dummy [224],\$dummy [225],\$dummy [226],
           \$dummy [227],\$dummy [228],\$dummy [229],\$dummy [230],\$dummy [231]
           ,\$dummy [232],\$dummy [233],\$dummy [234],\$dummy [235],
           \$dummy [236],\$dummy [237],\$dummy [238],\$dummy [239],\$dummy [240]
           ,\$dummy [241],\$dummy [242],\$dummy [243],\$dummy [244],
           \$dummy [245],\$dummy [246],\$dummy [247],\$dummy [248],\$dummy [249]
           ,\$dummy [250],\$dummy [251],\$dummy [252],\$dummy [253],
           \$dummy [254],\$dummy [255],\$dummy [256],\$dummy [257],\$dummy [258]
           ,\$dummy [259],\$dummy [260],\$dummy [261],\$dummy [262],
           \$dummy [263],\$dummy [264],\$dummy [265],\$dummy [266],\$dummy [267]
           ,\$dummy [268],\$dummy [269],\$dummy [270],\$dummy [271],
           \$dummy [272],\$dummy [273],\$dummy [274],\$dummy [275],\$dummy [276]
           ,\$dummy [277],\$dummy [278],\$dummy [279],\$dummy [280],
           \$dummy [281],\$dummy [282],\$dummy [283],\$dummy [284],\$dummy [285]
           ,\$dummy [286],\$dummy [287],\$dummy [288],\$dummy [289],
           \$dummy [290],\$dummy [291],\$dummy [292],\$dummy [293],\$dummy [294]
           ,\$dummy [295],\$dummy [296],\$dummy [297],\$dummy [298],
           \$dummy [299],\$dummy [300],\$dummy [301],\$dummy [302],\$dummy [303]
           ,\$dummy [304],\$dummy [305],\$dummy [306],\$dummy [307],
           \$dummy [308],\$dummy [309],\$dummy [310],\$dummy [311],\$dummy [312]
           ,\$dummy [313],\$dummy [314],\$dummy [315],\$dummy [316],
           \$dummy [317],\$dummy [318],\$dummy [319],\$dummy [320],\$dummy [321]
           ,\$dummy [322],\$dummy [323],\$dummy [324],\$dummy [325],
           \$dummy [326],\$dummy [327],\$dummy [328],\$dummy [329],\$dummy [330]
           ,\$dummy [331],\$dummy [332],\$dummy [333],\$dummy [334],
           \$dummy [335],\$dummy [336],\$dummy [337],\$dummy [338],\$dummy [339]
           ,\$dummy [340],\$dummy [341],\$dummy [342],\$dummy [343],
           \$dummy [344],\$dummy [345],\$dummy [346],\$dummy [347],\$dummy [348]
           ,\$dummy [349],\$dummy [350],\$dummy [351],\$dummy [352],
           \$dummy [353],\$dummy [354],\$dummy [355],\$dummy [356],\$dummy [357]
           ,\$dummy [358],\$dummy [359],\$dummy [360],\$dummy [361],
           \$dummy [362],\$dummy [363],\$dummy [364],\$dummy [365],\$dummy [366]
           ,\$dummy [367],\$dummy [368],\$dummy [369],\$dummy [370],
           \$dummy [371],\$dummy [372],\$dummy [373],\$dummy [374],\$dummy [375]
           ,\$dummy [376],\$dummy [377],\$dummy [378],\$dummy [379],
           \$dummy [380],\$dummy [381],\$dummy [382],\$dummy [383],\$dummy [384]
           ,\$dummy [385],\$dummy [386],\$dummy [387],\$dummy [388],
           \$dummy [389],\$dummy [390],\$dummy [391],\$dummy [392],\$dummy [393]
           ,\$dummy [394],\$dummy [395],\$dummy [396],\$dummy [397],
           \$dummy [398]}), .MFC (ACKF), .counterOut ({\$dummy [399],
           \$dummy [400],\$dummy [401],\$dummy [402]})) ;
    memoryDMA ImgMem (.resetEN (rst), .AddressIn ({AddressI_12,AddressI_11,
              AddressI_10,AddressI_9,AddressI_8,AddressI_7,AddressI_6,AddressI_5
              ,AddressI_4,AddressI_3,AddressI_2,AddressI_1,AddressI_0}), .dataIn (
              {DataIIn_15,DataIIn_14,DataIIn_13,DataIIn_12,DataIIn_11,DataIIn_10
              ,DataIIn_9,DataIIn_8,DataIIn_7,DataIIn_6,DataIIn_5,DataIIn_4,
              DataIIn_3,DataIIn_2,DataIIn_1,DataIIn_0}), .switcherEN (
              SwitchMEM_0), .ramSelector (ramSelector), .readEn (ReadI), .writeEn (
              WriteI), .CLK (nx10416), .Normal (zero_11), .MFC (ImgAddACKTriIN_0
              ), .counterOut ({\$dummy [403],\$dummy [404],\$dummy [405],
              \$dummy [406]}), .dataOut ({DataIOut_447,DataIOut_446,DataIOut_445
              ,DataIOut_444,DataIOut_443,DataIOut_442,DataIOut_441,DataIOut_440,
              DataIOut_439,DataIOut_438,DataIOut_437,DataIOut_436,DataIOut_435,
              DataIOut_434,DataIOut_433,DataIOut_432,DataIOut_431,DataIOut_430,
              DataIOut_429,DataIOut_428,DataIOut_427,DataIOut_426,DataIOut_425,
              DataIOut_424,DataIOut_423,DataIOut_422,DataIOut_421,DataIOut_420,
              DataIOut_419,DataIOut_418,DataIOut_417,DataIOut_416,DataIOut_415,
              DataIOut_414,DataIOut_413,DataIOut_412,DataIOut_411,DataIOut_410,
              DataIOut_409,DataIOut_408,DataIOut_407,DataIOut_406,DataIOut_405,
              DataIOut_404,DataIOut_403,DataIOut_402,DataIOut_401,DataIOut_400,
              DataIOut_399,DataIOut_398,DataIOut_397,DataIOut_396,DataIOut_395,
              DataIOut_394,DataIOut_393,DataIOut_392,DataIOut_391,DataIOut_390,
              DataIOut_389,DataIOut_388,DataIOut_387,DataIOut_386,DataIOut_385,
              DataIOut_384,DataIOut_383,DataIOut_382,DataIOut_381,DataIOut_380,
              DataIOut_379,DataIOut_378,DataIOut_377,DataIOut_376,DataIOut_375,
              DataIOut_374,DataIOut_373,DataIOut_372,DataIOut_371,DataIOut_370,
              DataIOut_369,DataIOut_368,DataIOut_367,DataIOut_366,DataIOut_365,
              DataIOut_364,DataIOut_363,DataIOut_362,DataIOut_361,DataIOut_360,
              DataIOut_359,DataIOut_358,DataIOut_357,DataIOut_356,DataIOut_355,
              DataIOut_354,DataIOut_353,DataIOut_352,DataIOut_351,DataIOut_350,
              DataIOut_349,DataIOut_348,DataIOut_347,DataIOut_346,DataIOut_345,
              DataIOut_344,DataIOut_343,DataIOut_342,DataIOut_341,DataIOut_340,
              DataIOut_339,DataIOut_338,DataIOut_337,DataIOut_336,DataIOut_335,
              DataIOut_334,DataIOut_333,DataIOut_332,DataIOut_331,DataIOut_330,
              DataIOut_329,DataIOut_328,DataIOut_327,DataIOut_326,DataIOut_325,
              DataIOut_324,DataIOut_323,DataIOut_322,DataIOut_321,DataIOut_320,
              DataIOut_319,DataIOut_318,DataIOut_317,DataIOut_316,DataIOut_315,
              DataIOut_314,DataIOut_313,DataIOut_312,DataIOut_311,DataIOut_310,
              DataIOut_309,DataIOut_308,DataIOut_307,DataIOut_306,DataIOut_305,
              DataIOut_304,DataIOut_303,DataIOut_302,DataIOut_301,DataIOut_300,
              DataIOut_299,DataIOut_298,DataIOut_297,DataIOut_296,DataIOut_295,
              DataIOut_294,DataIOut_293,DataIOut_292,DataIOut_291,DataIOut_290,
              DataIOut_289,DataIOut_288,DataIOut_287,DataIOut_286,DataIOut_285,
              DataIOut_284,DataIOut_283,DataIOut_282,DataIOut_281,DataIOut_280,
              DataIOut_279,DataIOut_278,DataIOut_277,DataIOut_276,DataIOut_275,
              DataIOut_274,DataIOut_273,DataIOut_272,DataIOut_271,DataIOut_270,
              DataIOut_269,DataIOut_268,DataIOut_267,DataIOut_266,DataIOut_265,
              DataIOut_264,DataIOut_263,DataIOut_262,DataIOut_261,DataIOut_260,
              DataIOut_259,DataIOut_258,DataIOut_257,DataIOut_256,DataIOut_255,
              DataIOut_254,DataIOut_253,DataIOut_252,DataIOut_251,DataIOut_250,
              DataIOut_249,DataIOut_248,DataIOut_247,DataIOut_246,DataIOut_245,
              DataIOut_244,DataIOut_243,DataIOut_242,DataIOut_241,DataIOut_240,
              DataIOut_239,DataIOut_238,DataIOut_237,DataIOut_236,DataIOut_235,
              DataIOut_234,DataIOut_233,DataIOut_232,DataIOut_231,DataIOut_230,
              DataIOut_229,DataIOut_228,DataIOut_227,DataIOut_226,DataIOut_225,
              DataIOut_224,DataIOut_223,DataIOut_222,DataIOut_221,DataIOut_220,
              DataIOut_219,DataIOut_218,DataIOut_217,DataIOut_216,DataIOut_215,
              DataIOut_214,DataIOut_213,DataIOut_212,DataIOut_211,DataIOut_210,
              DataIOut_209,DataIOut_208,DataIOut_207,DataIOut_206,DataIOut_205,
              DataIOut_204,DataIOut_203,DataIOut_202,DataIOut_201,DataIOut_200,
              DataIOut_199,DataIOut_198,DataIOut_197,DataIOut_196,DataIOut_195,
              DataIOut_194,DataIOut_193,DataIOut_192,DataIOut_191,DataIOut_190,
              DataIOut_189,DataIOut_188,DataIOut_187,DataIOut_186,DataIOut_185,
              DataIOut_184,DataIOut_183,DataIOut_182,DataIOut_181,DataIOut_180,
              DataIOut_179,DataIOut_178,DataIOut_177,DataIOut_176,DataIOut_175,
              DataIOut_174,DataIOut_173,DataIOut_172,DataIOut_171,DataIOut_170,
              DataIOut_169,DataIOut_168,DataIOut_167,DataIOut_166,DataIOut_165,
              DataIOut_164,DataIOut_163,DataIOut_162,DataIOut_161,DataIOut_160,
              DataIOut_159,DataIOut_158,DataIOut_157,DataIOut_156,DataIOut_155,
              DataIOut_154,DataIOut_153,DataIOut_152,DataIOut_151,DataIOut_150,
              DataIOut_149,DataIOut_148,DataIOut_147,DataIOut_146,DataIOut_145,
              DataIOut_144,DataIOut_143,DataIOut_142,DataIOut_141,DataIOut_140,
              DataIOut_139,DataIOut_138,DataIOut_137,DataIOut_136,DataIOut_135,
              DataIOut_134,DataIOut_133,DataIOut_132,DataIOut_131,DataIOut_130,
              DataIOut_129,DataIOut_128,DataIOut_127,DataIOut_126,DataIOut_125,
              DataIOut_124,DataIOut_123,DataIOut_122,DataIOut_121,DataIOut_120,
              DataIOut_119,DataIOut_118,DataIOut_117,DataIOut_116,DataIOut_115,
              DataIOut_114,DataIOut_113,DataIOut_112,DataIOut_111,DataIOut_110,
              DataIOut_109,DataIOut_108,DataIOut_107,DataIOut_106,DataIOut_105,
              DataIOut_104,DataIOut_103,DataIOut_102,DataIOut_101,DataIOut_100,
              DataIOut_99,DataIOut_98,DataIOut_97,DataIOut_96,DataIOut_95,
              DataIOut_94,DataIOut_93,DataIOut_92,DataIOut_91,DataIOut_90,
              DataIOut_89,DataIOut_88,DataIOut_87,DataIOut_86,DataIOut_85,
              DataIOut_84,DataIOut_83,DataIOut_82,DataIOut_81,DataIOut_80,
              DataIOut_79,DataIOut_78,DataIOut_77,DataIOut_76,DataIOut_75,
              DataIOut_74,DataIOut_73,DataIOut_72,DataIOut_71,DataIOut_70,
              DataIOut_69,DataIOut_68,DataIOut_67,DataIOut_66,DataIOut_65,
              DataIOut_64,DataIOut_63,DataIOut_62,DataIOut_61,DataIOut_60,
              DataIOut_59,DataIOut_58,DataIOut_57,DataIOut_56,DataIOut_55,
              DataIOut_54,DataIOut_53,DataIOut_52,DataIOut_51,DataIOut_50,
              DataIOut_49,DataIOut_48,DataIOut_47,DataIOut_46,DataIOut_45,
              DataIOut_44,DataIOut_43,DataIOut_42,DataIOut_41,DataIOut_40,
              DataIOut_39,DataIOut_38,DataIOut_37,DataIOut_36,DataIOut_35,
              DataIOut_34,DataIOut_33,DataIOut_32,DataIOut_31,DataIOut_30,
              DataIOut_29,DataIOut_28,DataIOut_27,DataIOut_26,DataIOut_25,
              DataIOut_24,DataIOut_23,DataIOut_22,DataIOut_21,DataIOut_20,
              DataIOut_19,DataIOut_18,DataIOut_17,DataIOut_16,DataIOut_15,
              DataIOut_14,DataIOut_13,DataIOut_12,DataIOut_11,DataIOut_10,
              DataIOut_9,DataIOut_8,DataIOut_7,DataIOut_6,DataIOut_5,DataIOut_4,
              DataIOut_3,DataIOut_2,DataIOut_1,DataIOut_0})) ;
    ReadInfoState ReadInf (.CLK (nx10418), .S ({zero_11,zero_11,zero_11,zero_11,
                  zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                  zero_11,zero_11,zero_11,current_state_0}), .reset (rst), .MFC (
                  zero_11), .filterAddressReg_out ({nx9974,nx9978,nx9982,nx9986,
                  nx9990,nx9994,nx9998,nx10002,nx10006,nx10010,nx10014,nx10018,
                  nx10022}), .filterRamData ({nx10256,nx10262,nx10268,nx10274,
                  nx10280,nx10286,nx10292,nx10292,nx10294,nx10294,nx10296,
                  nx10298,nx10300,nx10302,nx10302,nx10304}), .noOfLayersReg_out (
                  {\$dummy [407],\$dummy [408],\$dummy [409],\$dummy [410],
                  \$dummy [411],\$dummy [412],\$dummy [413],\$dummy [414],
                  \$dummy [415],\$dummy [416],\$dummy [417],\$dummy [418],
                  \$dummy [419],\$dummy [420],NoOfLayers_1,NoOfLayers_0}), .filterRamAddress (
                  {AddressF_12,AddressF_11,AddressF_10,AddressF_9,AddressF_8,
                  AddressF_7,AddressF_6,AddressF_5,AddressF_4,AddressF_3,
                  AddressF_2,AddressF_1,AddressF_0})) ;
    nBitRegister_13 FilterAddress (.D ({FilterAddressIN_12,FilterAddressIN_11,
                    FilterAddressIN_10,FilterAddressIN_9,FilterAddressIN_8,
                    FilterAddressIN_7,FilterAddressIN_6,FilterAddressIN_5,
                    FilterAddressIN_4,FilterAddressIN_3,FilterAddressIN_2,
                    FilterAddressIN_1,FilterAddressIN_0}), .CLK (nx10414), .RST (
                    rst), .EN (FilterAddressEN), .Q ({FilterAddressOut_12,
                    FilterAddressOut_11,FilterAddressOut_10,FilterAddressOut_9,
                    FilterAddressOut_8,FilterAddressOut_7,FilterAddressOut_6,
                    FilterAddressOut_5,FilterAddressOut_4,FilterAddressOut_3,
                    FilterAddressOut_2,FilterAddressOut_1,FilterAddressOut_0})
                    ) ;
    triStateBuffer_13 AdderTryState (.D ({TriStateCounterOUT_12,
                      TriStateCounterOUT_11,TriStateCounterOUT_10,
                      TriStateCounterOUT_9,TriStateCounterOUT_8,
                      TriStateCounterOUT_7,TriStateCounterOUT_6,
                      TriStateCounterOUT_5,TriStateCounterOUT_4,
                      TriStateCounterOUT_3,TriStateCounterOUT_2,
                      TriStateCounterOUT_1,TriStateCounterOUT_0}), .EN (
                      TriStateCounterEN), .F ({FilterAddressIN_12,
                      FilterAddressIN_11,FilterAddressIN_10,FilterAddressIN_9,
                      FilterAddressIN_8,FilterAddressIN_7,FilterAddressIN_6,
                      FilterAddressIN_5,FilterAddressIN_4,FilterAddressIN_3,
                      FilterAddressIN_2,FilterAddressIN_1,FilterAddressIN_0})) ;
    my_nadder_13 FilterAddressAdder (.a ({nx9974,nx9978,nx9982,nx9986,nx9990,
                 nx9994,nx9998,nx10002,nx10006,nx10010,nx10014,nx10018,nx10022})
                 , .b ({zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                 zero_11,zero_11,zero_11,zero_11,zero_11,zero_11}), .cin (PWR), 
                 .s ({TriStateCounterOUT_12,TriStateCounterOUT_11,
                 TriStateCounterOUT_10,TriStateCounterOUT_9,TriStateCounterOUT_8
                 ,TriStateCounterOUT_7,TriStateCounterOUT_6,TriStateCounterOUT_5
                 ,TriStateCounterOUT_4,TriStateCounterOUT_3,TriStateCounterOUT_2
                 ,TriStateCounterOUT_1,TriStateCounterOUT_0}), .cout (
                 \$dummy [421])) ;
    nBitRegister_13 ImgAddReg (.D ({ImgAddRegIN_12,ImgAddRegIN_11,ImgAddRegIN_10
                    ,ImgAddRegIN_9,ImgAddRegIN_8,ImgAddRegIN_7,ImgAddRegIN_6,
                    ImgAddRegIN_5,ImgAddRegIN_4,ImgAddRegIN_3,ImgAddRegIN_2,
                    ImgAddRegIN_1,ImgAddRegIN_0}), .CLK (nx10418), .RST (
                    ImgAddRST), .EN (ImgAddRegEN), .Q ({ImgAddRegOut_12,
                    ImgAddRegOut_11,ImgAddRegOut_10,ImgAddRegOut_9,
                    ImgAddRegOut_8,ImgAddRegOut_7,ImgAddRegOut_6,ImgAddRegOut_5,
                    ImgAddRegOut_4,ImgAddRegOut_3,ImgAddRegOut_2,ImgAddRegOut_1,
                    ImgAddRegOut_0})) ;
    triStateBuffer_13 ImgAddACKTri (.D ({zero_11,zero_11,zero_11,zero_11,zero_11
                      ,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                      nx10026}), .EN (nx9972), .F ({ImgAddRegIN_12,
                      ImgAddRegIN_11,ImgAddRegIN_10,ImgAddRegIN_9,ImgAddRegIN_8,
                      ImgAddRegIN_7,ImgAddRegIN_6,ImgAddRegIN_5,ImgAddRegIN_4,
                      ImgAddRegIN_3,ImgAddRegIN_2,ImgAddRegIN_1,ImgAddRegIN_0})
                      ) ;
    ReadLayerInfo ReadLayerInfo (.LayerInfoIn ({nx10258,nx10264,nx10270,nx10276,
                  nx10282,nx10288,nx10292,nx10292,nx10294,nx10296,nx10298,
                  nx10298,nx10300,nx10302,nx10302,nx10304}), .ImgWidthIn ({
                  nx10312,nx10316,nx10320,nx10324,nx10328,nx10332,nx10336,
                  nx10340,nx10344,nx10348,nx10352,nx10356,nx10360,nx10364,
                  nx10368,nx10372}), .FilterAdd ({nx9974,nx9978,nx9982,nx9986,
                  nx9990,nx9994,nx9998,nx10002,nx10006,nx10010,nx10014,nx10018,
                  nx10022}), .ImgAdd ({ImgAddRegOut_12,ImgAddRegOut_11,
                  ImgAddRegOut_10,ImgAddRegOut_9,ImgAddRegOut_8,ImgAddRegOut_7,
                  ImgAddRegOut_6,ImgAddRegOut_5,ImgAddRegOut_4,ImgAddRegOut_3,
                  ImgAddRegOut_2,ImgAddRegOut_1,ImgAddRegOut_0}), .clk (nx10420)
                  , .rst (rst), .ACKF (nx10308), .ACKI (nx10026), .current_state (
                  {zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                  zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,nx9970,zero_11
                  }), .LayerInfoOut ({LayerInfoOut_15,LayerInfoOut_14,
                  \$dummy [422],LayerInfoOut_12,LayerInfoOut_11,LayerInfoOut_10,
                  LayerInfoOut_9,LayerInfoOut_8,LayerInfoOut_7,LayerInfoOut_6,
                  LayerInfoOut_5,LayerInfoOut_4,LayerInfoOut_3,LayerInfoOut_2,
                  LayerInfoOut_1,LayerInfoOut_0}), .ImgWidthOut ({ImgWidthOut_15
                  ,ImgWidthOut_14,ImgWidthOut_13,ImgWidthOut_12,ImgWidthOut_11,
                  ImgWidthOut_10,ImgWidthOut_9,ImgWidthOut_8,ImgWidthOut_7,
                  ImgWidthOut_6,ImgWidthOut_5,ImgWidthOut_4,ImgWidthOut_3,
                  ImgWidthOut_2,ImgWidthOut_1,ImgWidthOut_0}), .FilterAddToDMA (
                  {AddressF_12,AddressF_11,AddressF_10,AddressF_9,AddressF_8,
                  AddressF_7,AddressF_6,AddressF_5,AddressF_4,AddressF_3,
                  AddressF_2,AddressF_1,AddressF_0}), .ImgAddToDMA ({AddressI_12
                  ,AddressI_11,AddressI_10,AddressI_9,AddressI_8,AddressI_7,
                  AddressI_6,AddressI_5,AddressI_4,AddressI_3,AddressI_2,
                  AddressI_1,AddressI_0})) ;
    CalculateInfo ClacInfo (.WSquareOut ({WidthSquareOut_9,WidthSquareOut_8,
                  WidthSquareOut_7,WidthSquareOut_6,WidthSquareOut_5,
                  WidthSquareOut_4,WidthSquareOut_3,WidthSquareOut_2,
                  WidthSquareOut_1,WidthSquareOut_0}), .CounOut ({\$dummy [423],
                  \$dummy [424]}), .LayerInfoIn ({zero_11,zero_11,zero_11,
                  zero_11,zero_11,zero_11,zero_11,nx10376,nx10380,nx10384,
                  nx10388,nx10392,zero_11,zero_11,zero_11,zero_11}), .clk (
                  nx10504), .rst (rst), .current_state ({zero_11,zero_11,zero_11
                  ,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                  nx9966,zero_11,current_state_2,zero_11,zero_11}), .ACK (
                  \$dummy [425]), .ACKI (nx10026), .Wmin1 ({\$dummy [426],
                  \$dummy [427],\$dummy [428],\$dummy [429],\$dummy [430]})) ;
    ReadBias RBias (.current_state ({zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,nx9968,zero_11,zero_11,
             zero_11,zero_11}), .BIAS ({zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,nx10032,nx10034,nx10036,nx10038,nx10040,
             nx10042,nx10044,nx10046,nx10048,nx10050,nx10052,nx10054,nx10056,
             nx10058,nx10060,nx10062,nx10064,nx10066,nx10068,nx10070,nx10072,
             nx10074,nx10076,nx10078,nx10080,nx10082,nx10084,nx10086,nx10088,
             nx10090,nx10092,nx10094,nx10096,nx10098,nx10100,nx10102,nx10104,
             nx10106,nx10108,nx10110,nx10112,nx10114,nx10116,nx10118,nx10120,
             nx10122,nx10124,nx10126,nx10128,nx10130,nx10132,nx10134,nx10136,
             nx10138,nx10140,nx10142,nx10144,nx10146,nx10148,nx10150,nx10152,
             nx10154,nx10156,nx10158,nx10160,nx10162,nx10164,nx10166,nx10168,
             nx10170,nx10172,nx10174,nx10176,nx10178,nx10180,nx10182,nx10184,
             nx10186,nx10188,nx10190,nx10192,nx10194,nx10196,nx10198,nx10200,
             nx10202,nx10204,nx10206,nx10208,nx10210,nx10212,nx10214,nx10216,
             nx10218,nx10220,nx10222,nx10224,nx10226,nx10228,nx10230,nx10232,
             nx10234,nx10236,nx10238,nx10240,nx10242,nx10244,nx10246,nx10248,
             nx10250,nx10252,nx10254,nx10260,nx10266,nx10272,nx10278,nx10284,
             nx10290,nx10292,nx10294,nx10294,nx10296,nx10298,nx10298,nx10300,
             nx10302,nx10304,nx10304}), .FilterAddress ({nx9976,nx9980,nx9984,
             nx9988,nx9992,nx9996,nx10000,nx10004,nx10008,nx10012,nx10016,
             nx10020,nx10024}), .DMAAddressToFilter ({AddressF_12,AddressF_11,
             AddressF_10,AddressF_9,AddressF_8,AddressF_7,AddressF_6,AddressF_5,
             AddressF_4,AddressF_3,AddressF_2,AddressF_1,AddressF_0}), .UpdatedAddress (
             {FilterAddressIN_12,FilterAddressIN_11,FilterAddressIN_10,
             FilterAddressIN_9,FilterAddressIN_8,FilterAddressIN_7,
             FilterAddressIN_6,FilterAddressIN_5,FilterAddressIN_4,
             FilterAddressIN_3,FilterAddressIN_2,FilterAddressIN_1,
             FilterAddressIN_0}), .changerAdd ({AddressChangerIN_12,
             AddressChangerIN_11,AddressChangerIN_10,AddressChangerIN_9,
             AddressChangerIN_8,AddressChangerIN_7,AddressChangerIN_6,
             AddressChangerIN_5,AddressChangerIN_4,AddressChangerIN_3,
             AddressChangerIN_2,AddressChangerIN_1,AddressChangerIN_0}), .CLK (
             nx10416), .RST (rst), .LayerInfo ({zero_11,zero_11,zero_11,zero_11,
             zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
             LayerInfoOut_3,LayerInfoOut_2,LayerInfoOut_1,LayerInfoOut_0}), .outBias0 (
             {Bias0_15,Bias0_14,Bias0_13,Bias0_12,Bias0_11,Bias0_10,Bias0_9,
             Bias0_8,Bias0_7,Bias0_6,Bias0_5,Bias0_4,Bias0_3,Bias0_2,Bias0_1,
             Bias0_0}), .outBias1 ({Bias1_15,Bias1_14,Bias1_13,Bias1_12,Bias1_11
             ,Bias1_10,Bias1_9,Bias1_8,Bias1_7,Bias1_6,Bias1_5,Bias1_4,Bias1_3,
             Bias1_2,Bias1_1,Bias1_0}), .outBias2 ({Bias2_15,Bias2_14,Bias2_13,
             Bias2_12,Bias2_11,Bias2_10,Bias2_9,Bias2_8,Bias2_7,Bias2_6,Bias2_5,
             Bias2_4,Bias2_3,Bias2_2,Bias2_1,Bias2_0}), .outBias3 ({Bias3_15,
             Bias3_14,Bias3_13,Bias3_12,Bias3_11,Bias3_10,Bias3_9,Bias3_8,
             Bias3_7,Bias3_6,Bias3_5,Bias3_4,Bias3_3,Bias3_2,Bias3_1,Bias3_0}), 
             .outBias4 ({Bias4_15,Bias4_14,Bias4_13,Bias4_12,Bias4_11,Bias4_10,
             Bias4_9,Bias4_8,Bias4_7,Bias4_6,Bias4_5,Bias4_4,Bias4_3,Bias4_2,
             Bias4_1,Bias4_0}), .outBias5 ({Bias5_15,Bias5_14,Bias5_13,Bias5_12,
             Bias5_11,Bias5_10,Bias5_9,Bias5_8,Bias5_7,Bias5_6,Bias5_5,Bias5_4,
             Bias5_3,Bias5_2,Bias5_1,Bias5_0}), .outBias6 ({Bias6_15,Bias6_14,
             Bias6_13,Bias6_12,Bias6_11,Bias6_10,Bias6_9,Bias6_8,Bias6_7,Bias6_6
             ,Bias6_5,Bias6_4,Bias6_3,Bias6_2,Bias6_1,Bias6_0}), .outBias7 ({
             Bias7_15,Bias7_14,Bias7_13,Bias7_12,Bias7_11,Bias7_10,Bias7_9,
             Bias7_8,Bias7_7,Bias7_6,Bias7_5,Bias7_4,Bias7_3,Bias7_2,Bias7_1,
             Bias7_0}), .ACKF (nx10308)) ;
    ReadFilter Rfilter (.current_state ({zero_11,zero_11,zero_11,zero_11,
               current_state_10,zero_11,zero_11,nx9962,zero_11,current_state_5,
               zero_11,zero_11,zero_11,zero_11,zero_11}), .LayerInfo ({zero_11,
               zero_11,zero_11,LayerInfoOut_12,LayerInfoOut_11,LayerInfoOut_10,
               LayerInfoOut_9,nx10378,nx10382,nx10386,nx10388,nx10392,
               LayerInfoOut_3,LayerInfoOut_2,LayerInfoOut_1,LayerInfoOut_0}), .depthcounter (
               {nx10406,nx10408,nx10410,nx10412}), .FilterCounter ({nx10398,
               nx10400,nx10402,nx10404}), .Heightcounter ({NumOfHeight_4,
               NumOfHeight_3,NumOfHeight_2,NumOfHeight_1,NumOfHeight_0}), .FILTER (
               {nx10032,nx10032,nx10032,nx10034,nx10034,nx10034,nx10036,nx10036,
               nx10036,nx10038,nx10038,nx10038,nx10040,nx10040,nx10040,nx10042,
               nx10042,nx10042,nx10044,nx10044,nx10044,nx10046,nx10046,nx10046,
               nx10048,nx10048,nx10048,nx10050,nx10050,nx10050,nx10052,nx10052,
               nx10052,nx10054,nx10054,nx10054,nx10056,nx10056,nx10056,nx10058,
               nx10058,nx10058,nx10060,nx10060,nx10060,nx10062,nx10062,nx10062,
               nx10064,nx10064,nx10064,nx10066,nx10066,nx10066,nx10068,nx10068,
               nx10068,nx10070,nx10070,nx10070,nx10072,nx10072,nx10072,nx10074,
               nx10074,nx10074,nx10076,nx10076,nx10076,nx10078,nx10078,nx10078,
               nx10080,nx10080,nx10080,nx10082,nx10082,nx10082,nx10084,nx10084,
               nx10084,nx10086,nx10086,nx10086,nx10088,nx10088,nx10088,nx10090,
               nx10090,nx10090,nx10092,nx10092,nx10092,nx10094,nx10094,nx10094,
               nx10096,nx10096,nx10096,nx10098,nx10098,nx10098,nx10100,nx10100,
               nx10100,nx10102,nx10102,nx10102,nx10104,nx10104,nx10104,nx10106,
               nx10106,nx10106,nx10108,nx10108,nx10108,nx10110,nx10110,nx10110,
               nx10112,nx10112,nx10112,nx10114,nx10114,nx10114,nx10116,nx10116,
               nx10116,nx10118,nx10118,nx10118,nx10120,nx10120,nx10120,nx10122,
               nx10122,nx10122,nx10124,nx10124,nx10124,nx10126,nx10126,nx10126,
               nx10128,nx10128,nx10128,nx10130,nx10130,nx10130,nx10132,nx10132,
               nx10132,nx10134,nx10134,nx10134,nx10136,nx10136,nx10136,nx10138,
               nx10138,nx10138,nx10140,nx10140,nx10140,nx10142,nx10142,nx10142,
               nx10144,nx10144,nx10144,nx10146,nx10146,nx10146,nx10148,nx10148,
               nx10148,nx10150,nx10150,nx10150,nx10152,nx10152,nx10152,nx10154,
               nx10154,nx10154,nx10156,nx10156,nx10156,nx10158,nx10158,nx10158,
               nx10160,nx10160,nx10160,nx10162,nx10162,nx10162,nx10164,nx10164,
               nx10164,nx10166,nx10166,nx10166,nx10168,nx10168,nx10168,nx10170,
               nx10170,nx10170,nx10172,nx10172,nx10172,nx10174,nx10174,nx10174,
               nx10176,nx10176,nx10176,nx10178,nx10178,nx10178,nx10180,nx10180,
               nx10180,nx10182,nx10182,nx10182,nx10184,nx10184,nx10184,nx10186,
               nx10186,nx10186,nx10188,nx10188,nx10188,nx10190,nx10190,nx10190,
               nx10192,nx10192,nx10192,nx10194,nx10194,nx10194,nx10196,nx10196,
               nx10196,nx10198,nx10198,nx10198,nx10200,nx10200,nx10200,nx10202,
               nx10202,nx10202,nx10204,nx10204,nx10204,nx10206,nx10206,nx10206,
               nx10208,nx10208,nx10208,nx10210,nx10210,nx10210,nx10212,nx10212,
               nx10212,nx10214,nx10214,nx10214,nx10216,nx10216,nx10216,nx10218,
               nx10218,nx10218,nx10220,nx10220,nx10220,nx10222,nx10222,nx10222,
               nx10224,nx10224,nx10224,nx10226,nx10226,nx10226,nx10228,nx10228,
               nx10228,nx10230,nx10230,nx10230,nx10232,nx10232,nx10232,nx10234,
               nx10234,nx10234,nx10236,nx10236,nx10236,nx10238,nx10238,nx10238,
               nx10240,nx10240,nx10240,nx10242,nx10242,nx10242,nx10244,nx10244,
               nx10244,nx10246,nx10246,nx10246,nx10248,nx10248,nx10248,nx10250,
               nx10250,nx10250,nx10252,nx10252,nx10252,nx10254,nx10254,nx10254,
               nx10256,nx10256,nx10256,nx10258,nx10258,nx10258,nx10260,nx10260,
               nx10260,nx10262,nx10262,nx10262,nx10264,nx10264,nx10264,nx10266,
               nx10266,nx10266,nx10268,nx10268,nx10268,nx10270,nx10270,nx10270,
               nx10272,nx10272,nx10272,nx10274,nx10274,nx10274,nx10276,nx10276,
               nx10276,nx10278,nx10278,nx10278,nx10280,nx10280,nx10280,nx10282,
               nx10282,nx10282,nx10284,nx10284,nx10284,nx10286,nx10286,nx10286,
               nx10288,nx10288,nx10288,nx10290,nx10290,nx10290,nx10292,nx10294,
               nx10296,nx10296,nx10298,nx10300,nx10300,nx10302,nx10304,nx10306})
               , .FilterAddress ({nx9976,nx9980,nx9984,nx9988,nx9992,nx9996,
               nx10000,nx10004,nx10008,nx10012,nx10016,nx10020,nx10024}), .msbNoOfFilters (
               nx10500), .CLK (nx10422), .RST (rst), .QImgStat (Q), .ACKF (
               nx10308), .IndicatorFilter ({IndicatorF_0}), .DMAAddress ({
               AddressF_12,AddressF_11,AddressF_10,AddressF_9,AddressF_8,
               AddressF_7,AddressF_6,AddressF_5,AddressF_4,AddressF_3,AddressF_2
               ,AddressF_1,AddressF_0}), .UpdatedAddress ({FilterAddressIN_12,
               FilterAddressIN_11,FilterAddressIN_10,FilterAddressIN_9,
               FilterAddressIN_8,FilterAddressIN_7,FilterAddressIN_6,
               FilterAddressIN_5,FilterAddressIN_4,FilterAddressIN_3,
               FilterAddressIN_2,FilterAddressIN_1,FilterAddressIN_0}), .outFilter0 (
               {Filter1_399,Filter1_398,Filter1_397,Filter1_396,Filter1_395,
               Filter1_394,Filter1_393,Filter1_392,Filter1_391,Filter1_390,
               Filter1_389,Filter1_388,Filter1_387,Filter1_386,Filter1_385,
               Filter1_384,Filter1_383,Filter1_382,Filter1_381,Filter1_380,
               Filter1_379,Filter1_378,Filter1_377,Filter1_376,Filter1_375,
               Filter1_374,Filter1_373,Filter1_372,Filter1_371,Filter1_370,
               Filter1_369,Filter1_368,Filter1_367,Filter1_366,Filter1_365,
               Filter1_364,Filter1_363,Filter1_362,Filter1_361,Filter1_360,
               Filter1_359,Filter1_358,Filter1_357,Filter1_356,Filter1_355,
               Filter1_354,Filter1_353,Filter1_352,Filter1_351,Filter1_350,
               Filter1_349,Filter1_348,Filter1_347,Filter1_346,Filter1_345,
               Filter1_344,Filter1_343,Filter1_342,Filter1_341,Filter1_340,
               Filter1_339,Filter1_338,Filter1_337,Filter1_336,Filter1_335,
               Filter1_334,Filter1_333,Filter1_332,Filter1_331,Filter1_330,
               Filter1_329,Filter1_328,Filter1_327,Filter1_326,Filter1_325,
               Filter1_324,Filter1_323,Filter1_322,Filter1_321,Filter1_320,
               Filter1_319,Filter1_318,Filter1_317,Filter1_316,Filter1_315,
               Filter1_314,Filter1_313,Filter1_312,Filter1_311,Filter1_310,
               Filter1_309,Filter1_308,Filter1_307,Filter1_306,Filter1_305,
               Filter1_304,Filter1_303,Filter1_302,Filter1_301,Filter1_300,
               Filter1_299,Filter1_298,Filter1_297,Filter1_296,Filter1_295,
               Filter1_294,Filter1_293,Filter1_292,Filter1_291,Filter1_290,
               Filter1_289,Filter1_288,Filter1_287,Filter1_286,Filter1_285,
               Filter1_284,Filter1_283,Filter1_282,Filter1_281,Filter1_280,
               Filter1_279,Filter1_278,Filter1_277,Filter1_276,Filter1_275,
               Filter1_274,Filter1_273,Filter1_272,Filter1_271,Filter1_270,
               Filter1_269,Filter1_268,Filter1_267,Filter1_266,Filter1_265,
               Filter1_264,Filter1_263,Filter1_262,Filter1_261,Filter1_260,
               Filter1_259,Filter1_258,Filter1_257,Filter1_256,Filter1_255,
               Filter1_254,Filter1_253,Filter1_252,Filter1_251,Filter1_250,
               Filter1_249,Filter1_248,Filter1_247,Filter1_246,Filter1_245,
               Filter1_244,Filter1_243,Filter1_242,Filter1_241,Filter1_240,
               Filter1_239,Filter1_238,Filter1_237,Filter1_236,Filter1_235,
               Filter1_234,Filter1_233,Filter1_232,Filter1_231,Filter1_230,
               Filter1_229,Filter1_228,Filter1_227,Filter1_226,Filter1_225,
               Filter1_224,Filter1_223,Filter1_222,Filter1_221,Filter1_220,
               Filter1_219,Filter1_218,Filter1_217,Filter1_216,Filter1_215,
               Filter1_214,Filter1_213,Filter1_212,Filter1_211,Filter1_210,
               Filter1_209,Filter1_208,Filter1_207,Filter1_206,Filter1_205,
               Filter1_204,Filter1_203,Filter1_202,Filter1_201,Filter1_200,
               Filter1_199,Filter1_198,Filter1_197,Filter1_196,Filter1_195,
               Filter1_194,Filter1_193,Filter1_192,Filter1_191,Filter1_190,
               Filter1_189,Filter1_188,Filter1_187,Filter1_186,Filter1_185,
               Filter1_184,Filter1_183,Filter1_182,Filter1_181,Filter1_180,
               Filter1_179,Filter1_178,Filter1_177,Filter1_176,Filter1_175,
               Filter1_174,Filter1_173,Filter1_172,Filter1_171,Filter1_170,
               Filter1_169,Filter1_168,Filter1_167,Filter1_166,Filter1_165,
               Filter1_164,Filter1_163,Filter1_162,Filter1_161,Filter1_160,
               Filter1_159,Filter1_158,Filter1_157,Filter1_156,Filter1_155,
               Filter1_154,Filter1_153,Filter1_152,Filter1_151,Filter1_150,
               Filter1_149,Filter1_148,Filter1_147,Filter1_146,Filter1_145,
               Filter1_144,Filter1_143,Filter1_142,Filter1_141,Filter1_140,
               Filter1_139,Filter1_138,Filter1_137,Filter1_136,Filter1_135,
               Filter1_134,Filter1_133,Filter1_132,Filter1_131,Filter1_130,
               Filter1_129,Filter1_128,Filter1_127,Filter1_126,Filter1_125,
               Filter1_124,Filter1_123,Filter1_122,Filter1_121,Filter1_120,
               Filter1_119,Filter1_118,Filter1_117,Filter1_116,Filter1_115,
               Filter1_114,Filter1_113,Filter1_112,Filter1_111,Filter1_110,
               Filter1_109,Filter1_108,Filter1_107,Filter1_106,Filter1_105,
               Filter1_104,Filter1_103,Filter1_102,Filter1_101,Filter1_100,
               Filter1_99,Filter1_98,Filter1_97,Filter1_96,Filter1_95,Filter1_94
               ,Filter1_93,Filter1_92,Filter1_91,Filter1_90,Filter1_89,
               Filter1_88,Filter1_87,Filter1_86,Filter1_85,Filter1_84,Filter1_83
               ,Filter1_82,Filter1_81,Filter1_80,Filter1_79,Filter1_78,
               Filter1_77,Filter1_76,Filter1_75,Filter1_74,Filter1_73,Filter1_72
               ,Filter1_71,Filter1_70,Filter1_69,Filter1_68,Filter1_67,
               Filter1_66,Filter1_65,Filter1_64,Filter1_63,Filter1_62,Filter1_61
               ,Filter1_60,Filter1_59,Filter1_58,Filter1_57,Filter1_56,
               Filter1_55,Filter1_54,Filter1_53,Filter1_52,Filter1_51,Filter1_50
               ,Filter1_49,Filter1_48,Filter1_47,Filter1_46,Filter1_45,
               Filter1_44,Filter1_43,Filter1_42,Filter1_41,Filter1_40,Filter1_39
               ,Filter1_38,Filter1_37,Filter1_36,Filter1_35,Filter1_34,
               Filter1_33,Filter1_32,Filter1_31,Filter1_30,Filter1_29,Filter1_28
               ,Filter1_27,Filter1_26,Filter1_25,Filter1_24,Filter1_23,
               Filter1_22,Filter1_21,Filter1_20,Filter1_19,Filter1_18,Filter1_17
               ,Filter1_16,Filter1_15,Filter1_14,Filter1_13,Filter1_12,
               Filter1_11,Filter1_10,Filter1_9,Filter1_8,Filter1_7,Filter1_6,
               Filter1_5,Filter1_4,Filter1_3,Filter1_2,Filter1_1,Filter1_0}), .outFilter1 (
               {Filter2_399,Filter2_398,Filter2_397,Filter2_396,Filter2_395,
               Filter2_394,Filter2_393,Filter2_392,Filter2_391,Filter2_390,
               Filter2_389,Filter2_388,Filter2_387,Filter2_386,Filter2_385,
               Filter2_384,Filter2_383,Filter2_382,Filter2_381,Filter2_380,
               Filter2_379,Filter2_378,Filter2_377,Filter2_376,Filter2_375,
               Filter2_374,Filter2_373,Filter2_372,Filter2_371,Filter2_370,
               Filter2_369,Filter2_368,Filter2_367,Filter2_366,Filter2_365,
               Filter2_364,Filter2_363,Filter2_362,Filter2_361,Filter2_360,
               Filter2_359,Filter2_358,Filter2_357,Filter2_356,Filter2_355,
               Filter2_354,Filter2_353,Filter2_352,Filter2_351,Filter2_350,
               Filter2_349,Filter2_348,Filter2_347,Filter2_346,Filter2_345,
               Filter2_344,Filter2_343,Filter2_342,Filter2_341,Filter2_340,
               Filter2_339,Filter2_338,Filter2_337,Filter2_336,Filter2_335,
               Filter2_334,Filter2_333,Filter2_332,Filter2_331,Filter2_330,
               Filter2_329,Filter2_328,Filter2_327,Filter2_326,Filter2_325,
               Filter2_324,Filter2_323,Filter2_322,Filter2_321,Filter2_320,
               Filter2_319,Filter2_318,Filter2_317,Filter2_316,Filter2_315,
               Filter2_314,Filter2_313,Filter2_312,Filter2_311,Filter2_310,
               Filter2_309,Filter2_308,Filter2_307,Filter2_306,Filter2_305,
               Filter2_304,Filter2_303,Filter2_302,Filter2_301,Filter2_300,
               Filter2_299,Filter2_298,Filter2_297,Filter2_296,Filter2_295,
               Filter2_294,Filter2_293,Filter2_292,Filter2_291,Filter2_290,
               Filter2_289,Filter2_288,Filter2_287,Filter2_286,Filter2_285,
               Filter2_284,Filter2_283,Filter2_282,Filter2_281,Filter2_280,
               Filter2_279,Filter2_278,Filter2_277,Filter2_276,Filter2_275,
               Filter2_274,Filter2_273,Filter2_272,Filter2_271,Filter2_270,
               Filter2_269,Filter2_268,Filter2_267,Filter2_266,Filter2_265,
               Filter2_264,Filter2_263,Filter2_262,Filter2_261,Filter2_260,
               Filter2_259,Filter2_258,Filter2_257,Filter2_256,Filter2_255,
               Filter2_254,Filter2_253,Filter2_252,Filter2_251,Filter2_250,
               Filter2_249,Filter2_248,Filter2_247,Filter2_246,Filter2_245,
               Filter2_244,Filter2_243,Filter2_242,Filter2_241,Filter2_240,
               Filter2_239,Filter2_238,Filter2_237,Filter2_236,Filter2_235,
               Filter2_234,Filter2_233,Filter2_232,Filter2_231,Filter2_230,
               Filter2_229,Filter2_228,Filter2_227,Filter2_226,Filter2_225,
               Filter2_224,Filter2_223,Filter2_222,Filter2_221,Filter2_220,
               Filter2_219,Filter2_218,Filter2_217,Filter2_216,Filter2_215,
               Filter2_214,Filter2_213,Filter2_212,Filter2_211,Filter2_210,
               Filter2_209,Filter2_208,Filter2_207,Filter2_206,Filter2_205,
               Filter2_204,Filter2_203,Filter2_202,Filter2_201,Filter2_200,
               Filter2_199,Filter2_198,Filter2_197,Filter2_196,Filter2_195,
               Filter2_194,Filter2_193,Filter2_192,Filter2_191,Filter2_190,
               Filter2_189,Filter2_188,Filter2_187,Filter2_186,Filter2_185,
               Filter2_184,Filter2_183,Filter2_182,Filter2_181,Filter2_180,
               Filter2_179,Filter2_178,Filter2_177,Filter2_176,Filter2_175,
               Filter2_174,Filter2_173,Filter2_172,Filter2_171,Filter2_170,
               Filter2_169,Filter2_168,Filter2_167,Filter2_166,Filter2_165,
               Filter2_164,Filter2_163,Filter2_162,Filter2_161,Filter2_160,
               Filter2_159,Filter2_158,Filter2_157,Filter2_156,Filter2_155,
               Filter2_154,Filter2_153,Filter2_152,Filter2_151,Filter2_150,
               Filter2_149,Filter2_148,Filter2_147,Filter2_146,Filter2_145,
               Filter2_144,Filter2_143,Filter2_142,Filter2_141,Filter2_140,
               Filter2_139,Filter2_138,Filter2_137,Filter2_136,Filter2_135,
               Filter2_134,Filter2_133,Filter2_132,Filter2_131,Filter2_130,
               Filter2_129,Filter2_128,Filter2_127,Filter2_126,Filter2_125,
               Filter2_124,Filter2_123,Filter2_122,Filter2_121,Filter2_120,
               Filter2_119,Filter2_118,Filter2_117,Filter2_116,Filter2_115,
               Filter2_114,Filter2_113,Filter2_112,Filter2_111,Filter2_110,
               Filter2_109,Filter2_108,Filter2_107,Filter2_106,Filter2_105,
               Filter2_104,Filter2_103,Filter2_102,Filter2_101,Filter2_100,
               Filter2_99,Filter2_98,Filter2_97,Filter2_96,Filter2_95,Filter2_94
               ,Filter2_93,Filter2_92,Filter2_91,Filter2_90,Filter2_89,
               Filter2_88,Filter2_87,Filter2_86,Filter2_85,Filter2_84,Filter2_83
               ,Filter2_82,Filter2_81,Filter2_80,Filter2_79,Filter2_78,
               Filter2_77,Filter2_76,Filter2_75,Filter2_74,Filter2_73,Filter2_72
               ,Filter2_71,Filter2_70,Filter2_69,Filter2_68,Filter2_67,
               Filter2_66,Filter2_65,Filter2_64,Filter2_63,Filter2_62,Filter2_61
               ,Filter2_60,Filter2_59,Filter2_58,Filter2_57,Filter2_56,
               Filter2_55,Filter2_54,Filter2_53,Filter2_52,Filter2_51,Filter2_50
               ,Filter2_49,Filter2_48,Filter2_47,Filter2_46,Filter2_45,
               Filter2_44,Filter2_43,Filter2_42,Filter2_41,Filter2_40,Filter2_39
               ,Filter2_38,Filter2_37,Filter2_36,Filter2_35,Filter2_34,
               Filter2_33,Filter2_32,Filter2_31,Filter2_30,Filter2_29,Filter2_28
               ,Filter2_27,Filter2_26,Filter2_25,Filter2_24,Filter2_23,
               Filter2_22,Filter2_21,Filter2_20,Filter2_19,Filter2_18,Filter2_17
               ,Filter2_16,Filter2_15,Filter2_14,Filter2_13,Filter2_12,
               Filter2_11,Filter2_10,Filter2_9,Filter2_8,Filter2_7,Filter2_6,
               Filter2_5,Filter2_4,Filter2_3,Filter2_2,Filter2_1,Filter2_0}), .donttrust (
               DontRstIndicator), .LastFilterIND (lastFilter), .LastHeightOut (
               \$dummy [431]), .lastDepthOut (lastDepthOut)) ;
    ReadImage RImg (.WI (WriteI), .current_state ({zero_11,zero_11,nx9954,
              current_state_11,current_state_10,zero_11,current_state_8,nx9962,
              current_state_6,current_state_5,nx9966,current_state_3,
              current_state_2,zero_11,zero_11}), .CLK (nx10418), .RST (rst), .ACK (
              nx10026), .ImgAddress ({ImgAddRegOut_12,ImgAddRegOut_11,
              ImgAddRegOut_10,ImgAddRegOut_9,ImgAddRegOut_8,ImgAddRegOut_7,
              ImgAddRegOut_6,ImgAddRegOut_5,ImgAddRegOut_4,ImgAddRegOut_3,
              ImgAddRegOut_2,ImgAddRegOut_1,ImgAddRegOut_0}), .ImgWidth ({
              ImgWidthOut_15,ImgWidthOut_14,ImgWidthOut_13,ImgWidthOut_12,
              ImgWidthOut_11,ImgWidthOut_10,ImgWidthOut_9,ImgWidthOut_8,
              ImgWidthOut_7,ImgWidthOut_6,ImgWidthOut_5,ImgWidthOut_4,
              ImgWidthOut_3,ImgWidthOut_2,ImgWidthOut_1,ImgWidthOut_0}), .DATA (
              {DataIOut_447,DataIOut_446,DataIOut_445,DataIOut_444,DataIOut_443,
              DataIOut_442,DataIOut_441,DataIOut_440,DataIOut_439,DataIOut_438,
              DataIOut_437,DataIOut_436,DataIOut_435,DataIOut_434,DataIOut_433,
              DataIOut_432,DataIOut_431,DataIOut_430,DataIOut_429,DataIOut_428,
              DataIOut_427,DataIOut_426,DataIOut_425,DataIOut_424,DataIOut_423,
              DataIOut_422,DataIOut_421,DataIOut_420,DataIOut_419,DataIOut_418,
              DataIOut_417,DataIOut_416,DataIOut_415,DataIOut_414,DataIOut_413,
              DataIOut_412,DataIOut_411,DataIOut_410,DataIOut_409,DataIOut_408,
              DataIOut_407,DataIOut_406,DataIOut_405,DataIOut_404,DataIOut_403,
              DataIOut_402,DataIOut_401,DataIOut_400,DataIOut_399,DataIOut_398,
              DataIOut_397,DataIOut_396,DataIOut_395,DataIOut_394,DataIOut_393,
              DataIOut_392,DataIOut_391,DataIOut_390,DataIOut_389,DataIOut_388,
              DataIOut_387,DataIOut_386,DataIOut_385,DataIOut_384,DataIOut_383,
              DataIOut_382,DataIOut_381,DataIOut_380,DataIOut_379,DataIOut_378,
              DataIOut_377,DataIOut_376,DataIOut_375,DataIOut_374,DataIOut_373,
              DataIOut_372,DataIOut_371,DataIOut_370,DataIOut_369,DataIOut_368,
              DataIOut_367,DataIOut_366,DataIOut_365,DataIOut_364,DataIOut_363,
              DataIOut_362,DataIOut_361,DataIOut_360,DataIOut_359,DataIOut_358,
              DataIOut_357,DataIOut_356,DataIOut_355,DataIOut_354,DataIOut_353,
              DataIOut_352,DataIOut_351,DataIOut_350,DataIOut_349,DataIOut_348,
              DataIOut_347,DataIOut_346,DataIOut_345,DataIOut_344,DataIOut_343,
              DataIOut_342,DataIOut_341,DataIOut_340,DataIOut_339,DataIOut_338,
              DataIOut_337,DataIOut_336,DataIOut_335,DataIOut_334,DataIOut_333,
              DataIOut_332,DataIOut_331,DataIOut_330,DataIOut_329,DataIOut_328,
              DataIOut_327,DataIOut_326,DataIOut_325,DataIOut_324,DataIOut_323,
              DataIOut_322,DataIOut_321,DataIOut_320,DataIOut_319,DataIOut_318,
              DataIOut_317,DataIOut_316,DataIOut_315,DataIOut_314,DataIOut_313,
              DataIOut_312,DataIOut_311,DataIOut_310,DataIOut_309,DataIOut_308,
              DataIOut_307,DataIOut_306,DataIOut_305,DataIOut_304,DataIOut_303,
              DataIOut_302,DataIOut_301,DataIOut_300,DataIOut_299,DataIOut_298,
              DataIOut_297,DataIOut_296,DataIOut_295,DataIOut_294,DataIOut_293,
              DataIOut_292,DataIOut_291,DataIOut_290,DataIOut_289,DataIOut_288,
              DataIOut_287,DataIOut_286,DataIOut_285,DataIOut_284,DataIOut_283,
              DataIOut_282,DataIOut_281,DataIOut_280,DataIOut_279,DataIOut_278,
              DataIOut_277,DataIOut_276,DataIOut_275,DataIOut_274,DataIOut_273,
              DataIOut_272,DataIOut_271,DataIOut_270,DataIOut_269,DataIOut_268,
              DataIOut_267,DataIOut_266,DataIOut_265,DataIOut_264,DataIOut_263,
              DataIOut_262,DataIOut_261,DataIOut_260,DataIOut_259,DataIOut_258,
              DataIOut_257,DataIOut_256,DataIOut_255,DataIOut_254,DataIOut_253,
              DataIOut_252,DataIOut_251,DataIOut_250,DataIOut_249,DataIOut_248,
              DataIOut_247,DataIOut_246,DataIOut_245,DataIOut_244,DataIOut_243,
              DataIOut_242,DataIOut_241,DataIOut_240,DataIOut_239,DataIOut_238,
              DataIOut_237,DataIOut_236,DataIOut_235,DataIOut_234,DataIOut_233,
              DataIOut_232,DataIOut_231,DataIOut_230,DataIOut_229,DataIOut_228,
              DataIOut_227,DataIOut_226,DataIOut_225,DataIOut_224,DataIOut_223,
              DataIOut_222,DataIOut_221,DataIOut_220,DataIOut_219,DataIOut_218,
              DataIOut_217,DataIOut_216,DataIOut_215,DataIOut_214,DataIOut_213,
              DataIOut_212,DataIOut_211,DataIOut_210,DataIOut_209,DataIOut_208,
              DataIOut_207,DataIOut_206,DataIOut_205,DataIOut_204,DataIOut_203,
              DataIOut_202,DataIOut_201,DataIOut_200,DataIOut_199,DataIOut_198,
              DataIOut_197,DataIOut_196,DataIOut_195,DataIOut_194,DataIOut_193,
              DataIOut_192,DataIOut_191,DataIOut_190,DataIOut_189,DataIOut_188,
              DataIOut_187,DataIOut_186,DataIOut_185,DataIOut_184,DataIOut_183,
              DataIOut_182,DataIOut_181,DataIOut_180,DataIOut_179,DataIOut_178,
              DataIOut_177,DataIOut_176,DataIOut_175,DataIOut_174,DataIOut_173,
              DataIOut_172,DataIOut_171,DataIOut_170,DataIOut_169,DataIOut_168,
              DataIOut_167,DataIOut_166,DataIOut_165,DataIOut_164,DataIOut_163,
              DataIOut_162,DataIOut_161,DataIOut_160,DataIOut_159,DataIOut_158,
              DataIOut_157,DataIOut_156,DataIOut_155,DataIOut_154,DataIOut_153,
              DataIOut_152,DataIOut_151,DataIOut_150,DataIOut_149,DataIOut_148,
              DataIOut_147,DataIOut_146,DataIOut_145,DataIOut_144,DataIOut_143,
              DataIOut_142,DataIOut_141,DataIOut_140,DataIOut_139,DataIOut_138,
              DataIOut_137,DataIOut_136,DataIOut_135,DataIOut_134,DataIOut_133,
              DataIOut_132,DataIOut_131,DataIOut_130,DataIOut_129,DataIOut_128,
              DataIOut_127,DataIOut_126,DataIOut_125,DataIOut_124,DataIOut_123,
              DataIOut_122,DataIOut_121,DataIOut_120,DataIOut_119,DataIOut_118,
              DataIOut_117,DataIOut_116,DataIOut_115,DataIOut_114,DataIOut_113,
              DataIOut_112,DataIOut_111,DataIOut_110,DataIOut_109,DataIOut_108,
              DataIOut_107,DataIOut_106,DataIOut_105,DataIOut_104,DataIOut_103,
              DataIOut_102,DataIOut_101,DataIOut_100,DataIOut_99,DataIOut_98,
              DataIOut_97,DataIOut_96,DataIOut_95,DataIOut_94,DataIOut_93,
              DataIOut_92,DataIOut_91,DataIOut_90,DataIOut_89,DataIOut_88,
              DataIOut_87,DataIOut_86,DataIOut_85,DataIOut_84,DataIOut_83,
              DataIOut_82,DataIOut_81,DataIOut_80,DataIOut_79,DataIOut_78,
              DataIOut_77,DataIOut_76,DataIOut_75,DataIOut_74,DataIOut_73,
              DataIOut_72,DataIOut_71,DataIOut_70,DataIOut_69,DataIOut_68,
              DataIOut_67,DataIOut_66,DataIOut_65,DataIOut_64,DataIOut_63,
              DataIOut_62,DataIOut_61,DataIOut_60,DataIOut_59,DataIOut_58,
              DataIOut_57,DataIOut_56,DataIOut_55,DataIOut_54,DataIOut_53,
              DataIOut_52,DataIOut_51,DataIOut_50,DataIOut_49,DataIOut_48,
              DataIOut_47,DataIOut_46,DataIOut_45,DataIOut_44,DataIOut_43,
              DataIOut_42,DataIOut_41,DataIOut_40,DataIOut_39,DataIOut_38,
              DataIOut_37,DataIOut_36,DataIOut_35,DataIOut_34,DataIOut_33,
              DataIOut_32,DataIOut_31,DataIOut_30,DataIOut_29,DataIOut_28,
              DataIOut_27,DataIOut_26,DataIOut_25,DataIOut_24,DataIOut_23,
              DataIOut_22,DataIOut_21,DataIOut_20,DataIOut_19,DataIOut_18,
              DataIOut_17,DataIOut_16,nx10312,nx10316,nx10320,nx10324,nx10328,
              nx10332,nx10336,nx10340,nx10344,nx10348,nx10352,nx10356,nx10360,
              nx10364,nx10368,nx10372}), .OutputImg0 ({\$dummy [432],
              \$dummy [433],\$dummy [434],\$dummy [435],\$dummy [436],
              \$dummy [437],\$dummy [438],\$dummy [439],\$dummy [440],
              \$dummy [441],\$dummy [442],\$dummy [443],\$dummy [444],
              \$dummy [445],\$dummy [446],\$dummy [447],\$dummy [448],
              \$dummy [449],\$dummy [450],\$dummy [451],\$dummy [452],
              \$dummy [453],\$dummy [454],\$dummy [455],\$dummy [456],
              \$dummy [457],\$dummy [458],\$dummy [459],\$dummy [460],
              \$dummy [461],\$dummy [462],\$dummy [463],\$dummy [464],
              \$dummy [465],\$dummy [466],\$dummy [467],\$dummy [468],
              \$dummy [469],\$dummy [470],\$dummy [471],\$dummy [472],
              \$dummy [473],\$dummy [474],\$dummy [475],\$dummy [476],
              \$dummy [477],\$dummy [478],\$dummy [479],\$dummy [480],
              \$dummy [481],\$dummy [482],\$dummy [483],\$dummy [484],
              \$dummy [485],\$dummy [486],\$dummy [487],\$dummy [488],
              \$dummy [489],\$dummy [490],\$dummy [491],\$dummy [492],
              \$dummy [493],\$dummy [494],\$dummy [495],\$dummy [496],
              \$dummy [497],\$dummy [498],\$dummy [499],\$dummy [500],
              \$dummy [501],\$dummy [502],\$dummy [503],\$dummy [504],
              \$dummy [505],\$dummy [506],\$dummy [507],\$dummy [508],
              \$dummy [509],\$dummy [510],\$dummy [511],\$dummy [512],
              \$dummy [513],\$dummy [514],\$dummy [515],\$dummy [516],
              \$dummy [517],\$dummy [518],\$dummy [519],\$dummy [520],
              \$dummy [521],\$dummy [522],\$dummy [523],\$dummy [524],
              \$dummy [525],\$dummy [526],\$dummy [527],\$dummy [528],
              \$dummy [529],\$dummy [530],\$dummy [531],\$dummy [532],
              \$dummy [533],\$dummy [534],\$dummy [535],\$dummy [536],
              \$dummy [537],\$dummy [538],\$dummy [539],\$dummy [540],
              \$dummy [541],\$dummy [542],\$dummy [543],\$dummy [544],
              \$dummy [545],\$dummy [546],\$dummy [547],\$dummy [548],
              \$dummy [549],\$dummy [550],\$dummy [551],\$dummy [552],
              \$dummy [553],\$dummy [554],\$dummy [555],\$dummy [556],
              \$dummy [557],\$dummy [558],\$dummy [559],\$dummy [560],
              \$dummy [561],\$dummy [562],\$dummy [563],\$dummy [564],
              \$dummy [565],\$dummy [566],\$dummy [567],\$dummy [568],
              \$dummy [569],\$dummy [570],\$dummy [571],\$dummy [572],
              \$dummy [573],\$dummy [574],\$dummy [575],\$dummy [576],
              \$dummy [577],\$dummy [578],\$dummy [579],\$dummy [580],
              \$dummy [581],\$dummy [582],\$dummy [583],\$dummy [584],
              \$dummy [585],\$dummy [586],\$dummy [587],\$dummy [588],
              \$dummy [589],\$dummy [590],\$dummy [591],\$dummy [592],
              \$dummy [593],\$dummy [594],\$dummy [595],\$dummy [596],
              \$dummy [597],\$dummy [598],\$dummy [599],\$dummy [600],
              \$dummy [601],\$dummy [602],\$dummy [603],\$dummy [604],
              \$dummy [605],\$dummy [606],\$dummy [607],\$dummy [608],
              \$dummy [609],\$dummy [610],\$dummy [611],\$dummy [612],
              \$dummy [613],\$dummy [614],\$dummy [615],\$dummy [616],
              \$dummy [617],\$dummy [618],\$dummy [619],\$dummy [620],
              \$dummy [621],\$dummy [622],\$dummy [623],\$dummy [624],
              \$dummy [625],\$dummy [626],\$dummy [627],\$dummy [628],
              \$dummy [629],\$dummy [630],\$dummy [631],\$dummy [632],
              \$dummy [633],\$dummy [634],\$dummy [635],\$dummy [636],
              \$dummy [637],\$dummy [638],\$dummy [639],\$dummy [640],
              \$dummy [641],\$dummy [642],\$dummy [643],\$dummy [644],
              \$dummy [645],\$dummy [646],\$dummy [647],\$dummy [648],
              \$dummy [649],\$dummy [650],\$dummy [651],\$dummy [652],
              \$dummy [653],\$dummy [654],\$dummy [655],\$dummy [656],
              \$dummy [657],\$dummy [658],\$dummy [659],\$dummy [660],
              \$dummy [661],\$dummy [662],\$dummy [663],\$dummy [664],
              \$dummy [665],\$dummy [666],\$dummy [667],\$dummy [668],
              \$dummy [669],\$dummy [670],\$dummy [671],\$dummy [672],
              \$dummy [673],\$dummy [674],\$dummy [675],\$dummy [676],
              \$dummy [677],\$dummy [678],\$dummy [679],\$dummy [680],
              \$dummy [681],\$dummy [682],\$dummy [683],\$dummy [684],
              \$dummy [685],\$dummy [686],\$dummy [687],\$dummy [688],
              \$dummy [689],\$dummy [690],\$dummy [691],\$dummy [692],
              \$dummy [693],\$dummy [694],\$dummy [695],\$dummy [696],
              \$dummy [697],\$dummy [698],\$dummy [699],\$dummy [700],
              \$dummy [701],\$dummy [702],\$dummy [703],\$dummy [704],
              \$dummy [705],\$dummy [706],\$dummy [707],\$dummy [708],
              \$dummy [709],\$dummy [710],\$dummy [711],\$dummy [712],
              \$dummy [713],\$dummy [714],\$dummy [715],\$dummy [716],
              \$dummy [717],\$dummy [718],\$dummy [719],\$dummy [720],
              \$dummy [721],\$dummy [722],\$dummy [723],\$dummy [724],
              \$dummy [725],\$dummy [726],\$dummy [727],\$dummy [728],
              \$dummy [729],\$dummy [730],\$dummy [731],\$dummy [732],
              \$dummy [733],\$dummy [734],\$dummy [735],\$dummy [736],
              \$dummy [737],\$dummy [738],\$dummy [739],\$dummy [740],
              \$dummy [741],\$dummy [742],\$dummy [743],\$dummy [744],
              \$dummy [745],\$dummy [746],\$dummy [747],\$dummy [748],
              \$dummy [749],\$dummy [750],\$dummy [751],\$dummy [752],
              \$dummy [753],\$dummy [754],\$dummy [755],\$dummy [756],
              \$dummy [757],\$dummy [758],\$dummy [759],\$dummy [760],
              \$dummy [761],\$dummy [762],\$dummy [763],\$dummy [764],
              \$dummy [765],\$dummy [766],\$dummy [767],\$dummy [768],
              \$dummy [769],\$dummy [770],\$dummy [771],\$dummy [772],
              \$dummy [773],\$dummy [774],\$dummy [775],\$dummy [776],
              \$dummy [777],\$dummy [778],\$dummy [779],\$dummy [780],
              \$dummy [781],\$dummy [782],\$dummy [783],\$dummy [784],
              \$dummy [785],\$dummy [786],\$dummy [787],\$dummy [788],
              \$dummy [789],\$dummy [790],\$dummy [791],\$dummy [792],
              \$dummy [793],\$dummy [794],\$dummy [795],\$dummy [796],
              \$dummy [797],\$dummy [798],\$dummy [799],OutputImg0_79,
              OutputImg0_78,OutputImg0_77,OutputImg0_76,OutputImg0_75,
              OutputImg0_74,OutputImg0_73,OutputImg0_72,OutputImg0_71,
              OutputImg0_70,OutputImg0_69,OutputImg0_68,OutputImg0_67,
              OutputImg0_66,OutputImg0_65,OutputImg0_64,OutputImg0_63,
              OutputImg0_62,OutputImg0_61,OutputImg0_60,OutputImg0_59,
              OutputImg0_58,OutputImg0_57,OutputImg0_56,OutputImg0_55,
              OutputImg0_54,OutputImg0_53,OutputImg0_52,OutputImg0_51,
              OutputImg0_50,OutputImg0_49,OutputImg0_48,OutputImg0_47,
              OutputImg0_46,OutputImg0_45,OutputImg0_44,OutputImg0_43,
              OutputImg0_42,OutputImg0_41,OutputImg0_40,OutputImg0_39,
              OutputImg0_38,OutputImg0_37,OutputImg0_36,OutputImg0_35,
              OutputImg0_34,OutputImg0_33,OutputImg0_32,OutputImg0_31,
              OutputImg0_30,OutputImg0_29,OutputImg0_28,OutputImg0_27,
              OutputImg0_26,OutputImg0_25,OutputImg0_24,OutputImg0_23,
              OutputImg0_22,OutputImg0_21,OutputImg0_20,OutputImg0_19,
              OutputImg0_18,OutputImg0_17,OutputImg0_16,OutputImg0_15,
              OutputImg0_14,OutputImg0_13,OutputImg0_12,OutputImg0_11,
              OutputImg0_10,OutputImg0_9,OutputImg0_8,OutputImg0_7,OutputImg0_6,
              OutputImg0_5,OutputImg0_4,OutputImg0_3,OutputImg0_2,OutputImg0_1,
              OutputImg0_0}), .OutputImg1 ({\$dummy [800],\$dummy [801],
              \$dummy [802],\$dummy [803],\$dummy [804],\$dummy [805],
              \$dummy [806],\$dummy [807],\$dummy [808],\$dummy [809],
              \$dummy [810],\$dummy [811],\$dummy [812],\$dummy [813],
              \$dummy [814],\$dummy [815],\$dummy [816],\$dummy [817],
              \$dummy [818],\$dummy [819],\$dummy [820],\$dummy [821],
              \$dummy [822],\$dummy [823],\$dummy [824],\$dummy [825],
              \$dummy [826],\$dummy [827],\$dummy [828],\$dummy [829],
              \$dummy [830],\$dummy [831],\$dummy [832],\$dummy [833],
              \$dummy [834],\$dummy [835],\$dummy [836],\$dummy [837],
              \$dummy [838],\$dummy [839],\$dummy [840],\$dummy [841],
              \$dummy [842],\$dummy [843],\$dummy [844],\$dummy [845],
              \$dummy [846],\$dummy [847],\$dummy [848],\$dummy [849],
              \$dummy [850],\$dummy [851],\$dummy [852],\$dummy [853],
              \$dummy [854],\$dummy [855],\$dummy [856],\$dummy [857],
              \$dummy [858],\$dummy [859],\$dummy [860],\$dummy [861],
              \$dummy [862],\$dummy [863],\$dummy [864],\$dummy [865],
              \$dummy [866],\$dummy [867],\$dummy [868],\$dummy [869],
              \$dummy [870],\$dummy [871],\$dummy [872],\$dummy [873],
              \$dummy [874],\$dummy [875],\$dummy [876],\$dummy [877],
              \$dummy [878],\$dummy [879],\$dummy [880],\$dummy [881],
              \$dummy [882],\$dummy [883],\$dummy [884],\$dummy [885],
              \$dummy [886],\$dummy [887],\$dummy [888],\$dummy [889],
              \$dummy [890],\$dummy [891],\$dummy [892],\$dummy [893],
              \$dummy [894],\$dummy [895],\$dummy [896],\$dummy [897],
              \$dummy [898],\$dummy [899],\$dummy [900],\$dummy [901],
              \$dummy [902],\$dummy [903],\$dummy [904],\$dummy [905],
              \$dummy [906],\$dummy [907],\$dummy [908],\$dummy [909],
              \$dummy [910],\$dummy [911],\$dummy [912],\$dummy [913],
              \$dummy [914],\$dummy [915],\$dummy [916],\$dummy [917],
              \$dummy [918],\$dummy [919],\$dummy [920],\$dummy [921],
              \$dummy [922],\$dummy [923],\$dummy [924],\$dummy [925],
              \$dummy [926],\$dummy [927],\$dummy [928],\$dummy [929],
              \$dummy [930],\$dummy [931],\$dummy [932],\$dummy [933],
              \$dummy [934],\$dummy [935],\$dummy [936],\$dummy [937],
              \$dummy [938],\$dummy [939],\$dummy [940],\$dummy [941],
              \$dummy [942],\$dummy [943],\$dummy [944],\$dummy [945],
              \$dummy [946],\$dummy [947],\$dummy [948],\$dummy [949],
              \$dummy [950],\$dummy [951],\$dummy [952],\$dummy [953],
              \$dummy [954],\$dummy [955],\$dummy [956],\$dummy [957],
              \$dummy [958],\$dummy [959],\$dummy [960],\$dummy [961],
              \$dummy [962],\$dummy [963],\$dummy [964],\$dummy [965],
              \$dummy [966],\$dummy [967],\$dummy [968],\$dummy [969],
              \$dummy [970],\$dummy [971],\$dummy [972],\$dummy [973],
              \$dummy [974],\$dummy [975],\$dummy [976],\$dummy [977],
              \$dummy [978],\$dummy [979],\$dummy [980],\$dummy [981],
              \$dummy [982],\$dummy [983],\$dummy [984],\$dummy [985],
              \$dummy [986],\$dummy [987],\$dummy [988],\$dummy [989],
              \$dummy [990],\$dummy [991],\$dummy [992],\$dummy [993],
              \$dummy [994],\$dummy [995],\$dummy [996],\$dummy [997],
              \$dummy [998],\$dummy [999],\$dummy [1000],\$dummy [1001],
              \$dummy [1002],\$dummy [1003],\$dummy [1004],\$dummy [1005],
              \$dummy [1006],\$dummy [1007],\$dummy [1008],\$dummy [1009],
              \$dummy [1010],\$dummy [1011],\$dummy [1012],\$dummy [1013],
              \$dummy [1014],\$dummy [1015],\$dummy [1016],\$dummy [1017],
              \$dummy [1018],\$dummy [1019],\$dummy [1020],\$dummy [1021],
              \$dummy [1022],\$dummy [1023],\$dummy [1024],\$dummy [1025],
              \$dummy [1026],\$dummy [1027],\$dummy [1028],\$dummy [1029],
              \$dummy [1030],\$dummy [1031],\$dummy [1032],\$dummy [1033],
              \$dummy [1034],\$dummy [1035],\$dummy [1036],\$dummy [1037],
              \$dummy [1038],\$dummy [1039],\$dummy [1040],\$dummy [1041],
              \$dummy [1042],\$dummy [1043],\$dummy [1044],\$dummy [1045],
              \$dummy [1046],\$dummy [1047],\$dummy [1048],\$dummy [1049],
              \$dummy [1050],\$dummy [1051],\$dummy [1052],\$dummy [1053],
              \$dummy [1054],\$dummy [1055],\$dummy [1056],\$dummy [1057],
              \$dummy [1058],\$dummy [1059],\$dummy [1060],\$dummy [1061],
              \$dummy [1062],\$dummy [1063],\$dummy [1064],\$dummy [1065],
              \$dummy [1066],\$dummy [1067],\$dummy [1068],\$dummy [1069],
              \$dummy [1070],\$dummy [1071],\$dummy [1072],\$dummy [1073],
              \$dummy [1074],\$dummy [1075],\$dummy [1076],\$dummy [1077],
              \$dummy [1078],\$dummy [1079],\$dummy [1080],\$dummy [1081],
              \$dummy [1082],\$dummy [1083],\$dummy [1084],\$dummy [1085],
              \$dummy [1086],\$dummy [1087],\$dummy [1088],\$dummy [1089],
              \$dummy [1090],\$dummy [1091],\$dummy [1092],\$dummy [1093],
              \$dummy [1094],\$dummy [1095],\$dummy [1096],\$dummy [1097],
              \$dummy [1098],\$dummy [1099],\$dummy [1100],\$dummy [1101],
              \$dummy [1102],\$dummy [1103],\$dummy [1104],\$dummy [1105],
              \$dummy [1106],\$dummy [1107],\$dummy [1108],\$dummy [1109],
              \$dummy [1110],\$dummy [1111],\$dummy [1112],\$dummy [1113],
              \$dummy [1114],\$dummy [1115],\$dummy [1116],\$dummy [1117],
              \$dummy [1118],\$dummy [1119],\$dummy [1120],\$dummy [1121],
              \$dummy [1122],\$dummy [1123],\$dummy [1124],\$dummy [1125],
              \$dummy [1126],\$dummy [1127],\$dummy [1128],\$dummy [1129],
              \$dummy [1130],\$dummy [1131],\$dummy [1132],\$dummy [1133],
              \$dummy [1134],\$dummy [1135],\$dummy [1136],\$dummy [1137],
              \$dummy [1138],\$dummy [1139],\$dummy [1140],\$dummy [1141],
              \$dummy [1142],\$dummy [1143],\$dummy [1144],\$dummy [1145],
              \$dummy [1146],\$dummy [1147],\$dummy [1148],\$dummy [1149],
              \$dummy [1150],\$dummy [1151],\$dummy [1152],\$dummy [1153],
              \$dummy [1154],\$dummy [1155],\$dummy [1156],\$dummy [1157],
              \$dummy [1158],\$dummy [1159],\$dummy [1160],\$dummy [1161],
              \$dummy [1162],\$dummy [1163],\$dummy [1164],\$dummy [1165],
              \$dummy [1166],\$dummy [1167],OutputImg1_79,OutputImg1_78,
              OutputImg1_77,OutputImg1_76,OutputImg1_75,OutputImg1_74,
              OutputImg1_73,OutputImg1_72,OutputImg1_71,OutputImg1_70,
              OutputImg1_69,OutputImg1_68,OutputImg1_67,OutputImg1_66,
              OutputImg1_65,OutputImg1_64,OutputImg1_63,OutputImg1_62,
              OutputImg1_61,OutputImg1_60,OutputImg1_59,OutputImg1_58,
              OutputImg1_57,OutputImg1_56,OutputImg1_55,OutputImg1_54,
              OutputImg1_53,OutputImg1_52,OutputImg1_51,OutputImg1_50,
              OutputImg1_49,OutputImg1_48,OutputImg1_47,OutputImg1_46,
              OutputImg1_45,OutputImg1_44,OutputImg1_43,OutputImg1_42,
              OutputImg1_41,OutputImg1_40,OutputImg1_39,OutputImg1_38,
              OutputImg1_37,OutputImg1_36,OutputImg1_35,OutputImg1_34,
              OutputImg1_33,OutputImg1_32,OutputImg1_31,OutputImg1_30,
              OutputImg1_29,OutputImg1_28,OutputImg1_27,OutputImg1_26,
              OutputImg1_25,OutputImg1_24,OutputImg1_23,OutputImg1_22,
              OutputImg1_21,OutputImg1_20,OutputImg1_19,OutputImg1_18,
              OutputImg1_17,OutputImg1_16,OutputImg1_15,OutputImg1_14,
              OutputImg1_13,OutputImg1_12,OutputImg1_11,OutputImg1_10,
              OutputImg1_9,OutputImg1_8,OutputImg1_7,OutputImg1_6,OutputImg1_5,
              OutputImg1_4,OutputImg1_3,OutputImg1_2,OutputImg1_1,OutputImg1_0})
              , .OutputImg2 ({\$dummy [1168],\$dummy [1169],\$dummy [1170],
              \$dummy [1171],\$dummy [1172],\$dummy [1173],\$dummy [1174],
              \$dummy [1175],\$dummy [1176],\$dummy [1177],\$dummy [1178],
              \$dummy [1179],\$dummy [1180],\$dummy [1181],\$dummy [1182],
              \$dummy [1183],\$dummy [1184],\$dummy [1185],\$dummy [1186],
              \$dummy [1187],\$dummy [1188],\$dummy [1189],\$dummy [1190],
              \$dummy [1191],\$dummy [1192],\$dummy [1193],\$dummy [1194],
              \$dummy [1195],\$dummy [1196],\$dummy [1197],\$dummy [1198],
              \$dummy [1199],\$dummy [1200],\$dummy [1201],\$dummy [1202],
              \$dummy [1203],\$dummy [1204],\$dummy [1205],\$dummy [1206],
              \$dummy [1207],\$dummy [1208],\$dummy [1209],\$dummy [1210],
              \$dummy [1211],\$dummy [1212],\$dummy [1213],\$dummy [1214],
              \$dummy [1215],\$dummy [1216],\$dummy [1217],\$dummy [1218],
              \$dummy [1219],\$dummy [1220],\$dummy [1221],\$dummy [1222],
              \$dummy [1223],\$dummy [1224],\$dummy [1225],\$dummy [1226],
              \$dummy [1227],\$dummy [1228],\$dummy [1229],\$dummy [1230],
              \$dummy [1231],\$dummy [1232],\$dummy [1233],\$dummy [1234],
              \$dummy [1235],\$dummy [1236],\$dummy [1237],\$dummy [1238],
              \$dummy [1239],\$dummy [1240],\$dummy [1241],\$dummy [1242],
              \$dummy [1243],\$dummy [1244],\$dummy [1245],\$dummy [1246],
              \$dummy [1247],\$dummy [1248],\$dummy [1249],\$dummy [1250],
              \$dummy [1251],\$dummy [1252],\$dummy [1253],\$dummy [1254],
              \$dummy [1255],\$dummy [1256],\$dummy [1257],\$dummy [1258],
              \$dummy [1259],\$dummy [1260],\$dummy [1261],\$dummy [1262],
              \$dummy [1263],\$dummy [1264],\$dummy [1265],\$dummy [1266],
              \$dummy [1267],\$dummy [1268],\$dummy [1269],\$dummy [1270],
              \$dummy [1271],\$dummy [1272],\$dummy [1273],\$dummy [1274],
              \$dummy [1275],\$dummy [1276],\$dummy [1277],\$dummy [1278],
              \$dummy [1279],\$dummy [1280],\$dummy [1281],\$dummy [1282],
              \$dummy [1283],\$dummy [1284],\$dummy [1285],\$dummy [1286],
              \$dummy [1287],\$dummy [1288],\$dummy [1289],\$dummy [1290],
              \$dummy [1291],\$dummy [1292],\$dummy [1293],\$dummy [1294],
              \$dummy [1295],\$dummy [1296],\$dummy [1297],\$dummy [1298],
              \$dummy [1299],\$dummy [1300],\$dummy [1301],\$dummy [1302],
              \$dummy [1303],\$dummy [1304],\$dummy [1305],\$dummy [1306],
              \$dummy [1307],\$dummy [1308],\$dummy [1309],\$dummy [1310],
              \$dummy [1311],\$dummy [1312],\$dummy [1313],\$dummy [1314],
              \$dummy [1315],\$dummy [1316],\$dummy [1317],\$dummy [1318],
              \$dummy [1319],\$dummy [1320],\$dummy [1321],\$dummy [1322],
              \$dummy [1323],\$dummy [1324],\$dummy [1325],\$dummy [1326],
              \$dummy [1327],\$dummy [1328],\$dummy [1329],\$dummy [1330],
              \$dummy [1331],\$dummy [1332],\$dummy [1333],\$dummy [1334],
              \$dummy [1335],\$dummy [1336],\$dummy [1337],\$dummy [1338],
              \$dummy [1339],\$dummy [1340],\$dummy [1341],\$dummy [1342],
              \$dummy [1343],\$dummy [1344],\$dummy [1345],\$dummy [1346],
              \$dummy [1347],\$dummy [1348],\$dummy [1349],\$dummy [1350],
              \$dummy [1351],\$dummy [1352],\$dummy [1353],\$dummy [1354],
              \$dummy [1355],\$dummy [1356],\$dummy [1357],\$dummy [1358],
              \$dummy [1359],\$dummy [1360],\$dummy [1361],\$dummy [1362],
              \$dummy [1363],\$dummy [1364],\$dummy [1365],\$dummy [1366],
              \$dummy [1367],\$dummy [1368],\$dummy [1369],\$dummy [1370],
              \$dummy [1371],\$dummy [1372],\$dummy [1373],\$dummy [1374],
              \$dummy [1375],\$dummy [1376],\$dummy [1377],\$dummy [1378],
              \$dummy [1379],\$dummy [1380],\$dummy [1381],\$dummy [1382],
              \$dummy [1383],\$dummy [1384],\$dummy [1385],\$dummy [1386],
              \$dummy [1387],\$dummy [1388],\$dummy [1389],\$dummy [1390],
              \$dummy [1391],\$dummy [1392],\$dummy [1393],\$dummy [1394],
              \$dummy [1395],\$dummy [1396],\$dummy [1397],\$dummy [1398],
              \$dummy [1399],\$dummy [1400],\$dummy [1401],\$dummy [1402],
              \$dummy [1403],\$dummy [1404],\$dummy [1405],\$dummy [1406],
              \$dummy [1407],\$dummy [1408],\$dummy [1409],\$dummy [1410],
              \$dummy [1411],\$dummy [1412],\$dummy [1413],\$dummy [1414],
              \$dummy [1415],\$dummy [1416],\$dummy [1417],\$dummy [1418],
              \$dummy [1419],\$dummy [1420],\$dummy [1421],\$dummy [1422],
              \$dummy [1423],\$dummy [1424],\$dummy [1425],\$dummy [1426],
              \$dummy [1427],\$dummy [1428],\$dummy [1429],\$dummy [1430],
              \$dummy [1431],\$dummy [1432],\$dummy [1433],\$dummy [1434],
              \$dummy [1435],\$dummy [1436],\$dummy [1437],\$dummy [1438],
              \$dummy [1439],\$dummy [1440],\$dummy [1441],\$dummy [1442],
              \$dummy [1443],\$dummy [1444],\$dummy [1445],\$dummy [1446],
              \$dummy [1447],\$dummy [1448],\$dummy [1449],\$dummy [1450],
              \$dummy [1451],\$dummy [1452],\$dummy [1453],\$dummy [1454],
              \$dummy [1455],\$dummy [1456],\$dummy [1457],\$dummy [1458],
              \$dummy [1459],\$dummy [1460],\$dummy [1461],\$dummy [1462],
              \$dummy [1463],\$dummy [1464],\$dummy [1465],\$dummy [1466],
              \$dummy [1467],\$dummy [1468],\$dummy [1469],\$dummy [1470],
              \$dummy [1471],\$dummy [1472],\$dummy [1473],\$dummy [1474],
              \$dummy [1475],\$dummy [1476],\$dummy [1477],\$dummy [1478],
              \$dummy [1479],\$dummy [1480],\$dummy [1481],\$dummy [1482],
              \$dummy [1483],\$dummy [1484],\$dummy [1485],\$dummy [1486],
              \$dummy [1487],\$dummy [1488],\$dummy [1489],\$dummy [1490],
              \$dummy [1491],\$dummy [1492],\$dummy [1493],\$dummy [1494],
              \$dummy [1495],\$dummy [1496],\$dummy [1497],\$dummy [1498],
              \$dummy [1499],\$dummy [1500],\$dummy [1501],\$dummy [1502],
              \$dummy [1503],\$dummy [1504],\$dummy [1505],\$dummy [1506],
              \$dummy [1507],\$dummy [1508],\$dummy [1509],\$dummy [1510],
              \$dummy [1511],\$dummy [1512],\$dummy [1513],\$dummy [1514],
              \$dummy [1515],\$dummy [1516],\$dummy [1517],\$dummy [1518],
              \$dummy [1519],\$dummy [1520],\$dummy [1521],\$dummy [1522],
              \$dummy [1523],\$dummy [1524],\$dummy [1525],\$dummy [1526],
              \$dummy [1527],\$dummy [1528],\$dummy [1529],\$dummy [1530],
              \$dummy [1531],\$dummy [1532],\$dummy [1533],\$dummy [1534],
              \$dummy [1535],OutputImg2_79,OutputImg2_78,OutputImg2_77,
              OutputImg2_76,OutputImg2_75,OutputImg2_74,OutputImg2_73,
              OutputImg2_72,OutputImg2_71,OutputImg2_70,OutputImg2_69,
              OutputImg2_68,OutputImg2_67,OutputImg2_66,OutputImg2_65,
              OutputImg2_64,OutputImg2_63,OutputImg2_62,OutputImg2_61,
              OutputImg2_60,OutputImg2_59,OutputImg2_58,OutputImg2_57,
              OutputImg2_56,OutputImg2_55,OutputImg2_54,OutputImg2_53,
              OutputImg2_52,OutputImg2_51,OutputImg2_50,OutputImg2_49,
              OutputImg2_48,OutputImg2_47,OutputImg2_46,OutputImg2_45,
              OutputImg2_44,OutputImg2_43,OutputImg2_42,OutputImg2_41,
              OutputImg2_40,OutputImg2_39,OutputImg2_38,OutputImg2_37,
              OutputImg2_36,OutputImg2_35,OutputImg2_34,OutputImg2_33,
              OutputImg2_32,OutputImg2_31,OutputImg2_30,OutputImg2_29,
              OutputImg2_28,OutputImg2_27,OutputImg2_26,OutputImg2_25,
              OutputImg2_24,OutputImg2_23,OutputImg2_22,OutputImg2_21,
              OutputImg2_20,OutputImg2_19,OutputImg2_18,OutputImg2_17,
              OutputImg2_16,OutputImg2_15,OutputImg2_14,OutputImg2_13,
              OutputImg2_12,OutputImg2_11,OutputImg2_10,OutputImg2_9,
              OutputImg2_8,OutputImg2_7,OutputImg2_6,OutputImg2_5,OutputImg2_4,
              OutputImg2_3,OutputImg2_2,OutputImg2_1,OutputImg2_0}), .OutputImg3 (
              {\$dummy [1536],\$dummy [1537],\$dummy [1538],\$dummy [1539],
              \$dummy [1540],\$dummy [1541],\$dummy [1542],\$dummy [1543],
              \$dummy [1544],\$dummy [1545],\$dummy [1546],\$dummy [1547],
              \$dummy [1548],\$dummy [1549],\$dummy [1550],\$dummy [1551],
              \$dummy [1552],\$dummy [1553],\$dummy [1554],\$dummy [1555],
              \$dummy [1556],\$dummy [1557],\$dummy [1558],\$dummy [1559],
              \$dummy [1560],\$dummy [1561],\$dummy [1562],\$dummy [1563],
              \$dummy [1564],\$dummy [1565],\$dummy [1566],\$dummy [1567],
              \$dummy [1568],\$dummy [1569],\$dummy [1570],\$dummy [1571],
              \$dummy [1572],\$dummy [1573],\$dummy [1574],\$dummy [1575],
              \$dummy [1576],\$dummy [1577],\$dummy [1578],\$dummy [1579],
              \$dummy [1580],\$dummy [1581],\$dummy [1582],\$dummy [1583],
              \$dummy [1584],\$dummy [1585],\$dummy [1586],\$dummy [1587],
              \$dummy [1588],\$dummy [1589],\$dummy [1590],\$dummy [1591],
              \$dummy [1592],\$dummy [1593],\$dummy [1594],\$dummy [1595],
              \$dummy [1596],\$dummy [1597],\$dummy [1598],\$dummy [1599],
              \$dummy [1600],\$dummy [1601],\$dummy [1602],\$dummy [1603],
              \$dummy [1604],\$dummy [1605],\$dummy [1606],\$dummy [1607],
              \$dummy [1608],\$dummy [1609],\$dummy [1610],\$dummy [1611],
              \$dummy [1612],\$dummy [1613],\$dummy [1614],\$dummy [1615],
              \$dummy [1616],\$dummy [1617],\$dummy [1618],\$dummy [1619],
              \$dummy [1620],\$dummy [1621],\$dummy [1622],\$dummy [1623],
              \$dummy [1624],\$dummy [1625],\$dummy [1626],\$dummy [1627],
              \$dummy [1628],\$dummy [1629],\$dummy [1630],\$dummy [1631],
              \$dummy [1632],\$dummy [1633],\$dummy [1634],\$dummy [1635],
              \$dummy [1636],\$dummy [1637],\$dummy [1638],\$dummy [1639],
              \$dummy [1640],\$dummy [1641],\$dummy [1642],\$dummy [1643],
              \$dummy [1644],\$dummy [1645],\$dummy [1646],\$dummy [1647],
              \$dummy [1648],\$dummy [1649],\$dummy [1650],\$dummy [1651],
              \$dummy [1652],\$dummy [1653],\$dummy [1654],\$dummy [1655],
              \$dummy [1656],\$dummy [1657],\$dummy [1658],\$dummy [1659],
              \$dummy [1660],\$dummy [1661],\$dummy [1662],\$dummy [1663],
              \$dummy [1664],\$dummy [1665],\$dummy [1666],\$dummy [1667],
              \$dummy [1668],\$dummy [1669],\$dummy [1670],\$dummy [1671],
              \$dummy [1672],\$dummy [1673],\$dummy [1674],\$dummy [1675],
              \$dummy [1676],\$dummy [1677],\$dummy [1678],\$dummy [1679],
              \$dummy [1680],\$dummy [1681],\$dummy [1682],\$dummy [1683],
              \$dummy [1684],\$dummy [1685],\$dummy [1686],\$dummy [1687],
              \$dummy [1688],\$dummy [1689],\$dummy [1690],\$dummy [1691],
              \$dummy [1692],\$dummy [1693],\$dummy [1694],\$dummy [1695],
              \$dummy [1696],\$dummy [1697],\$dummy [1698],\$dummy [1699],
              \$dummy [1700],\$dummy [1701],\$dummy [1702],\$dummy [1703],
              \$dummy [1704],\$dummy [1705],\$dummy [1706],\$dummy [1707],
              \$dummy [1708],\$dummy [1709],\$dummy [1710],\$dummy [1711],
              \$dummy [1712],\$dummy [1713],\$dummy [1714],\$dummy [1715],
              \$dummy [1716],\$dummy [1717],\$dummy [1718],\$dummy [1719],
              \$dummy [1720],\$dummy [1721],\$dummy [1722],\$dummy [1723],
              \$dummy [1724],\$dummy [1725],\$dummy [1726],\$dummy [1727],
              \$dummy [1728],\$dummy [1729],\$dummy [1730],\$dummy [1731],
              \$dummy [1732],\$dummy [1733],\$dummy [1734],\$dummy [1735],
              \$dummy [1736],\$dummy [1737],\$dummy [1738],\$dummy [1739],
              \$dummy [1740],\$dummy [1741],\$dummy [1742],\$dummy [1743],
              \$dummy [1744],\$dummy [1745],\$dummy [1746],\$dummy [1747],
              \$dummy [1748],\$dummy [1749],\$dummy [1750],\$dummy [1751],
              \$dummy [1752],\$dummy [1753],\$dummy [1754],\$dummy [1755],
              \$dummy [1756],\$dummy [1757],\$dummy [1758],\$dummy [1759],
              \$dummy [1760],\$dummy [1761],\$dummy [1762],\$dummy [1763],
              \$dummy [1764],\$dummy [1765],\$dummy [1766],\$dummy [1767],
              \$dummy [1768],\$dummy [1769],\$dummy [1770],\$dummy [1771],
              \$dummy [1772],\$dummy [1773],\$dummy [1774],\$dummy [1775],
              \$dummy [1776],\$dummy [1777],\$dummy [1778],\$dummy [1779],
              \$dummy [1780],\$dummy [1781],\$dummy [1782],\$dummy [1783],
              \$dummy [1784],\$dummy [1785],\$dummy [1786],\$dummy [1787],
              \$dummy [1788],\$dummy [1789],\$dummy [1790],\$dummy [1791],
              \$dummy [1792],\$dummy [1793],\$dummy [1794],\$dummy [1795],
              \$dummy [1796],\$dummy [1797],\$dummy [1798],\$dummy [1799],
              \$dummy [1800],\$dummy [1801],\$dummy [1802],\$dummy [1803],
              \$dummy [1804],\$dummy [1805],\$dummy [1806],\$dummy [1807],
              \$dummy [1808],\$dummy [1809],\$dummy [1810],\$dummy [1811],
              \$dummy [1812],\$dummy [1813],\$dummy [1814],\$dummy [1815],
              \$dummy [1816],\$dummy [1817],\$dummy [1818],\$dummy [1819],
              \$dummy [1820],\$dummy [1821],\$dummy [1822],\$dummy [1823],
              \$dummy [1824],\$dummy [1825],\$dummy [1826],\$dummy [1827],
              \$dummy [1828],\$dummy [1829],\$dummy [1830],\$dummy [1831],
              \$dummy [1832],\$dummy [1833],\$dummy [1834],\$dummy [1835],
              \$dummy [1836],\$dummy [1837],\$dummy [1838],\$dummy [1839],
              \$dummy [1840],\$dummy [1841],\$dummy [1842],\$dummy [1843],
              \$dummy [1844],\$dummy [1845],\$dummy [1846],\$dummy [1847],
              \$dummy [1848],\$dummy [1849],\$dummy [1850],\$dummy [1851],
              \$dummy [1852],\$dummy [1853],\$dummy [1854],\$dummy [1855],
              \$dummy [1856],\$dummy [1857],\$dummy [1858],\$dummy [1859],
              \$dummy [1860],\$dummy [1861],\$dummy [1862],\$dummy [1863],
              \$dummy [1864],\$dummy [1865],\$dummy [1866],\$dummy [1867],
              \$dummy [1868],\$dummy [1869],\$dummy [1870],\$dummy [1871],
              \$dummy [1872],\$dummy [1873],\$dummy [1874],\$dummy [1875],
              \$dummy [1876],\$dummy [1877],\$dummy [1878],\$dummy [1879],
              \$dummy [1880],\$dummy [1881],\$dummy [1882],\$dummy [1883],
              \$dummy [1884],\$dummy [1885],\$dummy [1886],\$dummy [1887],
              \$dummy [1888],\$dummy [1889],\$dummy [1890],\$dummy [1891],
              \$dummy [1892],\$dummy [1893],\$dummy [1894],\$dummy [1895],
              \$dummy [1896],\$dummy [1897],\$dummy [1898],\$dummy [1899],
              \$dummy [1900],\$dummy [1901],\$dummy [1902],\$dummy [1903],
              OutputImg3_79,OutputImg3_78,OutputImg3_77,OutputImg3_76,
              OutputImg3_75,OutputImg3_74,OutputImg3_73,OutputImg3_72,
              OutputImg3_71,OutputImg3_70,OutputImg3_69,OutputImg3_68,
              OutputImg3_67,OutputImg3_66,OutputImg3_65,OutputImg3_64,
              OutputImg3_63,OutputImg3_62,OutputImg3_61,OutputImg3_60,
              OutputImg3_59,OutputImg3_58,OutputImg3_57,OutputImg3_56,
              OutputImg3_55,OutputImg3_54,OutputImg3_53,OutputImg3_52,
              OutputImg3_51,OutputImg3_50,OutputImg3_49,OutputImg3_48,
              OutputImg3_47,OutputImg3_46,OutputImg3_45,OutputImg3_44,
              OutputImg3_43,OutputImg3_42,OutputImg3_41,OutputImg3_40,
              OutputImg3_39,OutputImg3_38,OutputImg3_37,OutputImg3_36,
              OutputImg3_35,OutputImg3_34,OutputImg3_33,OutputImg3_32,
              OutputImg3_31,OutputImg3_30,OutputImg3_29,OutputImg3_28,
              OutputImg3_27,OutputImg3_26,OutputImg3_25,OutputImg3_24,
              OutputImg3_23,OutputImg3_22,OutputImg3_21,OutputImg3_20,
              OutputImg3_19,OutputImg3_18,OutputImg3_17,OutputImg3_16,
              OutputImg3_15,OutputImg3_14,OutputImg3_13,OutputImg3_12,
              OutputImg3_11,OutputImg3_10,OutputImg3_9,OutputImg3_8,OutputImg3_7
              ,OutputImg3_6,OutputImg3_5,OutputImg3_4,OutputImg3_3,OutputImg3_2,
              OutputImg3_1,OutputImg3_0}), .OutputImg4 ({\$dummy [1904],
              \$dummy [1905],\$dummy [1906],\$dummy [1907],\$dummy [1908],
              \$dummy [1909],\$dummy [1910],\$dummy [1911],\$dummy [1912],
              \$dummy [1913],\$dummy [1914],\$dummy [1915],\$dummy [1916],
              \$dummy [1917],\$dummy [1918],\$dummy [1919],\$dummy [1920],
              \$dummy [1921],\$dummy [1922],\$dummy [1923],\$dummy [1924],
              \$dummy [1925],\$dummy [1926],\$dummy [1927],\$dummy [1928],
              \$dummy [1929],\$dummy [1930],\$dummy [1931],\$dummy [1932],
              \$dummy [1933],\$dummy [1934],\$dummy [1935],\$dummy [1936],
              \$dummy [1937],\$dummy [1938],\$dummy [1939],\$dummy [1940],
              \$dummy [1941],\$dummy [1942],\$dummy [1943],\$dummy [1944],
              \$dummy [1945],\$dummy [1946],\$dummy [1947],\$dummy [1948],
              \$dummy [1949],\$dummy [1950],\$dummy [1951],\$dummy [1952],
              \$dummy [1953],\$dummy [1954],\$dummy [1955],\$dummy [1956],
              \$dummy [1957],\$dummy [1958],\$dummy [1959],\$dummy [1960],
              \$dummy [1961],\$dummy [1962],\$dummy [1963],\$dummy [1964],
              \$dummy [1965],\$dummy [1966],\$dummy [1967],\$dummy [1968],
              \$dummy [1969],\$dummy [1970],\$dummy [1971],\$dummy [1972],
              \$dummy [1973],\$dummy [1974],\$dummy [1975],\$dummy [1976],
              \$dummy [1977],\$dummy [1978],\$dummy [1979],\$dummy [1980],
              \$dummy [1981],\$dummy [1982],\$dummy [1983],\$dummy [1984],
              \$dummy [1985],\$dummy [1986],\$dummy [1987],\$dummy [1988],
              \$dummy [1989],\$dummy [1990],\$dummy [1991],\$dummy [1992],
              \$dummy [1993],\$dummy [1994],\$dummy [1995],\$dummy [1996],
              \$dummy [1997],\$dummy [1998],\$dummy [1999],\$dummy [2000],
              \$dummy [2001],\$dummy [2002],\$dummy [2003],\$dummy [2004],
              \$dummy [2005],\$dummy [2006],\$dummy [2007],\$dummy [2008],
              \$dummy [2009],\$dummy [2010],\$dummy [2011],\$dummy [2012],
              \$dummy [2013],\$dummy [2014],\$dummy [2015],\$dummy [2016],
              \$dummy [2017],\$dummy [2018],\$dummy [2019],\$dummy [2020],
              \$dummy [2021],\$dummy [2022],\$dummy [2023],\$dummy [2024],
              \$dummy [2025],\$dummy [2026],\$dummy [2027],\$dummy [2028],
              \$dummy [2029],\$dummy [2030],\$dummy [2031],\$dummy [2032],
              \$dummy [2033],\$dummy [2034],\$dummy [2035],\$dummy [2036],
              \$dummy [2037],\$dummy [2038],\$dummy [2039],\$dummy [2040],
              \$dummy [2041],\$dummy [2042],\$dummy [2043],\$dummy [2044],
              \$dummy [2045],\$dummy [2046],\$dummy [2047],\$dummy [2048],
              \$dummy [2049],\$dummy [2050],\$dummy [2051],\$dummy [2052],
              \$dummy [2053],\$dummy [2054],\$dummy [2055],\$dummy [2056],
              \$dummy [2057],\$dummy [2058],\$dummy [2059],\$dummy [2060],
              \$dummy [2061],\$dummy [2062],\$dummy [2063],\$dummy [2064],
              \$dummy [2065],\$dummy [2066],\$dummy [2067],\$dummy [2068],
              \$dummy [2069],\$dummy [2070],\$dummy [2071],\$dummy [2072],
              \$dummy [2073],\$dummy [2074],\$dummy [2075],\$dummy [2076],
              \$dummy [2077],\$dummy [2078],\$dummy [2079],\$dummy [2080],
              \$dummy [2081],\$dummy [2082],\$dummy [2083],\$dummy [2084],
              \$dummy [2085],\$dummy [2086],\$dummy [2087],\$dummy [2088],
              \$dummy [2089],\$dummy [2090],\$dummy [2091],\$dummy [2092],
              \$dummy [2093],\$dummy [2094],\$dummy [2095],\$dummy [2096],
              \$dummy [2097],\$dummy [2098],\$dummy [2099],\$dummy [2100],
              \$dummy [2101],\$dummy [2102],\$dummy [2103],\$dummy [2104],
              \$dummy [2105],\$dummy [2106],\$dummy [2107],\$dummy [2108],
              \$dummy [2109],\$dummy [2110],\$dummy [2111],\$dummy [2112],
              \$dummy [2113],\$dummy [2114],\$dummy [2115],\$dummy [2116],
              \$dummy [2117],\$dummy [2118],\$dummy [2119],\$dummy [2120],
              \$dummy [2121],\$dummy [2122],\$dummy [2123],\$dummy [2124],
              \$dummy [2125],\$dummy [2126],\$dummy [2127],\$dummy [2128],
              \$dummy [2129],\$dummy [2130],\$dummy [2131],\$dummy [2132],
              \$dummy [2133],\$dummy [2134],\$dummy [2135],\$dummy [2136],
              \$dummy [2137],\$dummy [2138],\$dummy [2139],\$dummy [2140],
              \$dummy [2141],\$dummy [2142],\$dummy [2143],\$dummy [2144],
              \$dummy [2145],\$dummy [2146],\$dummy [2147],\$dummy [2148],
              \$dummy [2149],\$dummy [2150],\$dummy [2151],\$dummy [2152],
              \$dummy [2153],\$dummy [2154],\$dummy [2155],\$dummy [2156],
              \$dummy [2157],\$dummy [2158],\$dummy [2159],\$dummy [2160],
              \$dummy [2161],\$dummy [2162],\$dummy [2163],\$dummy [2164],
              \$dummy [2165],\$dummy [2166],\$dummy [2167],\$dummy [2168],
              \$dummy [2169],\$dummy [2170],\$dummy [2171],\$dummy [2172],
              \$dummy [2173],\$dummy [2174],\$dummy [2175],\$dummy [2176],
              \$dummy [2177],\$dummy [2178],\$dummy [2179],\$dummy [2180],
              \$dummy [2181],\$dummy [2182],\$dummy [2183],\$dummy [2184],
              \$dummy [2185],\$dummy [2186],\$dummy [2187],\$dummy [2188],
              \$dummy [2189],\$dummy [2190],\$dummy [2191],\$dummy [2192],
              \$dummy [2193],\$dummy [2194],\$dummy [2195],\$dummy [2196],
              \$dummy [2197],\$dummy [2198],\$dummy [2199],\$dummy [2200],
              \$dummy [2201],\$dummy [2202],\$dummy [2203],\$dummy [2204],
              \$dummy [2205],\$dummy [2206],\$dummy [2207],\$dummy [2208],
              \$dummy [2209],\$dummy [2210],\$dummy [2211],\$dummy [2212],
              \$dummy [2213],\$dummy [2214],\$dummy [2215],\$dummy [2216],
              \$dummy [2217],\$dummy [2218],\$dummy [2219],\$dummy [2220],
              \$dummy [2221],\$dummy [2222],\$dummy [2223],\$dummy [2224],
              \$dummy [2225],\$dummy [2226],\$dummy [2227],\$dummy [2228],
              \$dummy [2229],\$dummy [2230],\$dummy [2231],\$dummy [2232],
              \$dummy [2233],\$dummy [2234],\$dummy [2235],\$dummy [2236],
              \$dummy [2237],\$dummy [2238],\$dummy [2239],\$dummy [2240],
              \$dummy [2241],\$dummy [2242],\$dummy [2243],\$dummy [2244],
              \$dummy [2245],\$dummy [2246],\$dummy [2247],\$dummy [2248],
              \$dummy [2249],\$dummy [2250],\$dummy [2251],\$dummy [2252],
              \$dummy [2253],\$dummy [2254],\$dummy [2255],\$dummy [2256],
              \$dummy [2257],\$dummy [2258],\$dummy [2259],\$dummy [2260],
              \$dummy [2261],\$dummy [2262],\$dummy [2263],\$dummy [2264],
              \$dummy [2265],\$dummy [2266],\$dummy [2267],\$dummy [2268],
              \$dummy [2269],\$dummy [2270],\$dummy [2271],OutputImg4_79,
              OutputImg4_78,OutputImg4_77,OutputImg4_76,OutputImg4_75,
              OutputImg4_74,OutputImg4_73,OutputImg4_72,OutputImg4_71,
              OutputImg4_70,OutputImg4_69,OutputImg4_68,OutputImg4_67,
              OutputImg4_66,OutputImg4_65,OutputImg4_64,OutputImg4_63,
              OutputImg4_62,OutputImg4_61,OutputImg4_60,OutputImg4_59,
              OutputImg4_58,OutputImg4_57,OutputImg4_56,OutputImg4_55,
              OutputImg4_54,OutputImg4_53,OutputImg4_52,OutputImg4_51,
              OutputImg4_50,OutputImg4_49,OutputImg4_48,OutputImg4_47,
              OutputImg4_46,OutputImg4_45,OutputImg4_44,OutputImg4_43,
              OutputImg4_42,OutputImg4_41,OutputImg4_40,OutputImg4_39,
              OutputImg4_38,OutputImg4_37,OutputImg4_36,OutputImg4_35,
              OutputImg4_34,OutputImg4_33,OutputImg4_32,OutputImg4_31,
              OutputImg4_30,OutputImg4_29,OutputImg4_28,OutputImg4_27,
              OutputImg4_26,OutputImg4_25,OutputImg4_24,OutputImg4_23,
              OutputImg4_22,OutputImg4_21,OutputImg4_20,OutputImg4_19,
              OutputImg4_18,OutputImg4_17,OutputImg4_16,OutputImg4_15,
              OutputImg4_14,OutputImg4_13,OutputImg4_12,OutputImg4_11,
              OutputImg4_10,OutputImg4_9,OutputImg4_8,OutputImg4_7,OutputImg4_6,
              OutputImg4_5,OutputImg4_4,OutputImg4_3,OutputImg4_2,OutputImg4_1,
              OutputImg4_0}), .OutputImg5 ({\$dummy [2272],\$dummy [2273],
              \$dummy [2274],\$dummy [2275],\$dummy [2276],\$dummy [2277],
              \$dummy [2278],\$dummy [2279],\$dummy [2280],\$dummy [2281],
              \$dummy [2282],\$dummy [2283],\$dummy [2284],\$dummy [2285],
              \$dummy [2286],\$dummy [2287],\$dummy [2288],\$dummy [2289],
              \$dummy [2290],\$dummy [2291],\$dummy [2292],\$dummy [2293],
              \$dummy [2294],\$dummy [2295],\$dummy [2296],\$dummy [2297],
              \$dummy [2298],\$dummy [2299],\$dummy [2300],\$dummy [2301],
              \$dummy [2302],\$dummy [2303],\$dummy [2304],\$dummy [2305],
              \$dummy [2306],\$dummy [2307],\$dummy [2308],\$dummy [2309],
              \$dummy [2310],\$dummy [2311],\$dummy [2312],\$dummy [2313],
              \$dummy [2314],\$dummy [2315],\$dummy [2316],\$dummy [2317],
              \$dummy [2318],\$dummy [2319],\$dummy [2320],\$dummy [2321],
              \$dummy [2322],\$dummy [2323],\$dummy [2324],\$dummy [2325],
              \$dummy [2326],\$dummy [2327],\$dummy [2328],\$dummy [2329],
              \$dummy [2330],\$dummy [2331],\$dummy [2332],\$dummy [2333],
              \$dummy [2334],\$dummy [2335],\$dummy [2336],\$dummy [2337],
              \$dummy [2338],\$dummy [2339],\$dummy [2340],\$dummy [2341],
              \$dummy [2342],\$dummy [2343],\$dummy [2344],\$dummy [2345],
              \$dummy [2346],\$dummy [2347],\$dummy [2348],\$dummy [2349],
              \$dummy [2350],\$dummy [2351],\$dummy [2352],\$dummy [2353],
              \$dummy [2354],\$dummy [2355],\$dummy [2356],\$dummy [2357],
              \$dummy [2358],\$dummy [2359],\$dummy [2360],\$dummy [2361],
              \$dummy [2362],\$dummy [2363],\$dummy [2364],\$dummy [2365],
              \$dummy [2366],\$dummy [2367],\$dummy [2368],\$dummy [2369],
              \$dummy [2370],\$dummy [2371],\$dummy [2372],\$dummy [2373],
              \$dummy [2374],\$dummy [2375],\$dummy [2376],\$dummy [2377],
              \$dummy [2378],\$dummy [2379],\$dummy [2380],\$dummy [2381],
              \$dummy [2382],\$dummy [2383],\$dummy [2384],\$dummy [2385],
              \$dummy [2386],\$dummy [2387],\$dummy [2388],\$dummy [2389],
              \$dummy [2390],\$dummy [2391],\$dummy [2392],\$dummy [2393],
              \$dummy [2394],\$dummy [2395],\$dummy [2396],\$dummy [2397],
              \$dummy [2398],\$dummy [2399],\$dummy [2400],\$dummy [2401],
              \$dummy [2402],\$dummy [2403],\$dummy [2404],\$dummy [2405],
              \$dummy [2406],\$dummy [2407],\$dummy [2408],\$dummy [2409],
              \$dummy [2410],\$dummy [2411],\$dummy [2412],\$dummy [2413],
              \$dummy [2414],\$dummy [2415],\$dummy [2416],\$dummy [2417],
              \$dummy [2418],\$dummy [2419],\$dummy [2420],\$dummy [2421],
              \$dummy [2422],\$dummy [2423],\$dummy [2424],\$dummy [2425],
              \$dummy [2426],\$dummy [2427],\$dummy [2428],\$dummy [2429],
              \$dummy [2430],\$dummy [2431],\$dummy [2432],\$dummy [2433],
              \$dummy [2434],\$dummy [2435],\$dummy [2436],\$dummy [2437],
              \$dummy [2438],\$dummy [2439],\$dummy [2440],\$dummy [2441],
              \$dummy [2442],\$dummy [2443],\$dummy [2444],\$dummy [2445],
              \$dummy [2446],\$dummy [2447],\$dummy [2448],\$dummy [2449],
              \$dummy [2450],\$dummy [2451],\$dummy [2452],\$dummy [2453],
              \$dummy [2454],\$dummy [2455],\$dummy [2456],\$dummy [2457],
              \$dummy [2458],\$dummy [2459],\$dummy [2460],\$dummy [2461],
              \$dummy [2462],\$dummy [2463],\$dummy [2464],\$dummy [2465],
              \$dummy [2466],\$dummy [2467],\$dummy [2468],\$dummy [2469],
              \$dummy [2470],\$dummy [2471],\$dummy [2472],\$dummy [2473],
              \$dummy [2474],\$dummy [2475],\$dummy [2476],\$dummy [2477],
              \$dummy [2478],\$dummy [2479],\$dummy [2480],\$dummy [2481],
              \$dummy [2482],\$dummy [2483],\$dummy [2484],\$dummy [2485],
              \$dummy [2486],\$dummy [2487],\$dummy [2488],\$dummy [2489],
              \$dummy [2490],\$dummy [2491],\$dummy [2492],\$dummy [2493],
              \$dummy [2494],\$dummy [2495],\$dummy [2496],\$dummy [2497],
              \$dummy [2498],\$dummy [2499],\$dummy [2500],\$dummy [2501],
              \$dummy [2502],\$dummy [2503],\$dummy [2504],\$dummy [2505],
              \$dummy [2506],\$dummy [2507],\$dummy [2508],\$dummy [2509],
              \$dummy [2510],\$dummy [2511],\$dummy [2512],\$dummy [2513],
              \$dummy [2514],\$dummy [2515],\$dummy [2516],\$dummy [2517],
              \$dummy [2518],\$dummy [2519],\$dummy [2520],\$dummy [2521],
              \$dummy [2522],\$dummy [2523],\$dummy [2524],\$dummy [2525],
              \$dummy [2526],\$dummy [2527],\$dummy [2528],\$dummy [2529],
              \$dummy [2530],\$dummy [2531],\$dummy [2532],\$dummy [2533],
              \$dummy [2534],\$dummy [2535],\$dummy [2536],\$dummy [2537],
              \$dummy [2538],\$dummy [2539],\$dummy [2540],\$dummy [2541],
              \$dummy [2542],\$dummy [2543],\$dummy [2544],\$dummy [2545],
              \$dummy [2546],\$dummy [2547],\$dummy [2548],\$dummy [2549],
              \$dummy [2550],\$dummy [2551],\$dummy [2552],\$dummy [2553],
              \$dummy [2554],\$dummy [2555],\$dummy [2556],\$dummy [2557],
              \$dummy [2558],\$dummy [2559],\$dummy [2560],\$dummy [2561],
              \$dummy [2562],\$dummy [2563],\$dummy [2564],\$dummy [2565],
              \$dummy [2566],\$dummy [2567],\$dummy [2568],\$dummy [2569],
              \$dummy [2570],\$dummy [2571],\$dummy [2572],\$dummy [2573],
              \$dummy [2574],\$dummy [2575],\$dummy [2576],\$dummy [2577],
              \$dummy [2578],\$dummy [2579],\$dummy [2580],\$dummy [2581],
              \$dummy [2582],\$dummy [2583],\$dummy [2584],\$dummy [2585],
              \$dummy [2586],\$dummy [2587],\$dummy [2588],\$dummy [2589],
              \$dummy [2590],\$dummy [2591],\$dummy [2592],\$dummy [2593],
              \$dummy [2594],\$dummy [2595],\$dummy [2596],\$dummy [2597],
              \$dummy [2598],\$dummy [2599],\$dummy [2600],\$dummy [2601],
              \$dummy [2602],\$dummy [2603],\$dummy [2604],\$dummy [2605],
              \$dummy [2606],\$dummy [2607],\$dummy [2608],\$dummy [2609],
              \$dummy [2610],\$dummy [2611],\$dummy [2612],\$dummy [2613],
              \$dummy [2614],\$dummy [2615],\$dummy [2616],\$dummy [2617],
              \$dummy [2618],\$dummy [2619],\$dummy [2620],\$dummy [2621],
              \$dummy [2622],\$dummy [2623],\$dummy [2624],\$dummy [2625],
              \$dummy [2626],\$dummy [2627],\$dummy [2628],\$dummy [2629],
              \$dummy [2630],\$dummy [2631],\$dummy [2632],\$dummy [2633],
              \$dummy [2634],\$dummy [2635],\$dummy [2636],\$dummy [2637],
              \$dummy [2638],\$dummy [2639],\$dummy [2640],\$dummy [2641],
              \$dummy [2642],\$dummy [2643],\$dummy [2644],\$dummy [2645],
              \$dummy [2646],\$dummy [2647],\$dummy [2648],\$dummy [2649],
              \$dummy [2650],\$dummy [2651],\$dummy [2652],\$dummy [2653],
              \$dummy [2654],\$dummy [2655],\$dummy [2656],\$dummy [2657],
              \$dummy [2658],\$dummy [2659],\$dummy [2660],\$dummy [2661],
              \$dummy [2662],\$dummy [2663],\$dummy [2664],\$dummy [2665],
              \$dummy [2666],\$dummy [2667],\$dummy [2668],\$dummy [2669],
              \$dummy [2670],\$dummy [2671],\$dummy [2672],\$dummy [2673],
              \$dummy [2674],\$dummy [2675],\$dummy [2676],\$dummy [2677],
              \$dummy [2678],\$dummy [2679],\$dummy [2680],\$dummy [2681],
              \$dummy [2682],\$dummy [2683],\$dummy [2684],\$dummy [2685],
              \$dummy [2686],\$dummy [2687],\$dummy [2688],\$dummy [2689],
              \$dummy [2690],\$dummy [2691],\$dummy [2692],\$dummy [2693],
              \$dummy [2694],\$dummy [2695],\$dummy [2696],\$dummy [2697],
              \$dummy [2698],\$dummy [2699],\$dummy [2700],\$dummy [2701],
              \$dummy [2702],\$dummy [2703],\$dummy [2704],\$dummy [2705],
              \$dummy [2706],\$dummy [2707],\$dummy [2708],\$dummy [2709],
              \$dummy [2710],\$dummy [2711],\$dummy [2712],\$dummy [2713],
              \$dummy [2714],\$dummy [2715],\$dummy [2716],\$dummy [2717],
              \$dummy [2718],\$dummy [2719]}), .ImgCounterOuput ({
              ImgCounterOuput_2,ImgCounterOuput_1,ImgCounterOuput_0}), .ImgAddToDma (
              {AddressI_12,AddressI_11,AddressI_10,AddressI_9,AddressI_8,
              AddressI_7,AddressI_6,AddressI_5,AddressI_4,AddressI_3,AddressI_2,
              AddressI_1,AddressI_0}), .UpdatedAddress ({ImgAddRegIN_12,
              ImgAddRegIN_11,ImgAddRegIN_10,ImgAddRegIN_9,ImgAddRegIN_8,
              ImgAddRegIN_7,ImgAddRegIN_6,ImgAddRegIN_5,ImgAddRegIN_4,
              ImgAddRegIN_3,ImgAddRegIN_2,ImgAddRegIN_1,ImgAddRegIN_0}), .ImgIndic (
              {IndicatorI_0}), .ImgEn ({\$dummy [2720],\$dummy [2721],
              \$dummy [2722],\$dummy [2723],\$dummy [2724],\$dummy [2725]}), .dontTrust (
              DontRstIndicator)) ;
    Convolution Sconv (.current_state ({zero_11,zero_11,zero_11,zero_11,zero_11,
                zero_11,zero_11,nx9962,zero_11,zero_11,zero_11,zero_11,zero_11,
                zero_11,zero_11}), .CLK (nx10424), .RST (rst), .QImgStat (Q), .ACK (
                \$dummy [2726]), .LayerInfo ({LayerInfoOut_15,nx10500,zero_11,
                zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                zero_11,zero_11,zero_11,zero_11,zero_11}), .ImgAddress ({zero_11
                ,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11
                ,zero_11,zero_11,zero_11,zero_11}), .OutputImg0 ({OutputImg0_79,
                OutputImg0_78,OutputImg0_77,OutputImg0_76,OutputImg0_75,
                OutputImg0_74,OutputImg0_73,OutputImg0_72,OutputImg0_71,
                OutputImg0_70,OutputImg0_69,OutputImg0_68,OutputImg0_67,
                OutputImg0_66,OutputImg0_65,OutputImg0_64,OutputImg0_63,
                OutputImg0_62,OutputImg0_61,OutputImg0_60,OutputImg0_59,
                OutputImg0_58,OutputImg0_57,OutputImg0_56,OutputImg0_55,
                OutputImg0_54,OutputImg0_53,OutputImg0_52,OutputImg0_51,
                OutputImg0_50,OutputImg0_49,OutputImg0_48,OutputImg0_47,
                OutputImg0_46,OutputImg0_45,OutputImg0_44,OutputImg0_43,
                OutputImg0_42,OutputImg0_41,OutputImg0_40,OutputImg0_39,
                OutputImg0_38,OutputImg0_37,OutputImg0_36,OutputImg0_35,
                OutputImg0_34,OutputImg0_33,OutputImg0_32,OutputImg0_31,
                OutputImg0_30,OutputImg0_29,OutputImg0_28,OutputImg0_27,
                OutputImg0_26,OutputImg0_25,OutputImg0_24,OutputImg0_23,
                OutputImg0_22,OutputImg0_21,OutputImg0_20,OutputImg0_19,
                OutputImg0_18,OutputImg0_17,OutputImg0_16,OutputImg0_15,
                OutputImg0_14,OutputImg0_13,OutputImg0_12,OutputImg0_11,
                OutputImg0_10,OutputImg0_9,OutputImg0_8,OutputImg0_7,
                OutputImg0_6,OutputImg0_5,OutputImg0_4,OutputImg0_3,OutputImg0_2
                ,OutputImg0_1,OutputImg0_0}), .OutputImg1 ({OutputImg1_79,
                OutputImg1_78,OutputImg1_77,OutputImg1_76,OutputImg1_75,
                OutputImg1_74,OutputImg1_73,OutputImg1_72,OutputImg1_71,
                OutputImg1_70,OutputImg1_69,OutputImg1_68,OutputImg1_67,
                OutputImg1_66,OutputImg1_65,OutputImg1_64,OutputImg1_63,
                OutputImg1_62,OutputImg1_61,OutputImg1_60,OutputImg1_59,
                OutputImg1_58,OutputImg1_57,OutputImg1_56,OutputImg1_55,
                OutputImg1_54,OutputImg1_53,OutputImg1_52,OutputImg1_51,
                OutputImg1_50,OutputImg1_49,OutputImg1_48,OutputImg1_47,
                OutputImg1_46,OutputImg1_45,OutputImg1_44,OutputImg1_43,
                OutputImg1_42,OutputImg1_41,OutputImg1_40,OutputImg1_39,
                OutputImg1_38,OutputImg1_37,OutputImg1_36,OutputImg1_35,
                OutputImg1_34,OutputImg1_33,OutputImg1_32,OutputImg1_31,
                OutputImg1_30,OutputImg1_29,OutputImg1_28,OutputImg1_27,
                OutputImg1_26,OutputImg1_25,OutputImg1_24,OutputImg1_23,
                OutputImg1_22,OutputImg1_21,OutputImg1_20,OutputImg1_19,
                OutputImg1_18,OutputImg1_17,OutputImg1_16,OutputImg1_15,
                OutputImg1_14,OutputImg1_13,OutputImg1_12,OutputImg1_11,
                OutputImg1_10,OutputImg1_9,OutputImg1_8,OutputImg1_7,
                OutputImg1_6,OutputImg1_5,OutputImg1_4,OutputImg1_3,OutputImg1_2
                ,OutputImg1_1,OutputImg1_0}), .OutputImg2 ({OutputImg2_79,
                OutputImg2_78,OutputImg2_77,OutputImg2_76,OutputImg2_75,
                OutputImg2_74,OutputImg2_73,OutputImg2_72,OutputImg2_71,
                OutputImg2_70,OutputImg2_69,OutputImg2_68,OutputImg2_67,
                OutputImg2_66,OutputImg2_65,OutputImg2_64,OutputImg2_63,
                OutputImg2_62,OutputImg2_61,OutputImg2_60,OutputImg2_59,
                OutputImg2_58,OutputImg2_57,OutputImg2_56,OutputImg2_55,
                OutputImg2_54,OutputImg2_53,OutputImg2_52,OutputImg2_51,
                OutputImg2_50,OutputImg2_49,OutputImg2_48,OutputImg2_47,
                OutputImg2_46,OutputImg2_45,OutputImg2_44,OutputImg2_43,
                OutputImg2_42,OutputImg2_41,OutputImg2_40,OutputImg2_39,
                OutputImg2_38,OutputImg2_37,OutputImg2_36,OutputImg2_35,
                OutputImg2_34,OutputImg2_33,OutputImg2_32,OutputImg2_31,
                OutputImg2_30,OutputImg2_29,OutputImg2_28,OutputImg2_27,
                OutputImg2_26,OutputImg2_25,OutputImg2_24,OutputImg2_23,
                OutputImg2_22,OutputImg2_21,OutputImg2_20,OutputImg2_19,
                OutputImg2_18,OutputImg2_17,OutputImg2_16,OutputImg2_15,
                OutputImg2_14,OutputImg2_13,OutputImg2_12,OutputImg2_11,
                OutputImg2_10,OutputImg2_9,OutputImg2_8,OutputImg2_7,
                OutputImg2_6,OutputImg2_5,OutputImg2_4,OutputImg2_3,OutputImg2_2
                ,OutputImg2_1,OutputImg2_0}), .OutputImg3 ({OutputImg3_79,
                OutputImg3_78,OutputImg3_77,OutputImg3_76,OutputImg3_75,
                OutputImg3_74,OutputImg3_73,OutputImg3_72,OutputImg3_71,
                OutputImg3_70,OutputImg3_69,OutputImg3_68,OutputImg3_67,
                OutputImg3_66,OutputImg3_65,OutputImg3_64,OutputImg3_63,
                OutputImg3_62,OutputImg3_61,OutputImg3_60,OutputImg3_59,
                OutputImg3_58,OutputImg3_57,OutputImg3_56,OutputImg3_55,
                OutputImg3_54,OutputImg3_53,OutputImg3_52,OutputImg3_51,
                OutputImg3_50,OutputImg3_49,OutputImg3_48,OutputImg3_47,
                OutputImg3_46,OutputImg3_45,OutputImg3_44,OutputImg3_43,
                OutputImg3_42,OutputImg3_41,OutputImg3_40,OutputImg3_39,
                OutputImg3_38,OutputImg3_37,OutputImg3_36,OutputImg3_35,
                OutputImg3_34,OutputImg3_33,OutputImg3_32,OutputImg3_31,
                OutputImg3_30,OutputImg3_29,OutputImg3_28,OutputImg3_27,
                OutputImg3_26,OutputImg3_25,OutputImg3_24,OutputImg3_23,
                OutputImg3_22,OutputImg3_21,OutputImg3_20,OutputImg3_19,
                OutputImg3_18,OutputImg3_17,OutputImg3_16,OutputImg3_15,
                OutputImg3_14,OutputImg3_13,OutputImg3_12,OutputImg3_11,
                OutputImg3_10,OutputImg3_9,OutputImg3_8,OutputImg3_7,
                OutputImg3_6,OutputImg3_5,OutputImg3_4,OutputImg3_3,OutputImg3_2
                ,OutputImg3_1,OutputImg3_0}), .OutputImg4 ({OutputImg4_79,
                OutputImg4_78,OutputImg4_77,OutputImg4_76,OutputImg4_75,
                OutputImg4_74,OutputImg4_73,OutputImg4_72,OutputImg4_71,
                OutputImg4_70,OutputImg4_69,OutputImg4_68,OutputImg4_67,
                OutputImg4_66,OutputImg4_65,OutputImg4_64,OutputImg4_63,
                OutputImg4_62,OutputImg4_61,OutputImg4_60,OutputImg4_59,
                OutputImg4_58,OutputImg4_57,OutputImg4_56,OutputImg4_55,
                OutputImg4_54,OutputImg4_53,OutputImg4_52,OutputImg4_51,
                OutputImg4_50,OutputImg4_49,OutputImg4_48,OutputImg4_47,
                OutputImg4_46,OutputImg4_45,OutputImg4_44,OutputImg4_43,
                OutputImg4_42,OutputImg4_41,OutputImg4_40,OutputImg4_39,
                OutputImg4_38,OutputImg4_37,OutputImg4_36,OutputImg4_35,
                OutputImg4_34,OutputImg4_33,OutputImg4_32,OutputImg4_31,
                OutputImg4_30,OutputImg4_29,OutputImg4_28,OutputImg4_27,
                OutputImg4_26,OutputImg4_25,OutputImg4_24,OutputImg4_23,
                OutputImg4_22,OutputImg4_21,OutputImg4_20,OutputImg4_19,
                OutputImg4_18,OutputImg4_17,OutputImg4_16,OutputImg4_15,
                OutputImg4_14,OutputImg4_13,OutputImg4_12,OutputImg4_11,
                OutputImg4_10,OutputImg4_9,OutputImg4_8,OutputImg4_7,
                OutputImg4_6,OutputImg4_5,OutputImg4_4,OutputImg4_3,OutputImg4_2
                ,OutputImg4_1,OutputImg4_0}), .outFilter0 ({Filter1_399,
                Filter1_398,Filter1_397,Filter1_396,Filter1_395,Filter1_394,
                Filter1_393,Filter1_392,Filter1_391,Filter1_390,Filter1_389,
                Filter1_388,Filter1_387,Filter1_386,Filter1_385,Filter1_384,
                Filter1_383,Filter1_382,Filter1_381,Filter1_380,Filter1_379,
                Filter1_378,Filter1_377,Filter1_376,Filter1_375,Filter1_374,
                Filter1_373,Filter1_372,Filter1_371,Filter1_370,Filter1_369,
                Filter1_368,Filter1_367,Filter1_366,Filter1_365,Filter1_364,
                Filter1_363,Filter1_362,Filter1_361,Filter1_360,Filter1_359,
                Filter1_358,Filter1_357,Filter1_356,Filter1_355,Filter1_354,
                Filter1_353,Filter1_352,Filter1_351,Filter1_350,Filter1_349,
                Filter1_348,Filter1_347,Filter1_346,Filter1_345,Filter1_344,
                Filter1_343,Filter1_342,Filter1_341,Filter1_340,Filter1_339,
                Filter1_338,Filter1_337,Filter1_336,Filter1_335,Filter1_334,
                Filter1_333,Filter1_332,Filter1_331,Filter1_330,Filter1_329,
                Filter1_328,Filter1_327,Filter1_326,Filter1_325,Filter1_324,
                Filter1_323,Filter1_322,Filter1_321,Filter1_320,Filter1_319,
                Filter1_318,Filter1_317,Filter1_316,Filter1_315,Filter1_314,
                Filter1_313,Filter1_312,Filter1_311,Filter1_310,Filter1_309,
                Filter1_308,Filter1_307,Filter1_306,Filter1_305,Filter1_304,
                Filter1_303,Filter1_302,Filter1_301,Filter1_300,Filter1_299,
                Filter1_298,Filter1_297,Filter1_296,Filter1_295,Filter1_294,
                Filter1_293,Filter1_292,Filter1_291,Filter1_290,Filter1_289,
                Filter1_288,Filter1_287,Filter1_286,Filter1_285,Filter1_284,
                Filter1_283,Filter1_282,Filter1_281,Filter1_280,Filter1_279,
                Filter1_278,Filter1_277,Filter1_276,Filter1_275,Filter1_274,
                Filter1_273,Filter1_272,Filter1_271,Filter1_270,Filter1_269,
                Filter1_268,Filter1_267,Filter1_266,Filter1_265,Filter1_264,
                Filter1_263,Filter1_262,Filter1_261,Filter1_260,Filter1_259,
                Filter1_258,Filter1_257,Filter1_256,Filter1_255,Filter1_254,
                Filter1_253,Filter1_252,Filter1_251,Filter1_250,Filter1_249,
                Filter1_248,Filter1_247,Filter1_246,Filter1_245,Filter1_244,
                Filter1_243,Filter1_242,Filter1_241,Filter1_240,Filter1_239,
                Filter1_238,Filter1_237,Filter1_236,Filter1_235,Filter1_234,
                Filter1_233,Filter1_232,Filter1_231,Filter1_230,Filter1_229,
                Filter1_228,Filter1_227,Filter1_226,Filter1_225,Filter1_224,
                Filter1_223,Filter1_222,Filter1_221,Filter1_220,Filter1_219,
                Filter1_218,Filter1_217,Filter1_216,Filter1_215,Filter1_214,
                Filter1_213,Filter1_212,Filter1_211,Filter1_210,Filter1_209,
                Filter1_208,Filter1_207,Filter1_206,Filter1_205,Filter1_204,
                Filter1_203,Filter1_202,Filter1_201,Filter1_200,Filter1_199,
                Filter1_198,Filter1_197,Filter1_196,Filter1_195,Filter1_194,
                Filter1_193,Filter1_192,Filter1_191,Filter1_190,Filter1_189,
                Filter1_188,Filter1_187,Filter1_186,Filter1_185,Filter1_184,
                Filter1_183,Filter1_182,Filter1_181,Filter1_180,Filter1_179,
                Filter1_178,Filter1_177,Filter1_176,Filter1_175,Filter1_174,
                Filter1_173,Filter1_172,Filter1_171,Filter1_170,Filter1_169,
                Filter1_168,Filter1_167,Filter1_166,Filter1_165,Filter1_164,
                Filter1_163,Filter1_162,Filter1_161,Filter1_160,Filter1_159,
                Filter1_158,Filter1_157,Filter1_156,Filter1_155,Filter1_154,
                Filter1_153,Filter1_152,Filter1_151,Filter1_150,Filter1_149,
                Filter1_148,Filter1_147,Filter1_146,Filter1_145,Filter1_144,
                Filter1_143,Filter1_142,Filter1_141,Filter1_140,Filter1_139,
                Filter1_138,Filter1_137,Filter1_136,Filter1_135,Filter1_134,
                Filter1_133,Filter1_132,Filter1_131,Filter1_130,Filter1_129,
                Filter1_128,Filter1_127,Filter1_126,Filter1_125,Filter1_124,
                Filter1_123,Filter1_122,Filter1_121,Filter1_120,Filter1_119,
                Filter1_118,Filter1_117,Filter1_116,Filter1_115,Filter1_114,
                Filter1_113,Filter1_112,Filter1_111,Filter1_110,Filter1_109,
                Filter1_108,Filter1_107,Filter1_106,Filter1_105,Filter1_104,
                Filter1_103,Filter1_102,Filter1_101,Filter1_100,Filter1_99,
                Filter1_98,Filter1_97,Filter1_96,Filter1_95,Filter1_94,
                Filter1_93,Filter1_92,Filter1_91,Filter1_90,Filter1_89,
                Filter1_88,Filter1_87,Filter1_86,Filter1_85,Filter1_84,
                Filter1_83,Filter1_82,Filter1_81,Filter1_80,Filter1_79,
                Filter1_78,Filter1_77,Filter1_76,Filter1_75,Filter1_74,
                Filter1_73,Filter1_72,Filter1_71,Filter1_70,Filter1_69,
                Filter1_68,Filter1_67,Filter1_66,Filter1_65,Filter1_64,
                Filter1_63,Filter1_62,Filter1_61,Filter1_60,Filter1_59,
                Filter1_58,Filter1_57,Filter1_56,Filter1_55,Filter1_54,
                Filter1_53,Filter1_52,Filter1_51,Filter1_50,Filter1_49,
                Filter1_48,Filter1_47,Filter1_46,Filter1_45,Filter1_44,
                Filter1_43,Filter1_42,Filter1_41,Filter1_40,Filter1_39,
                Filter1_38,Filter1_37,Filter1_36,Filter1_35,Filter1_34,
                Filter1_33,Filter1_32,Filter1_31,Filter1_30,Filter1_29,
                Filter1_28,Filter1_27,Filter1_26,Filter1_25,Filter1_24,
                Filter1_23,Filter1_22,Filter1_21,Filter1_20,Filter1_19,
                Filter1_18,Filter1_17,Filter1_16,Filter1_15,Filter1_14,
                Filter1_13,Filter1_12,Filter1_11,Filter1_10,Filter1_9,Filter1_8,
                Filter1_7,Filter1_6,Filter1_5,Filter1_4,Filter1_3,Filter1_2,
                Filter1_1,Filter1_0}), .outFilter1 ({Filter2_399,Filter2_398,
                Filter2_397,Filter2_396,Filter2_395,Filter2_394,Filter2_393,
                Filter2_392,Filter2_391,Filter2_390,Filter2_389,Filter2_388,
                Filter2_387,Filter2_386,Filter2_385,Filter2_384,Filter2_383,
                Filter2_382,Filter2_381,Filter2_380,Filter2_379,Filter2_378,
                Filter2_377,Filter2_376,Filter2_375,Filter2_374,Filter2_373,
                Filter2_372,Filter2_371,Filter2_370,Filter2_369,Filter2_368,
                Filter2_367,Filter2_366,Filter2_365,Filter2_364,Filter2_363,
                Filter2_362,Filter2_361,Filter2_360,Filter2_359,Filter2_358,
                Filter2_357,Filter2_356,Filter2_355,Filter2_354,Filter2_353,
                Filter2_352,Filter2_351,Filter2_350,Filter2_349,Filter2_348,
                Filter2_347,Filter2_346,Filter2_345,Filter2_344,Filter2_343,
                Filter2_342,Filter2_341,Filter2_340,Filter2_339,Filter2_338,
                Filter2_337,Filter2_336,Filter2_335,Filter2_334,Filter2_333,
                Filter2_332,Filter2_331,Filter2_330,Filter2_329,Filter2_328,
                Filter2_327,Filter2_326,Filter2_325,Filter2_324,Filter2_323,
                Filter2_322,Filter2_321,Filter2_320,Filter2_319,Filter2_318,
                Filter2_317,Filter2_316,Filter2_315,Filter2_314,Filter2_313,
                Filter2_312,Filter2_311,Filter2_310,Filter2_309,Filter2_308,
                Filter2_307,Filter2_306,Filter2_305,Filter2_304,Filter2_303,
                Filter2_302,Filter2_301,Filter2_300,Filter2_299,Filter2_298,
                Filter2_297,Filter2_296,Filter2_295,Filter2_294,Filter2_293,
                Filter2_292,Filter2_291,Filter2_290,Filter2_289,Filter2_288,
                Filter2_287,Filter2_286,Filter2_285,Filter2_284,Filter2_283,
                Filter2_282,Filter2_281,Filter2_280,Filter2_279,Filter2_278,
                Filter2_277,Filter2_276,Filter2_275,Filter2_274,Filter2_273,
                Filter2_272,Filter2_271,Filter2_270,Filter2_269,Filter2_268,
                Filter2_267,Filter2_266,Filter2_265,Filter2_264,Filter2_263,
                Filter2_262,Filter2_261,Filter2_260,Filter2_259,Filter2_258,
                Filter2_257,Filter2_256,Filter2_255,Filter2_254,Filter2_253,
                Filter2_252,Filter2_251,Filter2_250,Filter2_249,Filter2_248,
                Filter2_247,Filter2_246,Filter2_245,Filter2_244,Filter2_243,
                Filter2_242,Filter2_241,Filter2_240,Filter2_239,Filter2_238,
                Filter2_237,Filter2_236,Filter2_235,Filter2_234,Filter2_233,
                Filter2_232,Filter2_231,Filter2_230,Filter2_229,Filter2_228,
                Filter2_227,Filter2_226,Filter2_225,Filter2_224,Filter2_223,
                Filter2_222,Filter2_221,Filter2_220,Filter2_219,Filter2_218,
                Filter2_217,Filter2_216,Filter2_215,Filter2_214,Filter2_213,
                Filter2_212,Filter2_211,Filter2_210,Filter2_209,Filter2_208,
                Filter2_207,Filter2_206,Filter2_205,Filter2_204,Filter2_203,
                Filter2_202,Filter2_201,Filter2_200,Filter2_199,Filter2_198,
                Filter2_197,Filter2_196,Filter2_195,Filter2_194,Filter2_193,
                Filter2_192,Filter2_191,Filter2_190,Filter2_189,Filter2_188,
                Filter2_187,Filter2_186,Filter2_185,Filter2_184,Filter2_183,
                Filter2_182,Filter2_181,Filter2_180,Filter2_179,Filter2_178,
                Filter2_177,Filter2_176,Filter2_175,Filter2_174,Filter2_173,
                Filter2_172,Filter2_171,Filter2_170,Filter2_169,Filter2_168,
                Filter2_167,Filter2_166,Filter2_165,Filter2_164,Filter2_163,
                Filter2_162,Filter2_161,Filter2_160,Filter2_159,Filter2_158,
                Filter2_157,Filter2_156,Filter2_155,Filter2_154,Filter2_153,
                Filter2_152,Filter2_151,Filter2_150,Filter2_149,Filter2_148,
                Filter2_147,Filter2_146,Filter2_145,Filter2_144,Filter2_143,
                Filter2_142,Filter2_141,Filter2_140,Filter2_139,Filter2_138,
                Filter2_137,Filter2_136,Filter2_135,Filter2_134,Filter2_133,
                Filter2_132,Filter2_131,Filter2_130,Filter2_129,Filter2_128,
                Filter2_127,Filter2_126,Filter2_125,Filter2_124,Filter2_123,
                Filter2_122,Filter2_121,Filter2_120,Filter2_119,Filter2_118,
                Filter2_117,Filter2_116,Filter2_115,Filter2_114,Filter2_113,
                Filter2_112,Filter2_111,Filter2_110,Filter2_109,Filter2_108,
                Filter2_107,Filter2_106,Filter2_105,Filter2_104,Filter2_103,
                Filter2_102,Filter2_101,Filter2_100,Filter2_99,Filter2_98,
                Filter2_97,Filter2_96,Filter2_95,Filter2_94,Filter2_93,
                Filter2_92,Filter2_91,Filter2_90,Filter2_89,Filter2_88,
                Filter2_87,Filter2_86,Filter2_85,Filter2_84,Filter2_83,
                Filter2_82,Filter2_81,Filter2_80,Filter2_79,Filter2_78,
                Filter2_77,Filter2_76,Filter2_75,Filter2_74,Filter2_73,
                Filter2_72,Filter2_71,Filter2_70,Filter2_69,Filter2_68,
                Filter2_67,Filter2_66,Filter2_65,Filter2_64,Filter2_63,
                Filter2_62,Filter2_61,Filter2_60,Filter2_59,Filter2_58,
                Filter2_57,Filter2_56,Filter2_55,Filter2_54,Filter2_53,
                Filter2_52,Filter2_51,Filter2_50,Filter2_49,Filter2_48,
                Filter2_47,Filter2_46,Filter2_45,Filter2_44,Filter2_43,
                Filter2_42,Filter2_41,Filter2_40,Filter2_39,Filter2_38,
                Filter2_37,Filter2_36,Filter2_35,Filter2_34,Filter2_33,
                Filter2_32,Filter2_31,Filter2_30,Filter2_29,Filter2_28,
                Filter2_27,Filter2_26,Filter2_25,Filter2_24,Filter2_23,
                Filter2_22,Filter2_21,Filter2_20,Filter2_19,Filter2_18,
                Filter2_17,Filter2_16,Filter2_15,Filter2_14,Filter2_13,
                Filter2_12,Filter2_11,Filter2_10,Filter2_9,Filter2_8,Filter2_7,
                Filter2_6,Filter2_5,Filter2_4,Filter2_3,Filter2_2,Filter2_1,
                Filter2_0}), .ConvOuput ({ConvOuput_15,ConvOuput_14,ConvOuput_13
                ,ConvOuput_12,ConvOuput_11,ConvOuput_10,ConvOuput_9,ConvOuput_8,
                ConvOuput_7,ConvOuput_6,ConvOuput_5,ConvOuput_4,ConvOuput_3,
                ConvOuput_2,ConvOuput_1,ConvOuput_0})) ;
    saveState Ssave (.DMAOutput ({nx10314,nx10318,nx10322,nx10326,nx10330,
              nx10334,nx10338,nx10342,nx10346,nx10350,nx10354,nx10358,nx10362,
              nx10366,nx10370,nx10374}), .RegisterOutput ({nx10396,ConvOuput_14,
              ConvOuput_13,ConvOuput_12,ConvOuput_11,ConvOuput_10,ConvOuput_9,
              ConvOuput_8,ConvOuput_7,ConvOuput_6,ConvOuput_5,ConvOuput_4,
              ConvOuput_3,ConvOuput_2,ConvOuput_1,ConvOuput_0}), .bias1 ({
              Bias0_15,Bias0_14,Bias0_13,Bias0_12,Bias0_11,Bias0_10,Bias0_9,
              Bias0_8,Bias0_7,Bias0_6,Bias0_5,Bias0_4,Bias0_3,Bias0_2,Bias0_1,
              Bias0_0}), .bias2 ({Bias1_15,Bias1_14,Bias1_13,Bias1_12,Bias1_11,
              Bias1_10,Bias1_9,Bias1_8,Bias1_7,Bias1_6,Bias1_5,Bias1_4,Bias1_3,
              Bias1_2,Bias1_1,Bias1_0}), .bias3 ({Bias2_15,Bias2_14,Bias2_13,
              Bias2_12,Bias2_11,Bias2_10,Bias2_9,Bias2_8,Bias2_7,Bias2_6,Bias2_5
              ,Bias2_4,Bias2_3,Bias2_2,Bias2_1,Bias2_0}), .bias4 ({Bias3_15,
              Bias3_14,Bias3_13,Bias3_12,Bias3_11,Bias3_10,Bias3_9,Bias3_8,
              Bias3_7,Bias3_6,Bias3_5,Bias3_4,Bias3_3,Bias3_2,Bias3_1,Bias3_0})
              , .bias5 ({Bias4_15,Bias4_14,Bias4_13,Bias4_12,Bias4_11,Bias4_10,
              Bias4_9,Bias4_8,Bias4_7,Bias4_6,Bias4_5,Bias4_4,Bias4_3,Bias4_2,
              Bias4_1,Bias4_0}), .bias6 ({Bias5_15,Bias5_14,Bias5_13,Bias5_12,
              Bias5_11,Bias5_10,Bias5_9,Bias5_8,Bias5_7,Bias5_6,Bias5_5,Bias5_4,
              Bias5_3,Bias5_2,Bias5_1,Bias5_0}), .bias7 ({Bias6_15,Bias6_14,
              Bias6_13,Bias6_12,Bias6_11,Bias6_10,Bias6_9,Bias6_8,Bias6_7,
              Bias6_6,Bias6_5,Bias6_4,Bias6_3,Bias6_2,Bias6_1,Bias6_0}), .bias8 (
              {Bias7_15,Bias7_14,Bias7_13,Bias7_12,Bias7_11,Bias7_10,Bias7_9,
              Bias7_8,Bias7_7,Bias7_6,Bias7_5,Bias7_4,Bias7_3,Bias7_2,Bias7_1,
              Bias7_0}), .Depth ({nx10406,nx10408,nx10410,nx10412}), .NumberOfFiltersCounter (
              {nx10398,nx10400,nx10402,nx10404}), .rst (rst), .stateinput ({
              zero_11,nx9950,nx9954,zero_11,current_state_10,nx9958,
              current_state_8,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
              zero_11,zero_11}), .clk (nx10424), .outputCounterToDma ({
              AddressI_12,AddressI_11,AddressI_10,AddressI_9,AddressI_8,
              AddressI_7,AddressI_6,AddressI_5,AddressI_4,AddressI_3,AddressI_2,
              AddressI_1,AddressI_0}), .RealOutputCounter ({RealOutputCounter_12
              ,RealOutputCounter_11,RealOutputCounter_10,RealOutputCounter_9,
              RealOutputCounter_8,RealOutputCounter_7,RealOutputCounter_6,
              RealOutputCounter_5,RealOutputCounter_4,RealOutputCounter_3,
              RealOutputCounter_2,RealOutputCounter_1,RealOutputCounter_0}), .\output  (
              {DataIIn_15,DataIIn_14,DataIIn_13,DataIIn_12,DataIIn_11,DataIIn_10
              ,DataIIn_9,DataIIn_8,DataIIn_7,DataIIn_6,DataIIn_5,DataIIn_4,
              DataIIn_3,DataIIn_2,DataIIn_1,DataIIn_0}), .ShiftLeftCounterOutput (
              {ShiftLeftCounterOutput_4,ShiftLeftCounterOutput_3,
              ShiftLeftCounterOutput_2,ShiftLeftCounterOutput_1,
              ShiftLeftCounterOutput_0}), .ShiftCounterRst (ShiftCounterRst), .AddresCounterLoad (
              {OutputCounterLoad_12,OutputCounterLoad_11,OutputCounterLoad_10,
              OutputCounterLoad_9,OutputCounterLoad_8,OutputCounterLoad_7,
              OutputCounterLoad_6,OutputCounterLoad_5,OutputCounterLoad_4,
              OutputCounterLoad_3,OutputCounterLoad_2,OutputCounterLoad_1,
              OutputCounterLoad_0}), .X (X), .Y (Y)) ;
    ImageState Istate (.current_state ({zero_11,nx9950,nx9954,current_state_11,
               zero_11,nx9958,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
               zero_11,zero_11,zero_11}), .WSquared ({WidthSquareOut_9,
               WidthSquareOut_8,WidthSquareOut_7,WidthSquareOut_6,
               WidthSquareOut_5,WidthSquareOut_4,WidthSquareOut_3,
               WidthSquareOut_2,WidthSquareOut_1,WidthSquareOut_0}), .AddresCounterIN (
               {RealOutputCounter_12,RealOutputCounter_11,RealOutputCounter_10,
               RealOutputCounter_9,RealOutputCounter_8,RealOutputCounter_7,
               RealOutputCounter_6,RealOutputCounter_5,RealOutputCounter_4,
               RealOutputCounter_3,RealOutputCounter_2,RealOutputCounter_1,
               RealOutputCounter_0}), .AddresCounterLoad ({OutputCounterLoad_12,
               OutputCounterLoad_11,OutputCounterLoad_10,OutputCounterLoad_9,
               OutputCounterLoad_8,OutputCounterLoad_7,OutputCounterLoad_6,
               OutputCounterLoad_5,OutputCounterLoad_4,OutputCounterLoad_3,
               OutputCounterLoad_2,OutputCounterLoad_1,OutputCounterLoad_0}), .NoOfShiftsCounter (
               {ShiftLeftCounterOutput_4,ShiftLeftCounterOutput_3,
               ShiftLeftCounterOutput_2,ShiftLeftCounterOutput_1,
               ShiftLeftCounterOutput_0}), .LayerInfoIn ({zero_11,zero_11,
               zero_11,zero_11,zero_11,zero_11,zero_11,nx10378,nx10382,nx10386,
               nx10388,nx10392,LayerInfoOut_3,LayerInfoOut_2,LayerInfoOut_1,
               LayerInfoOut_0}), .CLK (nx10426), .RST (rst), .Q (Q), .NumOfFilters (
               {NumOfFilters_3,NumOfFilters_2,NumOfFilters_1,NumOfFilters_0}), .NumOfHeight (
               {NumOfHeight_4,NumOfHeight_3,NumOfHeight_2,NumOfHeight_1,
               NumOfHeight_0}), .X1 (X), .Y1 (Y), .K1 (K)) ;
    StateChecks ChState (.current_state ({zero_11,nx9950,nx9956,zero_11,zero_11,
                zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                zero_11,zero_11}), .noOfLayers ({zero_11,zero_11,zero_11,zero_11
                ,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11
                ,zero_11,zero_11,NoOfLayers_1,NoOfLayers_0}), .LayerInfo ({
                zero_11,zero_11,zero_11,LayerInfoOut_12,LayerInfoOut_11,
                LayerInfoOut_10,LayerInfoOut_9,zero_11,zero_11,zero_11,zero_11,
                zero_11,zero_11,zero_11,zero_11,zero_11}), .CLK (zero_11), .RST (
                rst), .L (L), .D (D), .CNDoutput ({CNDepthoutput_3,
                CNDepthoutput_2,CNDepthoutput_1,CNDepthoutput_0}), .CNLoutput ({
                \$dummy [2727],\$dummy [2728]})) ;
    outWidthState Owidth (.currentState ({zero_11,nx9950,zero_11,zero_11,zero_11
                  ,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,zero_11,
                  zero_11,zero_11,zero_11}), .infoReg ({zero_11,zero_11,zero_11,
                  zero_11,zero_11,zero_11,zero_11,nx10378,nx10382,nx10386,
                  nx10388,nx10392,zero_11,zero_11,zero_11,zero_11}), .address ({
                  AddressI_12,AddressI_11,AddressI_10,AddressI_9,AddressI_8,
                  AddressI_7,AddressI_6,AddressI_5,AddressI_4,AddressI_3,
                  AddressI_2,AddressI_1,AddressI_0}), .outWidth ({DataIIn_15,
                  DataIIn_14,DataIIn_13,DataIIn_12,DataIIn_11,DataIIn_10,
                  DataIIn_9,DataIIn_8,DataIIn_7,DataIIn_6,DataIIn_5,DataIIn_4,
                  DataIIn_3,DataIIn_2,DataIIn_1,DataIIn_0})) ;
    fake_vcc ix9649 (.Y (PWR)) ;
    fake_gnd ix9647 (.Y (zero_11)) ;
    or02 ix399 (.Y (ramSelector), .A0 (current_state_8), .A1 (nx9950)) ;
    dffr reg_current_state_8 (.Q (current_state_8), .QB (\$dummy [2729]), .D (
         next_state_8), .CLK (nx10430), .R (rst)) ;
    latch lat_next_state_8 (.Q (next_state_8), .D (nx9962), .CLK (nx10434)) ;
    dffr reg_current_state_7 (.Q (\$dummy [2730]), .QB (nx9870), .D (
         next_state_7), .CLK (nx10428), .R (rst)) ;
    latch lat_next_state_7 (.Q (next_state_7), .D (nx154), .CLK (nx10434)) ;
    nand02 ix155 (.Y (nx154), .A0 (nx9760), .A1 (nx9814)) ;
    aoi22 ix9761 (.Y (nx9760), .A0 (K), .A1 (current_state_11), .B0 (X), .B1 (
          nx9960)) ;
    dffr reg_current_state_11 (.Q (current_state_11), .QB (\$dummy [2731]), .D (
         next_state_11), .CLK (nx10426), .R (rst)) ;
    latch lat_next_state_11 (.Q (next_state_11), .D (nx256), .CLK (nx10432)) ;
    nor03_2x ix257 (.Y (nx256), .A0 (nx9765), .A1 (Y), .A2 (nx9768)) ;
    nand04 ix9766 (.Y (nx9765), .A0 (ShiftLeftCounterOutput_2), .A1 (
           ShiftLeftCounterOutput_4), .A2 (ShiftLeftCounterOutput_3), .A3 (nx18)
           ) ;
    nor02_2x ix19 (.Y (nx18), .A0 (ShiftLeftCounterOutput_1), .A1 (
             ShiftLeftCounterOutput_0)) ;
    latch lat_next_state_10 (.Q (next_state_10), .D (nx240), .CLK (nx10432)) ;
    dffr reg_current_state_9 (.Q (current_state_9), .QB (\$dummy [2732]), .D (
         next_state_9), .CLK (nx10426), .R (rst)) ;
    latch lat_next_state_9 (.Q (next_state_9), .D (nx224), .CLK (nx10432)) ;
    and02 ix225 (.Y (nx224), .A0 (next_state_dup_124), .A1 (current_state_8)) ;
    dff reg_next_state_dup_124 (.Q (next_state_dup_124), .QB (\$dummy [2733]), .D (
        nx9738), .CLK (nx10028)) ;
    or02 ix9739 (.Y (nx9738), .A0 (next_state_dup_124), .A1 (WriteI)) ;
    nand02 ix217 (.Y (WriteI), .A0 (nx9780), .A1 (nx9792)) ;
    oai21 ix9781 (.Y (nx9780), .A0 (nx210), .A1 (SaveAckLatch), .B0 (
          current_state_8)) ;
    nor04 ix211 (.Y (nx210), .A0 (nx10406), .A1 (nx10408), .A2 (nx10410), .A3 (
          nx10412)) ;
    dffr ix9064 (.Q (nx9063), .QB (\$dummy [2734]), .D (PWR), .CLK (nx10436), .R (
         nx180)) ;
    nand02 ix9786 (.Y (NOT_nx0), .A0 (start), .A1 (cl)) ;
    nand02 ix181 (.Y (nx180), .A0 (current_state_8), .A1 (nx10026)) ;
    latch lat_next_state_13 (.Q (next_state_13), .D (nx9711), .CLK (nx10432)) ;
    aoi21 ix289 (.Y (nx9711), .A0 (L), .A1 (D), .B0 (nx9796)) ;
    dffr reg_current_state_12 (.Q (\$dummy [2735]), .QB (nx9796), .D (
         next_state_12), .CLK (nx10426), .R (rst)) ;
    latch lat_next_state_12 (.Q (next_state_12), .D (nx270), .CLK (nx10432)) ;
    nor02ii ix271 (.Y (nx270), .A0 (K), .A1 (current_state_11)) ;
    dffr reg_current_state_14 (.Q (done), .QB (\$dummy [2736]), .D (
         next_state_14), .CLK (nx10420), .R (rst)) ;
    latch lat_next_state_14 (.Q (next_state_14), .D (nx300), .CLK (nx10432)) ;
    dff reg_next_state_dup_134 (.Q (next_state_dup_134), .QB (\$dummy [2737]), .D (
        NOT_L), .CLK (nx10028)) ;
    inv01 ix9806 (.Y (NOT_L), .A (L)) ;
    dffr reg_current_state_13 (.Q (\$dummy [2738]), .QB (nx9792), .D (
         next_state_13), .CLK (nx10418), .R (rst)) ;
    dffr reg_current_state_10 (.Q (current_state_10), .QB (nx9768), .D (
         next_state_10), .CLK (nx10426), .R (rst)) ;
    aoi32 ix9815 (.Y (nx9814), .A0 (nx20), .A1 (Y), .A2 (current_state_10), .B0 (
          next_state_dup_96), .B1 (nx142)) ;
    dff reg_next_state_dup_96 (.Q (next_state_dup_96), .QB (\$dummy [2739]), .D (
        nx9718), .CLK (nx10028)) ;
    or02 ix9719 (.Y (nx9718), .A0 (next_state_dup_96), .A1 (nx48)) ;
    aoi21 ix49 (.Y (nx48), .A0 (nx9822), .A1 (nx9826), .B0 (ImgCounterOuput_0)
          ) ;
    nand03 ix9823 (.Y (nx9822), .A0 (nx10500), .A1 (ImgCounterOuput_2), .A2 (
           nx9824)) ;
    inv01 ix9825 (.Y (nx9824), .A (ImgCounterOuput_1)) ;
    or03 ix9827 (.Y (nx9826), .A0 (nx10502), .A1 (ImgCounterOuput_2), .A2 (
         nx9824)) ;
    dffr reg_current_state_3 (.Q (current_state_3), .QB (\$dummy [2740]), .D (
         next_state_3), .CLK (nx10428), .R (rst)) ;
    latch lat_next_state_3 (.Q (next_state_3), .D (nx130), .CLK (nx10434)) ;
    nand02 ix131 (.Y (nx130), .A0 (nx9833), .A1 (nx9835)) ;
    nand04 ix9834 (.Y (nx9833), .A0 (nx9954), .A1 (L), .A2 (D), .A3 (
           LayerInfoOut_15)) ;
    dffr reg_current_state_2 (.Q (current_state_2), .QB (nx9835), .D (
         next_state_2), .CLK (nx10428), .R (rst)) ;
    latch lat_next_state_2 (.Q (next_state_2), .D (nx112), .CLK (nx10434)) ;
    dff reg_next_state_dup_26 (.Q (next_state_dup_26), .QB (\$dummy [2741]), .D (
        nx9728), .CLK (nx10436)) ;
    mux21_ni ix9729 (.Y (nx9728), .A0 (next_state_dup_26), .A1 (nx10304), .S0 (
             nx10308)) ;
    dffr reg_current_state_1 (.Q (\$dummy [2742]), .QB (nx9849), .D (
         next_state_1), .CLK (nx10428), .R (rst)) ;
    latch lat_next_state_1 (.Q (next_state_1), .D (nx100), .CLK (nx10432)) ;
    ao21 ix101 (.Y (nx100), .A0 (next_state_dup_147), .A1 (nx9950), .B0 (
         current_state_0)) ;
    dff reg_next_state_dup_147 (.Q (next_state_dup_147), .QB (\$dummy [2743]), .D (
        L), .CLK (nx10028)) ;
    dffs_ni reg_current_state_0 (.Q (current_state_0), .QB (\$dummy [2744]), .D (
            zero_11), .CLK (nx10426), .S (rst)) ;
    dffr reg_current_state_6 (.Q (current_state_6), .QB (\$dummy [2745]), .D (
         next_state_6), .CLK (nx10428), .R (rst)) ;
    latch lat_next_state_6 (.Q (next_state_6), .D (nx66), .CLK (nx10434)) ;
    nand02 ix67 (.Y (nx66), .A0 (nx9854), .A1 (nx9858)) ;
    nand04 ix9855 (.Y (nx9854), .A0 (nx9954), .A1 (L), .A2 (D), .A3 (nx9856)) ;
    inv01 ix9857 (.Y (nx9856), .A (LayerInfoOut_15)) ;
    dffr reg_current_state_5 (.Q (current_state_5), .QB (nx9858), .D (
         next_state_5), .CLK (nx10428), .R (rst)) ;
    latch lat_next_state_5 (.Q (next_state_5), .D (nx9966), .CLK (nx10434)) ;
    dffr reg_current_state_4 (.Q (current_state_4), .QB (\$dummy [2746]), .D (
         next_state_4), .CLK (nx10428), .R (rst)) ;
    latch lat_next_state_4 (.Q (next_state_4), .D (nx322), .CLK (nx10434)) ;
    dff reg_next_state_dup_24 (.Q (next_state_dup_24), .QB (nx9866), .D (nx9748)
        , .CLK (nx10436)) ;
    or02 ix401 (.Y (ImgAddRST), .A0 (nx9952), .A1 (rst)) ;
    or02 ix403 (.Y (TriChnagerToaddEN), .A0 (current_state_6), .A1 (
         current_state_10)) ;
    oai21 ix455 (.Y (AddressChangerEN), .A0 (nx9875), .A1 (nx9883), .B0 (nx9893)
          ) ;
    nand04 ix9876 (.Y (nx9875), .A0 (DontRstIndicator), .A1 (nx9960), .A2 (nx418
           ), .A3 (nx9881)) ;
    or02 ix419 (.Y (nx418), .A0 (nx416), .A1 (lastFilter)) ;
    nor04 ix417 (.Y (nx416), .A0 (nx9879), .A1 (LayerInfoOut_3), .A2 (
          LayerInfoOut_2), .A3 (LayerInfoOut_1)) ;
    inv01 ix9880 (.Y (nx9879), .A (LayerInfoOut_0)) ;
    xnor2 ix9882 (.Y (nx9881), .A0 (ShiftLeftCounterOutput_4), .A1 (nx10378)) ;
    nand04 ix9884 (.Y (nx9883), .A0 (nx9885), .A1 (nx9887), .A2 (nx9889), .A3 (
           nx9891)) ;
    xnor2 ix9886 (.Y (nx9885), .A0 (ShiftLeftCounterOutput_0), .A1 (nx10392)) ;
    xnor2 ix9888 (.Y (nx9887), .A0 (ShiftLeftCounterOutput_1), .A1 (nx10388)) ;
    xnor2 ix9890 (.Y (nx9889), .A0 (ShiftLeftCounterOutput_2), .A1 (nx10386)) ;
    xnor2 ix9892 (.Y (nx9891), .A0 (ShiftLeftCounterOutput_3), .A1 (nx10382)) ;
    nand02 ix9894 (.Y (nx9893), .A0 (nx10310), .A1 (nx9966)) ;
    or03 ix461 (.Y (ShiftCounterRst), .A0 (nx456), .A1 (current_state_11), .A2 (
         rst)) ;
    and02 ix469 (.Y (ImgAddRegEN), .A0 (nx10028), .A1 (nx466)) ;
    nand04 ix467 (.Y (nx466), .A0 (nx9899), .A1 (nx9903), .A2 (nx9905), .A3 (
           nx9849)) ;
    aoi21 ix9900 (.Y (nx9899), .A0 (nx9901), .A1 (nx9964), .B0 (current_state_2)
          ) ;
    inv01 ix9902 (.Y (nx9901), .A (IndicatorI_0)) ;
    nor02_2x ix9904 (.Y (nx9903), .A0 (current_state_3), .A1 (current_state_6)
             ) ;
    aoi21 ix517 (.Y (FilterAddressEN), .A0 (nx9908), .A1 (nx9913), .B0 (
          LayerInfoOut_15)) ;
    aoi21 ix9909 (.Y (nx9908), .A0 (lastFilter), .A1 (current_state_6), .B0 (
          TriStateCounterEN)) ;
    inv01 ix507 (.Y (TriStateCounterEN), .A (nx9911)) ;
    oai21 ix9912 (.Y (nx9911), .A0 (current_state_0), .A1 (nx9972), .B0 (nx10310
          )) ;
    aoi32 ix9914 (.Y (nx9913), .A0 (nx494), .A1 (current_state_10), .A2 (nx418)
          , .B0 (nx10310), .B1 (nx350)) ;
    oai21 ix495 (.Y (nx494), .A0 (DontRstIndicator), .A1 (nx9916), .B0 (
          lastDepthOut)) ;
    nor03_2x ix9917 (.Y (nx9916), .A0 (nx482), .A1 (nx480), .A2 (nx478)) ;
    xor2 ix483 (.Y (nx482), .A0 (NumOfHeight_3), .A1 (nx10382)) ;
    xor2 ix481 (.Y (nx480), .A0 (NumOfHeight_2), .A1 (nx10386)) ;
    nand03 ix479 (.Y (nx478), .A0 (nx9921), .A1 (nx9923), .A2 (nx9925)) ;
    xnor2 ix9922 (.Y (nx9921), .A0 (NumOfHeight_0), .A1 (nx10394)) ;
    xnor2 ix9924 (.Y (nx9923), .A0 (NumOfHeight_4), .A1 (nx10378)) ;
    xnor2 ix9926 (.Y (nx9925), .A0 (NumOfHeight_1), .A1 (nx10390)) ;
    oai21 ix351 (.Y (nx350), .A0 (IndicatorF_0), .A1 (nx9870), .B0 (nx9905)) ;
    inv01 ix9930 (.Y (SwitchBar_0), .A (SwitchMEM_0)) ;
    nand04 ix397 (.Y (ReadI), .A0 (nx9932), .A1 (nx9934), .A2 (nx9899), .A3 (
           nx9903)) ;
    nor03_2x ix9933 (.Y (nx9932), .A0 (nx9966), .A1 (current_state_5), .A2 (
             nx9972)) ;
    nand03 ix9935 (.Y (nx9934), .A0 (nx382), .A1 (current_state_8), .A2 (nx9941)
           ) ;
    mux21 ix383 (.Y (nx382), .A0 (nx9937), .A1 (nx9939), .S0 (nx10406)) ;
    nor03_2x ix9938 (.Y (nx9937), .A0 (nx10410), .A1 (nx10408), .A2 (nx10412)) ;
    and03 ix9940 (.Y (nx9939), .A0 (nx10410), .A1 (nx10408), .A2 (nx10412)) ;
    or03 ix355 (.Y (ReadF), .A0 (current_state_0), .A1 (nx9972), .A2 (nx350)) ;
    tri01 tri_dmaStartSignal (.Y (dmaStartSignal), .A (PWR), .E (zero_11)) ;
    inv01 ix143 (.Y (nx142), .A (nx9903)) ;
    inv01 ix21 (.Y (nx20), .A (nx9765)) ;
    inv01 ix1 (.Y (CLK), .A (NOT_nx0)) ;
    inv01 ix9949 (.Y (nx9950), .A (nx9792)) ;
    inv01 ix9951 (.Y (nx9952), .A (nx9792)) ;
    inv01 ix9953 (.Y (nx9954), .A (nx9796)) ;
    inv01 ix9955 (.Y (nx9956), .A (nx9796)) ;
    buf02 ix9957 (.Y (nx9958), .A (current_state_9)) ;
    buf02 ix9959 (.Y (nx9960), .A (current_state_9)) ;
    inv01 ix9961 (.Y (nx9962), .A (nx9870)) ;
    inv01 ix9963 (.Y (nx9964), .A (nx9870)) ;
    buf02 ix9965 (.Y (nx9966), .A (current_state_4)) ;
    buf02 ix9967 (.Y (nx9968), .A (current_state_4)) ;
    inv02 ix9969 (.Y (nx9970), .A (nx9849)) ;
    inv02 ix9971 (.Y (nx9972), .A (nx9849)) ;
    buf02 ix9973 (.Y (nx9974), .A (FilterAddressOut_12)) ;
    buf02 ix9975 (.Y (nx9976), .A (FilterAddressOut_12)) ;
    buf02 ix9977 (.Y (nx9978), .A (FilterAddressOut_11)) ;
    buf02 ix9979 (.Y (nx9980), .A (FilterAddressOut_11)) ;
    buf02 ix9981 (.Y (nx9982), .A (FilterAddressOut_10)) ;
    buf02 ix9983 (.Y (nx9984), .A (FilterAddressOut_10)) ;
    buf02 ix9985 (.Y (nx9986), .A (FilterAddressOut_9)) ;
    buf02 ix9987 (.Y (nx9988), .A (FilterAddressOut_9)) ;
    buf02 ix9989 (.Y (nx9990), .A (FilterAddressOut_8)) ;
    buf02 ix9991 (.Y (nx9992), .A (FilterAddressOut_8)) ;
    buf02 ix9993 (.Y (nx9994), .A (FilterAddressOut_7)) ;
    buf02 ix9995 (.Y (nx9996), .A (FilterAddressOut_7)) ;
    buf02 ix9997 (.Y (nx9998), .A (FilterAddressOut_6)) ;
    buf02 ix9999 (.Y (nx10000), .A (FilterAddressOut_6)) ;
    buf02 ix10001 (.Y (nx10002), .A (FilterAddressOut_5)) ;
    buf02 ix10003 (.Y (nx10004), .A (FilterAddressOut_5)) ;
    buf02 ix10005 (.Y (nx10006), .A (FilterAddressOut_4)) ;
    buf02 ix10007 (.Y (nx10008), .A (FilterAddressOut_4)) ;
    buf02 ix10009 (.Y (nx10010), .A (FilterAddressOut_3)) ;
    buf02 ix10011 (.Y (nx10012), .A (FilterAddressOut_3)) ;
    buf02 ix10013 (.Y (nx10014), .A (FilterAddressOut_2)) ;
    buf02 ix10015 (.Y (nx10016), .A (FilterAddressOut_2)) ;
    buf02 ix10017 (.Y (nx10018), .A (FilterAddressOut_1)) ;
    buf02 ix10019 (.Y (nx10020), .A (FilterAddressOut_1)) ;
    buf02 ix10021 (.Y (nx10022), .A (FilterAddressOut_0)) ;
    buf02 ix10023 (.Y (nx10024), .A (FilterAddressOut_0)) ;
    buf02 ix10025 (.Y (nx10026), .A (ImgAddACKTriIN_0)) ;
    buf02 ix10027 (.Y (nx10028), .A (ImgAddACKTriIN_0)) ;
    inv02 ix10031 (.Y (nx10032), .A (nx10490)) ;
    inv02 ix10033 (.Y (nx10034), .A (nx10490)) ;
    inv02 ix10035 (.Y (nx10036), .A (nx10490)) ;
    inv02 ix10037 (.Y (nx10038), .A (nx10490)) ;
    inv02 ix10039 (.Y (nx10040), .A (nx10490)) ;
    inv02 ix10041 (.Y (nx10042), .A (nx10490)) ;
    inv02 ix10043 (.Y (nx10044), .A (nx10490)) ;
    inv02 ix10045 (.Y (nx10046), .A (nx10442)) ;
    inv02 ix10047 (.Y (nx10048), .A (nx10442)) ;
    inv02 ix10049 (.Y (nx10050), .A (nx10442)) ;
    inv02 ix10051 (.Y (nx10052), .A (nx10442)) ;
    inv02 ix10053 (.Y (nx10054), .A (nx10442)) ;
    inv02 ix10055 (.Y (nx10056), .A (nx10442)) ;
    inv02 ix10057 (.Y (nx10058), .A (nx10442)) ;
    inv02 ix10059 (.Y (nx10060), .A (nx10444)) ;
    inv02 ix10061 (.Y (nx10062), .A (nx10444)) ;
    inv02 ix10063 (.Y (nx10064), .A (nx10444)) ;
    inv02 ix10065 (.Y (nx10066), .A (nx10444)) ;
    inv02 ix10067 (.Y (nx10068), .A (nx10444)) ;
    inv02 ix10069 (.Y (nx10070), .A (nx10444)) ;
    inv02 ix10071 (.Y (nx10072), .A (nx10444)) ;
    inv02 ix10073 (.Y (nx10074), .A (nx10446)) ;
    inv02 ix10075 (.Y (nx10076), .A (nx10446)) ;
    inv02 ix10077 (.Y (nx10078), .A (nx10446)) ;
    inv02 ix10079 (.Y (nx10080), .A (nx10446)) ;
    inv02 ix10081 (.Y (nx10082), .A (nx10446)) ;
    inv02 ix10083 (.Y (nx10084), .A (nx10446)) ;
    inv02 ix10085 (.Y (nx10086), .A (nx10446)) ;
    inv02 ix10087 (.Y (nx10088), .A (nx10448)) ;
    inv02 ix10089 (.Y (nx10090), .A (nx10448)) ;
    inv02 ix10091 (.Y (nx10092), .A (nx10448)) ;
    inv02 ix10093 (.Y (nx10094), .A (nx10448)) ;
    inv02 ix10095 (.Y (nx10096), .A (nx10448)) ;
    inv02 ix10097 (.Y (nx10098), .A (nx10448)) ;
    inv02 ix10099 (.Y (nx10100), .A (nx10448)) ;
    inv02 ix10101 (.Y (nx10102), .A (nx10450)) ;
    inv02 ix10103 (.Y (nx10104), .A (nx10450)) ;
    inv02 ix10105 (.Y (nx10106), .A (nx10450)) ;
    inv02 ix10107 (.Y (nx10108), .A (nx10450)) ;
    inv02 ix10109 (.Y (nx10110), .A (nx10450)) ;
    inv02 ix10111 (.Y (nx10112), .A (nx10450)) ;
    inv02 ix10113 (.Y (nx10114), .A (nx10450)) ;
    inv02 ix10115 (.Y (nx10116), .A (nx10452)) ;
    inv02 ix10117 (.Y (nx10118), .A (nx10452)) ;
    inv02 ix10119 (.Y (nx10120), .A (nx10452)) ;
    inv02 ix10121 (.Y (nx10122), .A (nx10452)) ;
    inv02 ix10123 (.Y (nx10124), .A (nx10452)) ;
    inv02 ix10125 (.Y (nx10126), .A (nx10452)) ;
    inv02 ix10127 (.Y (nx10128), .A (nx10452)) ;
    inv02 ix10129 (.Y (nx10130), .A (nx10454)) ;
    inv02 ix10131 (.Y (nx10132), .A (nx10454)) ;
    inv02 ix10133 (.Y (nx10134), .A (nx10454)) ;
    inv02 ix10135 (.Y (nx10136), .A (nx10454)) ;
    inv02 ix10137 (.Y (nx10138), .A (nx10454)) ;
    inv02 ix10139 (.Y (nx10140), .A (nx10454)) ;
    inv02 ix10141 (.Y (nx10142), .A (nx10454)) ;
    inv02 ix10143 (.Y (nx10144), .A (nx10456)) ;
    inv02 ix10145 (.Y (nx10146), .A (nx10456)) ;
    inv02 ix10147 (.Y (nx10148), .A (nx10456)) ;
    inv02 ix10149 (.Y (nx10150), .A (nx10456)) ;
    inv02 ix10151 (.Y (nx10152), .A (nx10456)) ;
    inv02 ix10153 (.Y (nx10154), .A (nx10456)) ;
    inv02 ix10155 (.Y (nx10156), .A (nx10456)) ;
    inv02 ix10157 (.Y (nx10158), .A (nx10458)) ;
    inv02 ix10159 (.Y (nx10160), .A (nx10458)) ;
    inv02 ix10161 (.Y (nx10162), .A (nx10458)) ;
    inv02 ix10163 (.Y (nx10164), .A (nx10458)) ;
    inv02 ix10165 (.Y (nx10166), .A (nx10458)) ;
    inv02 ix10167 (.Y (nx10168), .A (nx10458)) ;
    inv02 ix10169 (.Y (nx10170), .A (nx10458)) ;
    inv02 ix10171 (.Y (nx10172), .A (nx10460)) ;
    inv02 ix10173 (.Y (nx10174), .A (nx10460)) ;
    inv02 ix10175 (.Y (nx10176), .A (nx10460)) ;
    inv02 ix10177 (.Y (nx10178), .A (nx10460)) ;
    inv02 ix10179 (.Y (nx10180), .A (nx10460)) ;
    inv02 ix10181 (.Y (nx10182), .A (nx10460)) ;
    inv02 ix10183 (.Y (nx10184), .A (nx10460)) ;
    inv02 ix10185 (.Y (nx10186), .A (nx10462)) ;
    inv02 ix10187 (.Y (nx10188), .A (nx10462)) ;
    inv02 ix10189 (.Y (nx10190), .A (nx10462)) ;
    inv02 ix10191 (.Y (nx10192), .A (nx10462)) ;
    inv02 ix10193 (.Y (nx10194), .A (nx10462)) ;
    inv02 ix10195 (.Y (nx10196), .A (nx10462)) ;
    inv02 ix10197 (.Y (nx10198), .A (nx10462)) ;
    inv02 ix10199 (.Y (nx10200), .A (nx10464)) ;
    inv02 ix10201 (.Y (nx10202), .A (nx10464)) ;
    inv02 ix10203 (.Y (nx10204), .A (nx10464)) ;
    inv02 ix10205 (.Y (nx10206), .A (nx10464)) ;
    inv02 ix10207 (.Y (nx10208), .A (nx10464)) ;
    inv02 ix10209 (.Y (nx10210), .A (nx10464)) ;
    inv02 ix10211 (.Y (nx10212), .A (nx10464)) ;
    inv02 ix10213 (.Y (nx10214), .A (nx10466)) ;
    inv02 ix10215 (.Y (nx10216), .A (nx10466)) ;
    inv02 ix10217 (.Y (nx10218), .A (nx10466)) ;
    inv02 ix10219 (.Y (nx10220), .A (nx10466)) ;
    inv02 ix10221 (.Y (nx10222), .A (nx10466)) ;
    inv02 ix10223 (.Y (nx10224), .A (nx10466)) ;
    inv02 ix10225 (.Y (nx10226), .A (nx10466)) ;
    inv02 ix10227 (.Y (nx10228), .A (nx10468)) ;
    inv02 ix10229 (.Y (nx10230), .A (nx10468)) ;
    inv02 ix10231 (.Y (nx10232), .A (nx10468)) ;
    inv02 ix10233 (.Y (nx10234), .A (nx10468)) ;
    inv02 ix10235 (.Y (nx10236), .A (nx10468)) ;
    inv02 ix10237 (.Y (nx10238), .A (nx10468)) ;
    inv02 ix10239 (.Y (nx10240), .A (nx10468)) ;
    inv02 ix10241 (.Y (nx10242), .A (nx10470)) ;
    inv02 ix10243 (.Y (nx10244), .A (nx10470)) ;
    inv02 ix10245 (.Y (nx10246), .A (nx10470)) ;
    inv02 ix10247 (.Y (nx10248), .A (nx10470)) ;
    inv02 ix10249 (.Y (nx10250), .A (nx10470)) ;
    inv02 ix10251 (.Y (nx10252), .A (nx10470)) ;
    inv02 ix10253 (.Y (nx10254), .A (nx10470)) ;
    inv02 ix10255 (.Y (nx10256), .A (nx10472)) ;
    inv02 ix10257 (.Y (nx10258), .A (nx10472)) ;
    inv02 ix10259 (.Y (nx10260), .A (nx10472)) ;
    inv02 ix10261 (.Y (nx10262), .A (nx10472)) ;
    inv02 ix10263 (.Y (nx10264), .A (nx10472)) ;
    inv02 ix10265 (.Y (nx10266), .A (nx10472)) ;
    inv02 ix10267 (.Y (nx10268), .A (nx10472)) ;
    inv02 ix10269 (.Y (nx10270), .A (nx10474)) ;
    inv02 ix10271 (.Y (nx10272), .A (nx10474)) ;
    inv02 ix10273 (.Y (nx10274), .A (nx10474)) ;
    inv02 ix10275 (.Y (nx10276), .A (nx10474)) ;
    inv02 ix10277 (.Y (nx10278), .A (nx10474)) ;
    inv02 ix10279 (.Y (nx10280), .A (nx10474)) ;
    inv02 ix10281 (.Y (nx10282), .A (nx10474)) ;
    inv02 ix10283 (.Y (nx10284), .A (nx10476)) ;
    inv02 ix10285 (.Y (nx10286), .A (nx10476)) ;
    inv02 ix10287 (.Y (nx10288), .A (nx10476)) ;
    inv02 ix10289 (.Y (nx10290), .A (nx10476)) ;
    inv02 ix10291 (.Y (nx10292), .A (nx10476)) ;
    inv02 ix10293 (.Y (nx10294), .A (nx10476)) ;
    inv02 ix10295 (.Y (nx10296), .A (nx10476)) ;
    inv02 ix10297 (.Y (nx10298), .A (nx10478)) ;
    inv02 ix10299 (.Y (nx10300), .A (nx10478)) ;
    inv02 ix10301 (.Y (nx10302), .A (nx10478)) ;
    inv02 ix10303 (.Y (nx10304), .A (nx10478)) ;
    inv02 ix10305 (.Y (nx10306), .A (nx10478)) ;
    buf02 ix10307 (.Y (nx10308), .A (ACKF)) ;
    buf02 ix10309 (.Y (nx10310), .A (ACKF)) ;
    buf02 ix10311 (.Y (nx10312), .A (DataIOut_15)) ;
    buf02 ix10313 (.Y (nx10314), .A (DataIOut_15)) ;
    buf02 ix10315 (.Y (nx10316), .A (DataIOut_14)) ;
    buf02 ix10317 (.Y (nx10318), .A (DataIOut_14)) ;
    buf02 ix10319 (.Y (nx10320), .A (DataIOut_13)) ;
    buf02 ix10321 (.Y (nx10322), .A (DataIOut_13)) ;
    buf02 ix10323 (.Y (nx10324), .A (DataIOut_12)) ;
    buf02 ix10325 (.Y (nx10326), .A (DataIOut_12)) ;
    buf02 ix10327 (.Y (nx10328), .A (DataIOut_11)) ;
    buf02 ix10329 (.Y (nx10330), .A (DataIOut_11)) ;
    buf02 ix10331 (.Y (nx10332), .A (DataIOut_10)) ;
    buf02 ix10333 (.Y (nx10334), .A (DataIOut_10)) ;
    buf02 ix10335 (.Y (nx10336), .A (DataIOut_9)) ;
    buf02 ix10337 (.Y (nx10338), .A (DataIOut_9)) ;
    buf02 ix10339 (.Y (nx10340), .A (DataIOut_8)) ;
    buf02 ix10341 (.Y (nx10342), .A (DataIOut_8)) ;
    buf02 ix10343 (.Y (nx10344), .A (DataIOut_7)) ;
    buf02 ix10345 (.Y (nx10346), .A (DataIOut_7)) ;
    buf02 ix10347 (.Y (nx10348), .A (DataIOut_6)) ;
    buf02 ix10349 (.Y (nx10350), .A (DataIOut_6)) ;
    buf02 ix10351 (.Y (nx10352), .A (DataIOut_5)) ;
    buf02 ix10353 (.Y (nx10354), .A (DataIOut_5)) ;
    buf02 ix10355 (.Y (nx10356), .A (DataIOut_4)) ;
    buf02 ix10357 (.Y (nx10358), .A (DataIOut_4)) ;
    buf02 ix10359 (.Y (nx10360), .A (DataIOut_3)) ;
    buf02 ix10361 (.Y (nx10362), .A (DataIOut_3)) ;
    buf02 ix10363 (.Y (nx10364), .A (DataIOut_2)) ;
    buf02 ix10365 (.Y (nx10366), .A (DataIOut_2)) ;
    buf02 ix10367 (.Y (nx10368), .A (DataIOut_1)) ;
    buf02 ix10369 (.Y (nx10370), .A (DataIOut_1)) ;
    buf02 ix10371 (.Y (nx10372), .A (DataIOut_0)) ;
    buf02 ix10373 (.Y (nx10374), .A (DataIOut_0)) ;
    buf02 ix10375 (.Y (nx10376), .A (LayerInfoOut_8)) ;
    buf02 ix10377 (.Y (nx10378), .A (LayerInfoOut_8)) ;
    buf02 ix10379 (.Y (nx10380), .A (LayerInfoOut_7)) ;
    buf02 ix10381 (.Y (nx10382), .A (LayerInfoOut_7)) ;
    buf02 ix10383 (.Y (nx10384), .A (LayerInfoOut_6)) ;
    buf02 ix10385 (.Y (nx10386), .A (LayerInfoOut_6)) ;
    buf02 ix10387 (.Y (nx10388), .A (LayerInfoOut_5)) ;
    buf02 ix10389 (.Y (nx10390), .A (LayerInfoOut_5)) ;
    buf02 ix10391 (.Y (nx10392), .A (LayerInfoOut_4)) ;
    buf02 ix10393 (.Y (nx10394), .A (LayerInfoOut_4)) ;
    buf02 ix10395 (.Y (nx10396), .A (ConvOuput_15)) ;
    buf02 ix10397 (.Y (nx10398), .A (NumOfFilters_3)) ;
    buf02 ix10399 (.Y (nx10400), .A (NumOfFilters_2)) ;
    buf02 ix10401 (.Y (nx10402), .A (NumOfFilters_1)) ;
    buf02 ix10403 (.Y (nx10404), .A (NumOfFilters_0)) ;
    buf02 ix10405 (.Y (nx10406), .A (CNDepthoutput_3)) ;
    buf02 ix10407 (.Y (nx10408), .A (CNDepthoutput_2)) ;
    buf02 ix10409 (.Y (nx10410), .A (CNDepthoutput_1)) ;
    buf02 ix10411 (.Y (nx10412), .A (CNDepthoutput_0)) ;
    inv02 ix10413 (.Y (nx10414), .A (nx10436)) ;
    inv02 ix10415 (.Y (nx10416), .A (nx10436)) ;
    inv02 ix10417 (.Y (nx10418), .A (nx10436)) ;
    inv02 ix10419 (.Y (nx10420), .A (nx10436)) ;
    inv02 ix10421 (.Y (nx10422), .A (nx10438)) ;
    inv02 ix10423 (.Y (nx10424), .A (nx10438)) ;
    inv02 ix10425 (.Y (nx10426), .A (nx10438)) ;
    inv02 ix10427 (.Y (nx10428), .A (nx10438)) ;
    inv02 ix10429 (.Y (nx10430), .A (nx10438)) ;
    inv02 ix10431 (.Y (nx10432), .A (done)) ;
    inv02 ix10433 (.Y (nx10434), .A (done)) ;
    inv02 ix10435 (.Y (nx10436), .A (CLK)) ;
    inv02 ix10437 (.Y (nx10438), .A (CLK)) ;
    inv02 ix10439 (.Y (nx10440), .A (DataFOut_399)) ;
    inv02 ix10441 (.Y (nx10442), .A (nx10484)) ;
    inv02 ix10443 (.Y (nx10444), .A (nx10484)) ;
    inv02 ix10445 (.Y (nx10446), .A (nx10484)) ;
    inv02 ix10447 (.Y (nx10448), .A (nx10484)) ;
    inv02 ix10449 (.Y (nx10450), .A (nx10484)) ;
    inv02 ix10451 (.Y (nx10452), .A (nx10484)) ;
    inv02 ix10453 (.Y (nx10454), .A (nx10484)) ;
    inv02 ix10455 (.Y (nx10456), .A (nx10486)) ;
    inv02 ix10457 (.Y (nx10458), .A (nx10486)) ;
    inv02 ix10459 (.Y (nx10460), .A (nx10486)) ;
    inv02 ix10461 (.Y (nx10462), .A (nx10486)) ;
    inv02 ix10463 (.Y (nx10464), .A (nx10486)) ;
    inv02 ix10465 (.Y (nx10466), .A (nx10486)) ;
    inv02 ix10467 (.Y (nx10468), .A (nx10486)) ;
    inv02 ix10469 (.Y (nx10470), .A (nx10488)) ;
    inv02 ix10471 (.Y (nx10472), .A (nx10488)) ;
    inv02 ix10473 (.Y (nx10474), .A (nx10488)) ;
    inv02 ix10475 (.Y (nx10476), .A (nx10488)) ;
    inv02 ix10477 (.Y (nx10478), .A (nx10488)) ;
    inv02 ix10483 (.Y (nx10484), .A (nx10440)) ;
    inv02 ix10485 (.Y (nx10486), .A (nx10440)) ;
    inv02 ix10487 (.Y (nx10488), .A (nx10440)) ;
    inv02 ix10489 (.Y (nx10490), .A (DataFOut_399)) ;
    oai22 ix241 (.Y (nx240), .A0 (X), .A1 (nx10496), .B0 (nx9768), .B1 (nx20)) ;
    inv01 ix10495 (.Y (nx10496), .A (nx9960)) ;
    nand03 ix187 (.Y (nx186), .A0 (nx9870), .A1 (nx10498), .A2 (nx180)) ;
    inv01 ix10497 (.Y (nx10498), .A (nx9958)) ;
    nor02ii ix301 (.Y (nx300), .A0 (nx9792), .A1 (next_state_dup_134)) ;
    nor02ii ix113 (.Y (nx112), .A0 (nx9849), .A1 (next_state_dup_26)) ;
    nor02_2x ix323 (.Y (nx322), .A0 (nx9866), .A1 (nx9849)) ;
    mux21_ni ix9749 (.Y (nx9748), .A0 (next_state_dup_24), .A1 (nx10478), .S0 (
             nx10308)) ;
    nor02_2x ix457 (.Y (nx456), .A0 (nx9765), .A1 (nx9870)) ;
    nor02ii ix9906 (.Y (nx9905), .A0 (nx9966), .A1 (nx9858)) ;
    nor02ii ix519 (.Y (SwitchClk), .A0 (nx9792), .A1 (nx10028)) ;
    latchr lat_SaveAckLatch_u1 (.QB (nx5), .D (nx9063), .CLK (nx186), .R (
           zero_11)) ;
    inv01 lat_SaveAckLatch_u2 (.Y (SaveAckLatch), .A (nx5)) ;
    buf02 lat_SaveAckLatch_u3 (.Y (nx9941), .A (nx5)) ;
    buf02 ix10499 (.Y (nx10500), .A (LayerInfoOut_14)) ;
    buf02 ix10501 (.Y (nx10502), .A (LayerInfoOut_14)) ;
    inv02 ix10503 (.Y (nx10504), .A (nx10438)) ;
endmodule


module outWidthState ( currentState, infoReg, address, outWidth ) ;

    input [14:0]currentState ;
    input [15:0]infoReg ;
    output [12:0]address ;
    output [15:0]outWidth ;

    wire nx263, nx268, nx271, nx274, nx277, nx280, nx311, nx313, nx315, nx317, 
         nx319, nx321;



    fake_vcc ix264 (.Y (nx263)) ;
    tri01 tri_outwidthbefore_0 (.Y (outWidth[0]), .A (nx268), .E (nx313)) ;
    inv01 ix269 (.Y (nx268), .A (infoReg[4])) ;
    tri01 tri_outwidthbefore_1 (.Y (outWidth[1]), .A (nx271), .E (nx313)) ;
    inv01 ix272 (.Y (nx271), .A (infoReg[5])) ;
    tri01 tri_outwidthbefore_2 (.Y (outWidth[2]), .A (nx274), .E (nx313)) ;
    inv01 ix275 (.Y (nx274), .A (infoReg[6])) ;
    tri01 tri_outwidthbefore_3 (.Y (outWidth[3]), .A (nx277), .E (nx313)) ;
    inv01 ix278 (.Y (nx277), .A (infoReg[7])) ;
    tri01 tri_outwidthbefore_4 (.Y (outWidth[4]), .A (nx280), .E (nx313)) ;
    inv01 ix281 (.Y (nx280), .A (infoReg[8])) ;
    tri01 tri_outwidthbefore_5 (.Y (outWidth[5]), .A (nx263), .E (nx313)) ;
    tri01 tri_outwidthbefore_6 (.Y (outWidth[6]), .A (nx263), .E (nx313)) ;
    tri01 tri_outwidthbefore_7 (.Y (outWidth[7]), .A (nx263), .E (nx315)) ;
    tri01 tri_outwidthbefore_8 (.Y (outWidth[8]), .A (nx263), .E (nx315)) ;
    tri01 tri_outwidthbefore_9 (.Y (outWidth[9]), .A (nx263), .E (nx315)) ;
    tri01 tri_outwidthbefore_10 (.Y (outWidth[10]), .A (nx263), .E (nx315)) ;
    tri01 tri_outwidthbefore_11 (.Y (outWidth[11]), .A (nx263), .E (nx315)) ;
    tri01 tri_outwidthbefore_12 (.Y (outWidth[12]), .A (nx263), .E (nx315)) ;
    tri01 tri_outwidthbefore_13 (.Y (outWidth[13]), .A (nx263), .E (nx315)) ;
    tri01 tri_outwidthbefore_14 (.Y (outWidth[14]), .A (nx263), .E (nx317)) ;
    tri01 tri_outwidthbefore_15 (.Y (outWidth[15]), .A (nx263), .E (nx317)) ;
    tri01 tri_address_0 (.Y (address[0]), .A (nx263), .E (nx317)) ;
    tri01 tri_address_1 (.Y (address[1]), .A (nx263), .E (nx317)) ;
    tri01 tri_address_2 (.Y (address[2]), .A (nx263), .E (nx317)) ;
    tri01 tri_address_3 (.Y (address[3]), .A (nx263), .E (nx317)) ;
    tri01 tri_address_4 (.Y (address[4]), .A (nx263), .E (nx317)) ;
    tri01 tri_address_5 (.Y (address[5]), .A (nx263), .E (nx319)) ;
    tri01 tri_address_6 (.Y (address[6]), .A (nx263), .E (nx319)) ;
    tri01 tri_address_7 (.Y (address[7]), .A (nx263), .E (nx319)) ;
    tri01 tri_address_8 (.Y (address[8]), .A (nx263), .E (nx319)) ;
    tri01 tri_address_9 (.Y (address[9]), .A (nx263), .E (nx319)) ;
    tri01 tri_address_10 (.Y (address[10]), .A (nx263), .E (nx319)) ;
    tri01 tri_address_11 (.Y (address[11]), .A (nx263), .E (nx319)) ;
    tri01 tri_address_12 (.Y (address[12]), .A (nx263), .E (nx321)) ;
    inv01 ix310 (.Y (nx311), .A (currentState[13])) ;
    inv01 ix312 (.Y (nx313), .A (nx311)) ;
    inv01 ix314 (.Y (nx315), .A (nx311)) ;
    inv01 ix316 (.Y (nx317), .A (nx311)) ;
    inv01 ix318 (.Y (nx319), .A (nx311)) ;
    inv01 ix320 (.Y (nx321), .A (nx311)) ;
endmodule


module StateChecks ( current_state, noOfLayers, LayerInfo, CLK, RST, L, D, 
                     CNDoutput, CNLoutput ) ;

    input [14:0]current_state ;
    input [15:0]noOfLayers ;
    input [15:0]LayerInfo ;
    input CLK ;
    input RST ;
    output L ;
    output D ;
    output [3:0]CNDoutput ;
    output [1:0]CNLoutput ;

    wire DepthCounterRst, SDbar, GND0, PWR, nx62, nx64, nx67, nx69, nx71, nx73;



    Counter_4 counterNoDepth0 (.enable (PWR), .reset (DepthCounterRst), .clk (
              current_state[12]), .load (GND0), .\output  ({CNDoutput[3],
              CNDoutput[2],CNDoutput[1],CNDoutput[0]}), .\input  ({GND0,GND0,
              GND0,PWR})) ;
    Counter_2 counterNoLayer0 (.enable (PWR), .reset (RST), .clk (SDbar), .load (
              GND0), .\output  ({CNLoutput[1],CNLoutput[0]}), .\input  ({GND0,
              PWR})) ;
    fake_vcc ix44 (.Y (PWR)) ;
    fake_gnd ix42 (.Y (GND0)) ;
    nand02 ix5 (.Y (L), .A0 (nx62), .A1 (nx64)) ;
    xnor2 ix63 (.Y (nx62), .A0 (CNLoutput[1]), .A1 (noOfLayers[1])) ;
    xnor2 ix65 (.Y (nx64), .A0 (CNLoutput[0]), .A1 (noOfLayers[0])) ;
    nand04 ix19 (.Y (D), .A0 (nx67), .A1 (nx69), .A2 (nx71), .A3 (nx73)) ;
    xnor2 ix68 (.Y (nx67), .A0 (CNDoutput[3]), .A1 (LayerInfo[12])) ;
    xnor2 ix70 (.Y (nx69), .A0 (CNDoutput[2]), .A1 (LayerInfo[11])) ;
    xnor2 ix72 (.Y (nx71), .A0 (CNDoutput[1]), .A1 (LayerInfo[10])) ;
    xnor2 ix74 (.Y (nx73), .A0 (CNDoutput[0]), .A1 (LayerInfo[9])) ;
    or02 ix23 (.Y (DepthCounterRst), .A0 (RST), .A1 (current_state[13])) ;
    inv01 ix76 (.Y (SDbar), .A (D)) ;
endmodule


module ImageState ( current_state, WSquared, AddresCounterIN, AddresCounterLoad, 
                    NoOfShiftsCounter, LayerInfoIn, CLK, RST, Q, NumOfFilters, 
                    NumOfHeight, X1, Y1, K1 ) ;

    input [14:0]current_state ;
    input [9:0]WSquared ;
    input [12:0]AddresCounterIN ;
    output [12:0]AddresCounterLoad ;
    input [4:0]NoOfShiftsCounter ;
    input [15:0]LayerInfoIn ;
    input CLK ;
    input RST ;
    output Q ;
    output [3:0]NumOfFilters ;
    output [4:0]NumOfHeight ;
    output X1 ;
    output Y1 ;
    output K1 ;

    wire Qbar_0, newSliceRegOUT_12, newSliceRegOUT_11, newSliceRegOUT_10, 
         newSliceRegOUT_9, newSliceRegOUT_8, newSliceRegOUT_7, newSliceRegOUT_6, 
         newSliceRegOUT_5, newSliceRegOUT_4, newSliceRegOUT_3, newSliceRegOUT_2, 
         newSliceRegOUT_1, newSliceRegOUT_0, adder0Out_12, adder0Out_11, 
         adder0Out_10, adder0Out_9, adder0Out_8, adder0Out_7, adder0Out_6, 
         adder0Out_5, adder0Out_4, adder0Out_3, adder0Out_2, adder0Out_1, 
         adder0Out_0, adder1Out_12, adder1Out_11, adder1Out_10, adder1Out_9, 
         adder1Out_8, adder1Out_7, adder1Out_6, adder1Out_5, adder1Out_4, 
         adder1Out_3, adder1Out_2, adder1Out_1, adder1Out_0, QRST, cnhRST, 
         cnfCLK, FilterCounterRst, newSliceRegRST, newSliceRegEn, 
         triStateBuffer1EN, PWR, adder0b_12, YBar, nx253, nx255, nx257, nx259, 
         nx264, nx266, nx268, nx270, nx272, nx274, nx278, nx280, nx282, nx284, 
         nx286, nx288, nx295, nx297, nx300, nx310, nx316, nx318, nx320, nx322, 
         nx324;
    wire [1:0] \$dummy ;




    nBitRegister_1 DDF0 (.D ({Qbar_0}), .CLK (nx310), .RST (QRST), .EN (PWR), .Q (
                   {Q})) ;
    Counter_5 counterNoHeight0 (.enable (PWR), .reset (cnhRST), .clk (YBar), .load (
              adder0b_12), .\output  ({NumOfHeight[4],NumOfHeight[3],
              NumOfHeight[2],NumOfHeight[1],NumOfHeight[0]}), .\input  ({
              adder0b_12,adder0b_12,adder0b_12,adder0b_12,PWR})) ;
    Counter_4 counterNoFilters0 (.enable (PWR), .reset (FilterCounterRst), .clk (
              nx310), .load (adder0b_12), .\output  ({NumOfFilters[3],
              NumOfFilters[2],NumOfFilters[1],NumOfFilters[0]}), .\input  ({
              adder0b_12,adder0b_12,adder0b_12,PWR})) ;
    nBitRegister_13 newSliceReg0 (.D ({adder0Out_12,adder0Out_11,adder0Out_10,
                    adder0Out_9,adder0Out_8,adder0Out_7,adder0Out_6,adder0Out_5,
                    adder0Out_4,adder0Out_3,adder0Out_2,adder0Out_1,adder0Out_0}
                    ), .CLK (CLK), .RST (newSliceRegRST), .EN (newSliceRegEn), .Q (
                    {newSliceRegOUT_12,newSliceRegOUT_11,newSliceRegOUT_10,
                    newSliceRegOUT_9,newSliceRegOUT_8,newSliceRegOUT_7,
                    newSliceRegOUT_6,newSliceRegOUT_5,newSliceRegOUT_4,
                    newSliceRegOUT_3,newSliceRegOUT_2,newSliceRegOUT_1,
                    newSliceRegOUT_0})) ;
    my_nadder_13 adder0 (.a ({newSliceRegOUT_12,newSliceRegOUT_11,
                 newSliceRegOUT_10,newSliceRegOUT_9,newSliceRegOUT_8,
                 newSliceRegOUT_7,newSliceRegOUT_6,newSliceRegOUT_5,
                 newSliceRegOUT_4,newSliceRegOUT_3,newSliceRegOUT_2,
                 newSliceRegOUT_1,newSliceRegOUT_0}), .b ({adder0b_12,adder0b_12
                 ,adder0b_12,adder0b_12,adder0b_12,adder0b_12,adder0b_12,
                 adder0b_12,nx316,nx318,nx320,nx322,nx324}), .cin (adder0b_12), 
                 .s ({adder0Out_12,adder0Out_11,adder0Out_10,adder0Out_9,
                 adder0Out_8,adder0Out_7,adder0Out_6,adder0Out_5,adder0Out_4,
                 adder0Out_3,adder0Out_2,adder0Out_1,adder0Out_0}), .cout (
                 \$dummy [0])) ;
    triStateBuffer_13 triStateBuffer0 (.D ({adder0Out_12,adder0Out_11,
                      adder0Out_10,adder0Out_9,adder0Out_8,adder0Out_7,
                      adder0Out_6,adder0Out_5,adder0Out_4,adder0Out_3,
                      adder0Out_2,adder0Out_1,adder0Out_0}), .EN (newSliceRegEn)
                      , .F ({AddresCounterLoad[12],AddresCounterLoad[11],
                      AddresCounterLoad[10],AddresCounterLoad[9],
                      AddresCounterLoad[8],AddresCounterLoad[7],
                      AddresCounterLoad[6],AddresCounterLoad[5],
                      AddresCounterLoad[4],AddresCounterLoad[3],
                      AddresCounterLoad[2],AddresCounterLoad[1],
                      AddresCounterLoad[0]})) ;
    my_nadder_13 adder1 (.a ({AddresCounterIN[12],AddresCounterIN[11],
                 AddresCounterIN[10],AddresCounterIN[9],AddresCounterIN[8],
                 AddresCounterIN[7],AddresCounterIN[6],AddresCounterIN[5],
                 AddresCounterIN[4],AddresCounterIN[3],AddresCounterIN[2],
                 AddresCounterIN[1],AddresCounterIN[0]}), .b ({adder0b_12,
                 adder0b_12,adder0b_12,WSquared[9],WSquared[8],WSquared[7],
                 WSquared[6],WSquared[5],WSquared[4],WSquared[3],WSquared[2],
                 WSquared[1],WSquared[0]}), .cin (adder0b_12), .s ({adder1Out_12
                 ,adder1Out_11,adder1Out_10,adder1Out_9,adder1Out_8,adder1Out_7,
                 adder1Out_6,adder1Out_5,adder1Out_4,adder1Out_3,adder1Out_2,
                 adder1Out_1,adder1Out_0}), .cout (\$dummy [1])) ;
    triStateBuffer_13 triStateBuffer1 (.D ({adder1Out_12,adder1Out_11,
                      adder1Out_10,adder1Out_9,adder1Out_8,adder1Out_7,
                      adder1Out_6,adder1Out_5,adder1Out_4,adder1Out_3,
                      adder1Out_2,adder1Out_1,adder1Out_0}), .EN (
                      triStateBuffer1EN), .F ({AddresCounterLoad[12],
                      AddresCounterLoad[11],AddresCounterLoad[10],
                      AddresCounterLoad[9],AddresCounterLoad[8],
                      AddresCounterLoad[7],AddresCounterLoad[6],
                      AddresCounterLoad[5],AddresCounterLoad[4],
                      AddresCounterLoad[3],AddresCounterLoad[2],
                      AddresCounterLoad[1],AddresCounterLoad[0]})) ;
    xnor2 ix254 (.Y (nx253), .A0 (LayerInfoIn[3]), .A1 (NumOfFilters[3])) ;
    xnor2 ix256 (.Y (nx255), .A0 (LayerInfoIn[2]), .A1 (NumOfFilters[2])) ;
    xnor2 ix258 (.Y (nx257), .A0 (LayerInfoIn[1]), .A1 (NumOfFilters[1])) ;
    xnor2 ix260 (.Y (nx259), .A0 (LayerInfoIn[0]), .A1 (NumOfFilters[0])) ;
    fake_gnd ix221 (.Y (adder0b_12)) ;
    fake_vcc ix219 (.Y (PWR)) ;
    nand04 ix17 (.Y (K1), .A0 (nx264), .A1 (nx270), .A2 (nx272), .A3 (nx274)) ;
    and02 ix265 (.Y (nx264), .A0 (nx266), .A1 (nx268)) ;
    xnor2 ix267 (.Y (nx266), .A0 (nx318), .A1 (NumOfHeight[3])) ;
    xnor2 ix269 (.Y (nx268), .A0 (nx320), .A1 (NumOfHeight[2])) ;
    xnor2 ix271 (.Y (nx270), .A0 (nx324), .A1 (NumOfHeight[0])) ;
    xnor2 ix273 (.Y (nx272), .A0 (nx316), .A1 (NumOfHeight[4])) ;
    xnor2 ix275 (.Y (nx274), .A0 (nx322), .A1 (NumOfHeight[1])) ;
    nand04 ix49 (.Y (Y1), .A0 (nx253), .A1 (nx255), .A2 (nx257), .A3 (nx259)) ;
    nand04 ix35 (.Y (X1), .A0 (nx278), .A1 (nx284), .A2 (nx286), .A3 (nx288)) ;
    and02 ix279 (.Y (nx278), .A0 (nx280), .A1 (nx282)) ;
    xnor2 ix281 (.Y (nx280), .A0 (nx318), .A1 (NoOfShiftsCounter[3])) ;
    xnor2 ix283 (.Y (nx282), .A0 (nx320), .A1 (NoOfShiftsCounter[2])) ;
    xnor2 ix285 (.Y (nx284), .A0 (nx324), .A1 (NoOfShiftsCounter[0])) ;
    xnor2 ix287 (.Y (nx286), .A0 (nx316), .A1 (NoOfShiftsCounter[4])) ;
    xnor2 ix289 (.Y (nx288), .A0 (nx322), .A1 (NoOfShiftsCounter[1])) ;
    nor02ii ix61 (.Y (triStateBuffer1EN), .A0 (newSliceRegEn), .A1 (nx310)) ;
    nor02ii ix53 (.Y (newSliceRegEn), .A0 (Y1), .A1 (current_state[9])) ;
    nor02ii ix57 (.Y (cnfCLK), .A0 (X1), .A1 (current_state[9])) ;
    or02 ix63 (.Y (newSliceRegRST), .A0 (RST), .A1 (current_state[12])) ;
    oai21 ix69 (.Y (FilterCounterRst), .A0 (nx295), .A1 (Y1), .B0 (nx297)) ;
    inv01 ix296 (.Y (nx295), .A (current_state[11])) ;
    inv01 ix298 (.Y (nx297), .A (RST)) ;
    oai21 ix77 (.Y (cnhRST), .A0 (nx300), .A1 (K1), .B0 (nx297)) ;
    inv01 ix301 (.Y (nx300), .A (current_state[12])) ;
    or02 ix79 (.Y (QRST), .A0 (RST), .A1 (current_state[13])) ;
    inv01 ix304 (.Y (Qbar_0), .A (Q)) ;
    inv01 ix252 (.Y (YBar), .A (Y1)) ;
    buf02 ix309 (.Y (nx310), .A (cnfCLK)) ;
    buf02 ix315 (.Y (nx316), .A (LayerInfoIn[8])) ;
    buf02 ix317 (.Y (nx318), .A (LayerInfoIn[7])) ;
    buf02 ix319 (.Y (nx320), .A (LayerInfoIn[6])) ;
    buf02 ix321 (.Y (nx322), .A (LayerInfoIn[5])) ;
    buf02 ix323 (.Y (nx324), .A (LayerInfoIn[4])) ;
endmodule


module Counter_4 ( enable, reset, clk, load, \output , \input  ) ;

    input enable ;
    input reset ;
    input clk ;
    input load ;
    output [3:0]\output  ;
    input [3:0]\input  ;

    wire addResult_3, addResult_2, addResult_1, addResult_0, one_0, one_3, nx52, 
         NOT_clk, nx8, nx12, nx46, nx20, nx24, nx40, nx32, nx36, nx34, nx45, 
         nx49, nx143, nx153, nx163, nx173, nx182, nx216;
    wire [8:0] \$dummy ;




    my_nadder_4 A1 (.a ({\output [3],\output [2],\output [1],\output [0]}), .b (
                {one_3,one_3,one_3,one_0}), .cin (one_3), .s ({addResult_3,
                addResult_2,addResult_1,addResult_0}), .cout (\$dummy [0])) ;
    fake_gnd ix120 (.Y (one_3)) ;
    fake_vcc ix118 (.Y (one_0)) ;
    dffsr_ni reg_toOutput_0__dup_1 (.Q (\output [0]), .QB (\$dummy [1]), .D (
             nx143), .CLK (clk), .S (nx8), .R (nx12)) ;
    mux21_ni ix144 (.Y (nx143), .A0 (\output [0]), .A1 (addResult_0), .S0 (
             enable)) ;
    nor02ii ix9 (.Y (nx8), .A0 (nx182), .A1 (nx52)) ;
    nor02_2x ix183 (.Y (nx182), .A0 (nx216), .A1 (load)) ;
    dffr ix53 (.Q (nx52), .QB (\$dummy [2]), .D (\input [0]), .CLK (NOT_clk), .R (
         nx216)) ;
    inv01 ix186 (.Y (NOT_clk), .A (clk)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (nx52), .A1 (nx182)) ;
    dffsr_ni reg_toOutput_1__dup_1 (.Q (\output [1]), .QB (\$dummy [3]), .D (
             nx153), .CLK (clk), .S (nx20), .R (nx24)) ;
    mux21_ni ix154 (.Y (nx153), .A0 (\output [1]), .A1 (addResult_1), .S0 (
             enable)) ;
    nor02ii ix21 (.Y (nx20), .A0 (nx182), .A1 (nx46)) ;
    dffr ix47 (.Q (nx46), .QB (\$dummy [4]), .D (\input [1]), .CLK (NOT_clk), .R (
         nx216)) ;
    nor02_2x ix25 (.Y (nx24), .A0 (nx46), .A1 (nx182)) ;
    dffsr_ni reg_toOutput_2__dup_1 (.Q (\output [2]), .QB (\$dummy [5]), .D (
             nx163), .CLK (clk), .S (nx32), .R (nx36)) ;
    mux21_ni ix164 (.Y (nx163), .A0 (\output [2]), .A1 (addResult_2), .S0 (
             enable)) ;
    nor02ii ix33 (.Y (nx32), .A0 (nx182), .A1 (nx40)) ;
    dffr ix41 (.Q (nx40), .QB (\$dummy [6]), .D (\input [2]), .CLK (NOT_clk), .R (
         nx216)) ;
    nor02_2x ix37 (.Y (nx36), .A0 (nx40), .A1 (nx182)) ;
    dffsr_ni reg_toOutput_3__dup_1 (.Q (\output [3]), .QB (\$dummy [7]), .D (
             nx173), .CLK (clk), .S (nx45), .R (nx49)) ;
    mux21_ni ix174 (.Y (nx173), .A0 (\output [3]), .A1 (addResult_3), .S0 (
             enable)) ;
    nor02ii ix46 (.Y (nx45), .A0 (nx182), .A1 (nx34)) ;
    dffr ix42 (.Q (nx34), .QB (\$dummy [8]), .D (\input [3]), .CLK (NOT_clk), .R (
         nx216)) ;
    nor02_2x ix50 (.Y (nx49), .A0 (nx34), .A1 (nx182)) ;
    buf02 ix215 (.Y (nx216), .A (reset)) ;
endmodule


module saveState ( DMAOutput, RegisterOutput, bias1, bias2, bias3, bias4, bias5, 
                   bias6, bias7, bias8, Depth, NumberOfFiltersCounter, rst, 
                   stateinput, clk, outputCounterToDma, RealOutputCounter, 
                   \output , ShiftLeftCounterOutput, ShiftCounterRst, 
                   AddresCounterLoad, X, Y ) ;

    input [15:0]DMAOutput ;
    input [15:0]RegisterOutput ;
    input [15:0]bias1 ;
    input [15:0]bias2 ;
    input [15:0]bias3 ;
    input [15:0]bias4 ;
    input [15:0]bias5 ;
    input [15:0]bias6 ;
    input [15:0]bias7 ;
    input [15:0]bias8 ;
    input [3:0]Depth ;
    input [3:0]NumberOfFiltersCounter ;
    input rst ;
    input [14:0]stateinput ;
    input clk ;
    output [12:0]outputCounterToDma ;
    output [12:0]RealOutputCounter ;
    output [15:0]\output  ;
    output [4:0]ShiftLeftCounterOutput ;
    input ShiftCounterRst ;
    input [12:0]AddresCounterLoad ;
    input X ;
    input Y ;

    wire ShiftRegClk, resetCounter, Enable, GND0, nx238, nx240;



    Counter_5 Scounter (.enable (Enable), .reset (ShiftCounterRst), .clk (
              ShiftRegClk), .load (GND0), .\output  ({ShiftLeftCounterOutput[4],
              ShiftLeftCounterOutput[3],ShiftLeftCounterOutput[2],
              ShiftLeftCounterOutput[1],ShiftLeftCounterOutput[0]}), .\input  ({
              GND0,GND0,GND0,GND0,GND0})) ;
    addressCounter first (.reset (resetCounter), .current_state ({GND0,GND0,
                   stateinput[12],GND0,GND0,stateinput[9],nx238,GND0,GND0,GND0,
                   GND0,GND0,GND0,GND0,GND0}), .outputAddress ({
                   outputCounterToDma[12],outputCounterToDma[11],
                   outputCounterToDma[10],outputCounterToDma[9],
                   outputCounterToDma[8],outputCounterToDma[7],
                   outputCounterToDma[6],outputCounterToDma[5],
                   outputCounterToDma[4],outputCounterToDma[3],
                   outputCounterToDma[2],outputCounterToDma[1],
                   outputCounterToDma[0]}), .RealOutputCounter ({
                   RealOutputCounter[12],RealOutputCounter[11],
                   RealOutputCounter[10],RealOutputCounter[9],
                   RealOutputCounter[8],RealOutputCounter[7],
                   RealOutputCounter[6],RealOutputCounter[5],
                   RealOutputCounter[4],RealOutputCounter[3],
                   RealOutputCounter[2],RealOutputCounter[1],
                   RealOutputCounter[0]}), .AddresCounterLoad ({
                   AddresCounterLoad[12],AddresCounterLoad[11],
                   AddresCounterLoad[10],AddresCounterLoad[9],
                   AddresCounterLoad[8],AddresCounterLoad[7],
                   AddresCounterLoad[6],AddresCounterLoad[5],
                   AddresCounterLoad[4],AddresCounterLoad[3],
                   AddresCounterLoad[2],AddresCounterLoad[1],
                   AddresCounterLoad[0]}), .X (X), .Y (Y), .clk (clk)) ;
    depthNotZero second (.fromOutDMA ({DMAOutput[15],DMAOutput[14],DMAOutput[13]
                 ,DMAOutput[12],DMAOutput[11],DMAOutput[10],DMAOutput[9],
                 DMAOutput[8],DMAOutput[7],DMAOutput[6],DMAOutput[5],
                 DMAOutput[4],DMAOutput[3],DMAOutput[2],DMAOutput[1],
                 DMAOutput[0]}), .fromOutReg ({RegisterOutput[15],
                 RegisterOutput[14],RegisterOutput[13],RegisterOutput[12],
                 RegisterOutput[11],RegisterOutput[10],RegisterOutput[9],
                 RegisterOutput[8],RegisterOutput[7],RegisterOutput[6],
                 RegisterOutput[5],RegisterOutput[4],RegisterOutput[3],
                 RegisterOutput[2],RegisterOutput[1],RegisterOutput[0]}), .Depth (
                 {Depth[3],Depth[2],Depth[1],Depth[0]}), .current_state ({GND0,
                 GND0,GND0,GND0,GND0,GND0,nx238,GND0,GND0,GND0,GND0,GND0,GND0,
                 GND0,GND0}), .\output  ({\output [15],\output [14],\output [13]
                 ,\output [12],\output [11],\output [10],\output [9],\output [8]
                 ,\output [7],\output [6],\output [5],\output [4],\output [3],
                 \output [2],\output [1],\output [0]})) ;
    depthZero third (.fromOutReg ({RegisterOutput[15],RegisterOutput[14],
              RegisterOutput[13],RegisterOutput[12],RegisterOutput[11],
              RegisterOutput[10],RegisterOutput[9],RegisterOutput[8],
              RegisterOutput[7],RegisterOutput[6],RegisterOutput[5],
              RegisterOutput[4],RegisterOutput[3],RegisterOutput[2],
              RegisterOutput[1],RegisterOutput[0]}), .bias1 ({bias1[15],
              bias1[14],bias1[13],bias1[12],bias1[11],bias1[10],bias1[9],
              bias1[8],bias1[7],bias1[6],bias1[5],bias1[4],bias1[3],bias1[2],
              bias1[1],bias1[0]}), .bias2 ({bias2[15],bias2[14],bias2[13],
              bias2[12],bias2[11],bias2[10],bias2[9],bias2[8],bias2[7],bias2[6],
              bias2[5],bias2[4],bias2[3],bias2[2],bias2[1],bias2[0]}), .bias3 ({
              bias3[15],bias3[14],bias3[13],bias3[12],bias3[11],bias3[10],
              bias3[9],bias3[8],bias3[7],bias3[6],bias3[5],bias3[4],bias3[3],
              bias3[2],bias3[1],bias3[0]}), .bias4 ({bias4[15],bias4[14],
              bias4[13],bias4[12],bias4[11],bias4[10],bias4[9],bias4[8],bias4[7]
              ,bias4[6],bias4[5],bias4[4],bias4[3],bias4[2],bias4[1],bias4[0]})
              , .bias5 ({bias5[15],bias5[14],bias5[13],bias5[12],bias5[11],
              bias5[10],bias5[9],bias5[8],bias5[7],bias5[6],bias5[5],bias5[4],
              bias5[3],bias5[2],bias5[1],bias5[0]}), .bias6 ({bias6[15],
              bias6[14],bias6[13],bias6[12],bias6[11],bias6[10],bias6[9],
              bias6[8],bias6[7],bias6[6],bias6[5],bias6[4],bias6[3],bias6[2],
              bias6[1],bias6[0]}), .bias7 ({bias7[15],bias7[14],bias7[13],
              bias7[12],bias7[11],bias7[10],bias7[9],bias7[8],bias7[7],bias7[6],
              bias7[5],bias7[4],bias7[3],bias7[2],bias7[1],bias7[0]}), .bias8 ({
              bias8[15],bias8[14],bias8[13],bias8[12],bias8[11],bias8[10],
              bias8[9],bias8[8],bias8[7],bias8[6],bias8[5],bias8[4],bias8[3],
              bias8[2],bias8[1],bias8[0]}), .counterNumber ({
              NumberOfFiltersCounter[3],NumberOfFiltersCounter[2],
              NumberOfFiltersCounter[1],NumberOfFiltersCounter[0]}), .Depth ({
              Depth[3],Depth[2],Depth[1],Depth[0]}), .current_state ({GND0,GND0,
              GND0,GND0,GND0,GND0,nx238,GND0,GND0,GND0,GND0,GND0,GND0,GND0,GND0}
              ), .\output  ({\output [15],\output [14],\output [13],\output [12]
              ,\output [11],\output [10],\output [9],\output [8],\output [7],
              \output [6],\output [5],\output [4],\output [3],\output [2],
              \output [1],\output [0]})) ;
    fake_gnd ix214 (.Y (GND0)) ;
    or02 ix5 (.Y (Enable), .A0 (nx240), .A1 (stateinput[10])) ;
    or02 ix7 (.Y (resetCounter), .A0 (rst), .A1 (stateinput[13])) ;
    ao21 ix3 (.Y (ShiftRegClk), .A0 (clk), .A1 (stateinput[10]), .B0 (nx240)) ;
    buf02 ix237 (.Y (nx238), .A (stateinput[8])) ;
    buf02 ix239 (.Y (nx240), .A (stateinput[8])) ;
endmodule


module depthZero ( fromOutReg, bias1, bias2, bias3, bias4, bias5, bias6, bias7, 
                   bias8, counterNumber, Depth, current_state, \output  ) ;

    input [15:0]fromOutReg ;
    input [15:0]bias1 ;
    input [15:0]bias2 ;
    input [15:0]bias3 ;
    input [15:0]bias4 ;
    input [15:0]bias5 ;
    input [15:0]bias6 ;
    input [15:0]bias7 ;
    input [15:0]bias8 ;
    input [3:0]counterNumber ;
    input [3:0]Depth ;
    input [14:0]current_state ;
    output [15:0]\output  ;

    wire outputMux_15, outputMux_14, outputMux_13, outputMux_12, outputMux_11, 
         outputMux_10, outputMux_9, outputMux_8, outputMux_7, outputMux_6, 
         outputMux_5, outputMux_4, outputMux_3, outputMux_2, outputMux_1, 
         outputMux_0, outputAdder_15, outputAdder_14, outputAdder_13, 
         outputAdder_12, outputAdder_11, outputAdder_10, outputAdder_9, 
         outputAdder_8, outputAdder_7, outputAdder_6, outputAdder_5, 
         outputAdder_4, outputAdder_3, outputAdder_2, outputAdder_1, 
         outputAdder_0, Enable, GND, nx163, nx165;
    wire [0:0] \$dummy ;




    mux7 myMux (.a1 ({bias1[15],bias1[14],bias1[13],bias1[12],bias1[11],
         bias1[10],bias1[9],bias1[8],bias1[7],bias1[6],bias1[5],bias1[4],
         bias1[3],bias1[2],bias1[1],bias1[0]}), .a2 ({bias2[15],bias2[14],
         bias2[13],bias2[12],bias2[11],bias2[10],bias2[9],bias2[8],bias2[7],
         bias2[6],bias2[5],bias2[4],bias2[3],bias2[2],bias2[1],bias2[0]}), .a3 (
         {bias3[15],bias3[14],bias3[13],bias3[12],bias3[11],bias3[10],bias3[9],
         bias3[8],bias3[7],bias3[6],bias3[5],bias3[4],bias3[3],bias3[2],bias3[1]
         ,bias3[0]}), .a4 ({bias4[15],bias4[14],bias4[13],bias4[12],bias4[11],
         bias4[10],bias4[9],bias4[8],bias4[7],bias4[6],bias4[5],bias4[4],
         bias4[3],bias4[2],bias4[1],bias4[0]}), .a5 ({bias5[15],bias5[14],
         bias5[13],bias5[12],bias5[11],bias5[10],bias5[9],bias5[8],bias5[7],
         bias5[6],bias5[5],bias5[4],bias5[3],bias5[2],bias5[1],bias5[0]}), .a6 (
         {bias6[15],bias6[14],bias6[13],bias6[12],bias6[11],bias6[10],bias6[9],
         bias6[8],bias6[7],bias6[6],bias6[5],bias6[4],bias6[3],bias6[2],bias6[1]
         ,bias6[0]}), .a7 ({bias7[15],bias7[14],bias7[13],bias7[12],bias7[11],
         bias7[10],bias7[9],bias7[8],bias7[7],bias7[6],bias7[5],bias7[4],
         bias7[3],bias7[2],bias7[1],bias7[0]}), .a8 ({bias8[15],bias8[14],
         bias8[13],bias8[12],bias8[11],bias8[10],bias8[9],bias8[8],bias8[7],
         bias8[6],bias8[5],bias8[4],bias8[3],bias8[2],bias8[1],bias8[0]}), .sel (
         {counterNumber[3],counterNumber[2],counterNumber[1],counterNumber[0]})
         , .\output  ({outputMux_15,outputMux_14,outputMux_13,outputMux_12,
         outputMux_11,outputMux_10,outputMux_9,outputMux_8,outputMux_7,
         outputMux_6,outputMux_5,outputMux_4,outputMux_3,outputMux_2,outputMux_1
         ,outputMux_0})) ;
    my_nadder_16 myNadder (.a ({fromOutReg[15],fromOutReg[14],fromOutReg[13],
                 fromOutReg[12],fromOutReg[11],fromOutReg[10],fromOutReg[9],
                 fromOutReg[8],fromOutReg[7],fromOutReg[6],fromOutReg[5],
                 fromOutReg[4],fromOutReg[3],fromOutReg[2],fromOutReg[1],
                 fromOutReg[0]}), .b ({outputMux_15,outputMux_14,outputMux_13,
                 outputMux_12,outputMux_11,outputMux_10,outputMux_9,outputMux_8,
                 outputMux_7,outputMux_6,outputMux_5,outputMux_4,outputMux_3,
                 outputMux_2,outputMux_1,outputMux_0}), .cin (GND), .s ({
                 outputAdder_15,outputAdder_14,outputAdder_13,outputAdder_12,
                 outputAdder_11,outputAdder_10,outputAdder_9,outputAdder_8,
                 outputAdder_7,outputAdder_6,outputAdder_5,outputAdder_4,
                 outputAdder_3,outputAdder_2,outputAdder_1,outputAdder_0}), .cout (
                 \$dummy [0])) ;
    triStateBuffer_16 depth0 (.D ({outputAdder_15,outputAdder_14,outputAdder_13,
                      outputAdder_12,outputAdder_11,outputAdder_10,outputAdder_9
                      ,outputAdder_8,outputAdder_7,outputAdder_6,outputAdder_5,
                      outputAdder_4,outputAdder_3,outputAdder_2,outputAdder_1,
                      outputAdder_0}), .EN (Enable), .F ({\output [15],
                      \output [14],\output [13],\output [12],\output [11],
                      \output [10],\output [9],\output [8],\output [7],
                      \output [6],\output [5],\output [4],\output [3],
                      \output [2],\output [1],\output [0]})) ;
    fake_gnd ix150 (.Y (GND)) ;
    nor04 ix15 (.Y (Enable), .A0 (Depth[1]), .A1 (Depth[3]), .A2 (Depth[2]), .A3 (
          nx163)) ;
    nand02 ix164 (.Y (nx163), .A0 (nx165), .A1 (current_state[8])) ;
    inv01 ix166 (.Y (nx165), .A (Depth[0])) ;
endmodule


module mux7 ( a1, a2, a3, a4, a5, a6, a7, a8, sel, \output  ) ;

    input [15:0]a1 ;
    input [15:0]a2 ;
    input [15:0]a3 ;
    input [15:0]a4 ;
    input [15:0]a5 ;
    input [15:0]a6 ;
    input [15:0]a7 ;
    input [15:0]a8 ;
    input [3:0]sel ;
    output [15:0]\output  ;

    wire nx12, nx18, nx80, nx217, nx221, nx223, nx227, nx231, nx233, nx239, 
         nx241, nx247, nx255, nx257, nx259, nx261, nx265, nx267, nx269, nx271, 
         nx275, nx277, nx279, nx281, nx285, nx287, nx289, nx291, nx295, nx297, 
         nx299, nx301, nx305, nx307, nx309, nx311, nx315, nx317, nx319, nx321, 
         nx325, nx327, nx329, nx331, nx335, nx337, nx339, nx341, nx345, nx347, 
         nx349, nx351, nx355, nx357, nx359, nx361, nx365, nx367, nx369, nx371, 
         nx375, nx377, nx379, nx381, nx385, nx387, nx389, nx391, nx395, nx397, 
         nx399, nx401, nx408, nx410, nx412, nx414, nx416, nx418, nx421, nx423, 
         nx425, nx427, nx429, nx431, nx433, nx435, nx437, nx439, nx441, nx443, 
         nx445, nx447, nx449, nx451, nx453, nx455, nx457, nx459, nx461, nx463, 
         nx465, nx467;



    nand04 ix89 (.Y (\output [0]), .A0 (nx217), .A1 (nx233), .A2 (nx241), .A3 (
           nx247)) ;
    aoi22 ix218 (.Y (nx217), .A0 (a7[0]), .A1 (nx459), .B0 (a8[0]), .B1 (nx465)
          ) ;
    inv01 ix222 (.Y (nx221), .A (sel[2])) ;
    inv01 ix224 (.Y (nx223), .A (sel[1])) ;
    nand02 ix81 (.Y (nx80), .A0 (nx227), .A1 (nx231)) ;
    nand03 ix228 (.Y (nx227), .A0 (nx18), .A1 (sel[2]), .A2 (sel[1])) ;
    nor02ii ix19 (.Y (nx18), .A0 (sel[3]), .A1 (sel[0])) ;
    inv01 ix232 (.Y (nx231), .A (sel[3])) ;
    aoi22 ix234 (.Y (nx233), .A0 (a3[0]), .A1 (nx451), .B0 (a2[0]), .B1 (nx443)
          ) ;
    aoi22 ix242 (.Y (nx241), .A0 (a5[0]), .A1 (nx435), .B0 (a6[0]), .B1 (nx427)
          ) ;
    aoi22 ix248 (.Y (nx247), .A0 (a1[0]), .A1 (nx410), .B0 (a4[0]), .B1 (nx418)
          ) ;
    nor04 ix13 (.Y (nx12), .A0 (sel[3]), .A1 (sel[0]), .A2 (sel[2]), .A3 (sel[1]
          )) ;
    nand04 ix119 (.Y (\output [1]), .A0 (nx255), .A1 (nx257), .A2 (nx259), .A3 (
           nx261)) ;
    aoi22 ix256 (.Y (nx255), .A0 (a7[1]), .A1 (nx459), .B0 (a8[1]), .B1 (nx465)
          ) ;
    aoi22 ix258 (.Y (nx257), .A0 (a3[1]), .A1 (nx451), .B0 (a2[1]), .B1 (nx443)
          ) ;
    aoi22 ix260 (.Y (nx259), .A0 (a5[1]), .A1 (nx435), .B0 (a6[1]), .B1 (nx427)
          ) ;
    aoi22 ix262 (.Y (nx261), .A0 (a1[1]), .A1 (nx410), .B0 (a4[1]), .B1 (nx418)
          ) ;
    nand04 ix149 (.Y (\output [2]), .A0 (nx265), .A1 (nx267), .A2 (nx269), .A3 (
           nx271)) ;
    aoi22 ix266 (.Y (nx265), .A0 (a7[2]), .A1 (nx459), .B0 (a8[2]), .B1 (nx465)
          ) ;
    aoi22 ix268 (.Y (nx267), .A0 (a3[2]), .A1 (nx451), .B0 (a2[2]), .B1 (nx443)
          ) ;
    aoi22 ix270 (.Y (nx269), .A0 (a5[2]), .A1 (nx435), .B0 (a6[2]), .B1 (nx427)
          ) ;
    aoi22 ix272 (.Y (nx271), .A0 (a1[2]), .A1 (nx410), .B0 (a4[2]), .B1 (nx418)
          ) ;
    nand04 ix179 (.Y (\output [3]), .A0 (nx275), .A1 (nx277), .A2 (nx279), .A3 (
           nx281)) ;
    aoi22 ix276 (.Y (nx275), .A0 (a7[3]), .A1 (nx459), .B0 (a8[3]), .B1 (nx465)
          ) ;
    aoi22 ix278 (.Y (nx277), .A0 (a3[3]), .A1 (nx451), .B0 (a2[3]), .B1 (nx443)
          ) ;
    aoi22 ix280 (.Y (nx279), .A0 (a5[3]), .A1 (nx435), .B0 (a6[3]), .B1 (nx427)
          ) ;
    aoi22 ix282 (.Y (nx281), .A0 (a1[3]), .A1 (nx410), .B0 (a4[3]), .B1 (nx418)
          ) ;
    nand04 ix209 (.Y (\output [4]), .A0 (nx285), .A1 (nx287), .A2 (nx289), .A3 (
           nx291)) ;
    aoi22 ix286 (.Y (nx285), .A0 (a7[4]), .A1 (nx459), .B0 (a8[4]), .B1 (nx465)
          ) ;
    aoi22 ix288 (.Y (nx287), .A0 (a3[4]), .A1 (nx451), .B0 (a2[4]), .B1 (nx443)
          ) ;
    aoi22 ix290 (.Y (nx289), .A0 (a5[4]), .A1 (nx435), .B0 (a6[4]), .B1 (nx427)
          ) ;
    aoi22 ix292 (.Y (nx291), .A0 (a1[4]), .A1 (nx410), .B0 (a4[4]), .B1 (nx418)
          ) ;
    nand04 ix239 (.Y (\output [5]), .A0 (nx295), .A1 (nx297), .A2 (nx299), .A3 (
           nx301)) ;
    aoi22 ix296 (.Y (nx295), .A0 (a7[5]), .A1 (nx459), .B0 (a8[5]), .B1 (nx465)
          ) ;
    aoi22 ix298 (.Y (nx297), .A0 (a3[5]), .A1 (nx451), .B0 (a2[5]), .B1 (nx443)
          ) ;
    aoi22 ix300 (.Y (nx299), .A0 (a5[5]), .A1 (nx435), .B0 (a6[5]), .B1 (nx427)
          ) ;
    aoi22 ix302 (.Y (nx301), .A0 (a1[5]), .A1 (nx410), .B0 (a4[5]), .B1 (nx418)
          ) ;
    nand04 ix269 (.Y (\output [6]), .A0 (nx305), .A1 (nx307), .A2 (nx309), .A3 (
           nx311)) ;
    aoi22 ix306 (.Y (nx305), .A0 (a7[6]), .A1 (nx459), .B0 (a8[6]), .B1 (nx465)
          ) ;
    aoi22 ix308 (.Y (nx307), .A0 (a3[6]), .A1 (nx451), .B0 (a2[6]), .B1 (nx443)
          ) ;
    aoi22 ix310 (.Y (nx309), .A0 (a5[6]), .A1 (nx435), .B0 (a6[6]), .B1 (nx427)
          ) ;
    aoi22 ix312 (.Y (nx311), .A0 (a1[6]), .A1 (nx410), .B0 (a4[6]), .B1 (nx418)
          ) ;
    nand04 ix299 (.Y (\output [7]), .A0 (nx315), .A1 (nx317), .A2 (nx319), .A3 (
           nx321)) ;
    aoi22 ix316 (.Y (nx315), .A0 (a7[7]), .A1 (nx461), .B0 (a8[7]), .B1 (nx467)
          ) ;
    aoi22 ix318 (.Y (nx317), .A0 (a3[7]), .A1 (nx453), .B0 (a2[7]), .B1 (nx445)
          ) ;
    aoi22 ix320 (.Y (nx319), .A0 (a5[7]), .A1 (nx437), .B0 (a6[7]), .B1 (nx429)
          ) ;
    aoi22 ix322 (.Y (nx321), .A0 (a1[7]), .A1 (nx412), .B0 (a4[7]), .B1 (nx421)
          ) ;
    nand04 ix329 (.Y (\output [8]), .A0 (nx325), .A1 (nx327), .A2 (nx329), .A3 (
           nx331)) ;
    aoi22 ix326 (.Y (nx325), .A0 (a7[8]), .A1 (nx461), .B0 (a8[8]), .B1 (nx467)
          ) ;
    aoi22 ix328 (.Y (nx327), .A0 (a3[8]), .A1 (nx453), .B0 (a2[8]), .B1 (nx445)
          ) ;
    aoi22 ix330 (.Y (nx329), .A0 (a5[8]), .A1 (nx437), .B0 (a6[8]), .B1 (nx429)
          ) ;
    aoi22 ix332 (.Y (nx331), .A0 (a1[8]), .A1 (nx412), .B0 (a4[8]), .B1 (nx421)
          ) ;
    nand04 ix359 (.Y (\output [9]), .A0 (nx335), .A1 (nx337), .A2 (nx339), .A3 (
           nx341)) ;
    aoi22 ix336 (.Y (nx335), .A0 (a7[9]), .A1 (nx461), .B0 (a8[9]), .B1 (nx467)
          ) ;
    aoi22 ix338 (.Y (nx337), .A0 (a3[9]), .A1 (nx453), .B0 (a2[9]), .B1 (nx445)
          ) ;
    aoi22 ix340 (.Y (nx339), .A0 (a5[9]), .A1 (nx437), .B0 (a6[9]), .B1 (nx429)
          ) ;
    aoi22 ix342 (.Y (nx341), .A0 (a1[9]), .A1 (nx412), .B0 (a4[9]), .B1 (nx421)
          ) ;
    nand04 ix389 (.Y (\output [10]), .A0 (nx345), .A1 (nx347), .A2 (nx349), .A3 (
           nx351)) ;
    aoi22 ix346 (.Y (nx345), .A0 (a7[10]), .A1 (nx461), .B0 (a8[10]), .B1 (nx467
          )) ;
    aoi22 ix348 (.Y (nx347), .A0 (a3[10]), .A1 (nx453), .B0 (a2[10]), .B1 (nx445
          )) ;
    aoi22 ix350 (.Y (nx349), .A0 (a5[10]), .A1 (nx437), .B0 (a6[10]), .B1 (nx429
          )) ;
    aoi22 ix352 (.Y (nx351), .A0 (a1[10]), .A1 (nx412), .B0 (a4[10]), .B1 (nx421
          )) ;
    nand04 ix419 (.Y (\output [11]), .A0 (nx355), .A1 (nx357), .A2 (nx359), .A3 (
           nx361)) ;
    aoi22 ix356 (.Y (nx355), .A0 (a7[11]), .A1 (nx461), .B0 (a8[11]), .B1 (nx467
          )) ;
    aoi22 ix358 (.Y (nx357), .A0 (a3[11]), .A1 (nx453), .B0 (a2[11]), .B1 (nx445
          )) ;
    aoi22 ix360 (.Y (nx359), .A0 (a5[11]), .A1 (nx437), .B0 (a6[11]), .B1 (nx429
          )) ;
    aoi22 ix362 (.Y (nx361), .A0 (a1[11]), .A1 (nx412), .B0 (a4[11]), .B1 (nx421
          )) ;
    nand04 ix449 (.Y (\output [12]), .A0 (nx365), .A1 (nx367), .A2 (nx369), .A3 (
           nx371)) ;
    aoi22 ix366 (.Y (nx365), .A0 (a7[12]), .A1 (nx461), .B0 (a8[12]), .B1 (nx467
          )) ;
    aoi22 ix368 (.Y (nx367), .A0 (a3[12]), .A1 (nx453), .B0 (a2[12]), .B1 (nx445
          )) ;
    aoi22 ix370 (.Y (nx369), .A0 (a5[12]), .A1 (nx437), .B0 (a6[12]), .B1 (nx429
          )) ;
    aoi22 ix372 (.Y (nx371), .A0 (a1[12]), .A1 (nx412), .B0 (a4[12]), .B1 (nx421
          )) ;
    nand04 ix479 (.Y (\output [13]), .A0 (nx375), .A1 (nx377), .A2 (nx379), .A3 (
           nx381)) ;
    aoi22 ix376 (.Y (nx375), .A0 (a7[13]), .A1 (nx461), .B0 (a8[13]), .B1 (nx467
          )) ;
    aoi22 ix378 (.Y (nx377), .A0 (a3[13]), .A1 (nx453), .B0 (a2[13]), .B1 (nx445
          )) ;
    aoi22 ix380 (.Y (nx379), .A0 (a5[13]), .A1 (nx437), .B0 (a6[13]), .B1 (nx429
          )) ;
    aoi22 ix382 (.Y (nx381), .A0 (a1[13]), .A1 (nx412), .B0 (a4[13]), .B1 (nx421
          )) ;
    nand04 ix509 (.Y (\output [14]), .A0 (nx385), .A1 (nx387), .A2 (nx389), .A3 (
           nx391)) ;
    aoi22 ix386 (.Y (nx385), .A0 (a7[14]), .A1 (nx463), .B0 (a8[14]), .B1 (nx80)
          ) ;
    aoi22 ix388 (.Y (nx387), .A0 (a3[14]), .A1 (nx455), .B0 (a2[14]), .B1 (nx447
          )) ;
    aoi22 ix390 (.Y (nx389), .A0 (a5[14]), .A1 (nx439), .B0 (a6[14]), .B1 (nx431
          )) ;
    aoi22 ix392 (.Y (nx391), .A0 (a1[14]), .A1 (nx414), .B0 (a4[14]), .B1 (nx423
          )) ;
    nand04 ix539 (.Y (\output [15]), .A0 (nx395), .A1 (nx397), .A2 (nx399), .A3 (
           nx401)) ;
    aoi22 ix396 (.Y (nx395), .A0 (a7[15]), .A1 (nx463), .B0 (a8[15]), .B1 (nx80)
          ) ;
    aoi22 ix398 (.Y (nx397), .A0 (a3[15]), .A1 (nx455), .B0 (a2[15]), .B1 (nx447
          )) ;
    aoi22 ix400 (.Y (nx399), .A0 (a5[15]), .A1 (nx439), .B0 (a6[15]), .B1 (nx431
          )) ;
    aoi22 ix402 (.Y (nx401), .A0 (a1[15]), .A1 (nx414), .B0 (a4[15]), .B1 (nx423
          )) ;
    inv01 ix240 (.Y (nx239), .A (nx18)) ;
    inv01 ix407 (.Y (nx408), .A (nx12)) ;
    inv02 ix409 (.Y (nx410), .A (nx408)) ;
    inv02 ix411 (.Y (nx412), .A (nx408)) ;
    inv02 ix413 (.Y (nx414), .A (nx408)) ;
    inv02 ix417 (.Y (nx418), .A (nx416)) ;
    inv02 ix420 (.Y (nx421), .A (nx416)) ;
    inv02 ix422 (.Y (nx423), .A (nx416)) ;
    inv02 ix426 (.Y (nx427), .A (nx425)) ;
    inv02 ix428 (.Y (nx429), .A (nx425)) ;
    inv02 ix430 (.Y (nx431), .A (nx425)) ;
    inv02 ix434 (.Y (nx435), .A (nx433)) ;
    inv02 ix436 (.Y (nx437), .A (nx433)) ;
    inv02 ix438 (.Y (nx439), .A (nx433)) ;
    inv02 ix442 (.Y (nx443), .A (nx441)) ;
    inv02 ix444 (.Y (nx445), .A (nx441)) ;
    inv02 ix446 (.Y (nx447), .A (nx441)) ;
    inv02 ix450 (.Y (nx451), .A (nx449)) ;
    inv02 ix452 (.Y (nx453), .A (nx449)) ;
    inv02 ix454 (.Y (nx455), .A (nx449)) ;
    inv02 ix458 (.Y (nx459), .A (nx457)) ;
    inv02 ix460 (.Y (nx461), .A (nx457)) ;
    inv02 ix462 (.Y (nx463), .A (nx457)) ;
    nand02 ix464 (.Y (nx465), .A0 (nx227), .A1 (nx231)) ;
    nand02 ix466 (.Y (nx467), .A0 (nx227), .A1 (nx231)) ;
    or04 ix73 (.Y (nx457), .A0 (sel[3]), .A1 (sel[0]), .A2 (nx221), .A3 (nx223)
         ) ;
    or04 ix68 (.Y (nx449), .A0 (sel[3]), .A1 (sel[0]), .A2 (sel[2]), .A3 (nx223)
         ) ;
    or03 ix57 (.Y (nx441), .A0 (nx239), .A1 (sel[2]), .A2 (sel[1])) ;
    or04 ix43 (.Y (nx433), .A0 (sel[3]), .A1 (sel[0]), .A2 (nx221), .A3 (sel[1])
         ) ;
    nand03 ix35 (.Y (nx425), .A0 (nx18), .A1 (sel[2]), .A2 (nx223)) ;
    nand03 ix25 (.Y (nx416), .A0 (nx18), .A1 (nx221), .A2 (sel[1])) ;
endmodule


module depthNotZero ( fromOutDMA, fromOutReg, Depth, current_state, \output  ) ;

    input [15:0]fromOutDMA ;
    input [15:0]fromOutReg ;
    input [3:0]Depth ;
    input [14:0]current_state ;
    output [15:0]\output  ;

    wire outputAdder_15, outputAdder_14, outputAdder_13, outputAdder_12, 
         outputAdder_11, outputAdder_10, outputAdder_9, outputAdder_8, 
         outputAdder_7, outputAdder_6, outputAdder_5, outputAdder_4, 
         outputAdder_3, outputAdder_2, outputAdder_1, outputAdder_0, Enable, GND, 
         nx117;
    wire [0:0] \$dummy ;




    my_nadder_16 myNadder (.a ({fromOutReg[15],fromOutReg[14],fromOutReg[13],
                 fromOutReg[12],fromOutReg[11],fromOutReg[10],fromOutReg[9],
                 fromOutReg[8],fromOutReg[7],fromOutReg[6],fromOutReg[5],
                 fromOutReg[4],fromOutReg[3],fromOutReg[2],fromOutReg[1],
                 fromOutReg[0]}), .b ({fromOutDMA[15],fromOutDMA[14],
                 fromOutDMA[13],fromOutDMA[12],fromOutDMA[11],fromOutDMA[10],
                 fromOutDMA[9],fromOutDMA[8],fromOutDMA[7],fromOutDMA[6],
                 fromOutDMA[5],fromOutDMA[4],fromOutDMA[3],fromOutDMA[2],
                 fromOutDMA[1],fromOutDMA[0]}), .cin (GND), .s ({outputAdder_15,
                 outputAdder_14,outputAdder_13,outputAdder_12,outputAdder_11,
                 outputAdder_10,outputAdder_9,outputAdder_8,outputAdder_7,
                 outputAdder_6,outputAdder_5,outputAdder_4,outputAdder_3,
                 outputAdder_2,outputAdder_1,outputAdder_0}), .cout (\$dummy [0]
                 )) ;
    triStateBuffer_16 depth0 (.D ({outputAdder_15,outputAdder_14,outputAdder_13,
                      outputAdder_12,outputAdder_11,outputAdder_10,outputAdder_9
                      ,outputAdder_8,outputAdder_7,outputAdder_6,outputAdder_5,
                      outputAdder_4,outputAdder_3,outputAdder_2,outputAdder_1,
                      outputAdder_0}), .EN (Enable), .F ({\output [15],
                      \output [14],\output [13],\output [12],\output [11],
                      \output [10],\output [9],\output [8],\output [7],
                      \output [6],\output [5],\output [4],\output [3],
                      \output [2],\output [1],\output [0]})) ;
    fake_gnd ix104 (.Y (GND)) ;
    nor02ii ix7 (.Y (Enable), .A0 (nx117), .A1 (current_state[8])) ;
    nor04 ix118 (.Y (nx117), .A0 (Depth[0]), .A1 (Depth[1]), .A2 (Depth[2]), .A3 (
          Depth[3])) ;
endmodule


module addressCounter ( reset, current_state, outputAddress, RealOutputCounter, 
                        AddresCounterLoad, X, Y, clk ) ;

    input reset ;
    input [14:0]current_state ;
    output [12:0]outputAddress ;
    output [12:0]RealOutputCounter ;
    input [12:0]AddresCounterLoad ;
    input X ;
    input Y ;
    input clk ;

    wire CounterClk, CounterRest, Load, nx110;



    Counter_13 myCounter (.enable (current_state[8]), .reset (CounterRest), .clk (
               CounterClk), .load (Load), .\output  ({RealOutputCounter[12],
               RealOutputCounter[11],RealOutputCounter[10],RealOutputCounter[9],
               RealOutputCounter[8],RealOutputCounter[7],RealOutputCounter[6],
               RealOutputCounter[5],RealOutputCounter[4],RealOutputCounter[3],
               RealOutputCounter[2],RealOutputCounter[1],RealOutputCounter[0]})
               , .\input  ({AddresCounterLoad[12],AddresCounterLoad[11],
               AddresCounterLoad[10],AddresCounterLoad[9],AddresCounterLoad[8],
               AddresCounterLoad[7],AddresCounterLoad[6],AddresCounterLoad[5],
               AddresCounterLoad[4],AddresCounterLoad[3],AddresCounterLoad[2],
               AddresCounterLoad[1],AddresCounterLoad[0]})) ;
    triStateBuffer_13 outOfAddressCounter (.D ({RealOutputCounter[12],
                      RealOutputCounter[11],RealOutputCounter[10],
                      RealOutputCounter[9],RealOutputCounter[8],
                      RealOutputCounter[7],RealOutputCounter[6],
                      RealOutputCounter[5],RealOutputCounter[4],
                      RealOutputCounter[3],RealOutputCounter[2],
                      RealOutputCounter[1],RealOutputCounter[0]}), .EN (
                      current_state[8]), .F ({outputAddress[12],
                      outputAddress[11],outputAddress[10],outputAddress[9],
                      outputAddress[8],outputAddress[7],outputAddress[6],
                      outputAddress[5],outputAddress[4],outputAddress[3],
                      outputAddress[2],outputAddress[1],outputAddress[0]})) ;
    aoi21 ix11 (.Y (Load), .A0 (X), .A1 (Y), .B0 (nx110)) ;
    inv01 ix111 (.Y (nx110), .A (current_state[9])) ;
    or02 ix13 (.Y (CounterRest), .A0 (reset), .A1 (current_state[12])) ;
    ao21 ix3 (.Y (CounterClk), .A0 (clk), .A1 (current_state[9]), .B0 (
         current_state[8])) ;
endmodule


module Counter_13 ( enable, reset, clk, load, \output , \input  ) ;

    input enable ;
    input reset ;
    input clk ;
    input load ;
    output [12:0]\output  ;
    input [12:0]\input  ;

    wire addResult_12, addResult_11, addResult_10, addResult_9, addResult_8, 
         addResult_7, addResult_6, addResult_5, addResult_4, addResult_3, 
         addResult_2, addResult_1, addResult_0, one_0, one_12, nx160, nx8, nx12, 
         nx154, nx20, nx24, nx148, nx32, nx36, nx142, nx44, nx48, nx136, nx56, 
         nx60, nx130, nx68, nx72, nx124, nx80, nx84, nx118, nx92, nx96, nx112, 
         nx104, nx108, nx106, nx117, nx121, nx100, nx129, nx133, nx94, nx141, 
         nx145, nx88, nx153, nx157, nx404, nx414, nx424, nx434, nx444, nx454, 
         nx464, nx474, nx484, nx494, nx504, nx514, nx524, nx533, nx630, nx632, 
         nx634, nx648, nx650, nx652, nx654, nx656, nx658, nx660, nx662, nx664, 
         nx666, nx668;
    wire [26:0] \$dummy ;




    my_nadder_13 A1 (.a ({\output [12],\output [11],\output [10],\output [9],
                 \output [8],\output [7],\output [6],\output [5],\output [4],
                 \output [3],\output [2],\output [1],\output [0]}), .b ({one_12,
                 one_12,one_12,one_12,one_12,one_12,one_12,one_12,one_12,one_12,
                 one_12,one_12,one_0}), .cin (one_12), .s ({addResult_12,
                 addResult_11,addResult_10,addResult_9,addResult_8,addResult_7,
                 addResult_6,addResult_5,addResult_4,addResult_3,addResult_2,
                 addResult_1,addResult_0}), .cout (\$dummy [0])) ;
    fake_gnd ix354 (.Y (one_12)) ;
    fake_vcc ix352 (.Y (one_0)) ;
    dffsr_ni reg_toOutput_0__dup_1 (.Q (\output [0]), .QB (\$dummy [1]), .D (
             nx404), .CLK (nx648), .S (nx8), .R (nx12)) ;
    mux21_ni ix405 (.Y (nx404), .A0 (\output [0]), .A1 (addResult_0), .S0 (nx658
             )) ;
    nor02_2x ix534 (.Y (nx533), .A0 (nx654), .A1 (load)) ;
    dffr ix161 (.Q (nx160), .QB (\$dummy [2]), .D (\input [0]), .CLK (nx662), .R (
         nx654)) ;
    dffsr_ni reg_toOutput_1__dup_1 (.Q (\output [1]), .QB (\$dummy [3]), .D (
             nx414), .CLK (nx648), .S (nx20), .R (nx24)) ;
    mux21_ni ix415 (.Y (nx414), .A0 (\output [1]), .A1 (addResult_1), .S0 (nx658
             )) ;
    dffr ix155 (.Q (nx154), .QB (\$dummy [4]), .D (\input [1]), .CLK (nx662), .R (
         nx654)) ;
    dffsr_ni reg_toOutput_2__dup_1 (.Q (\output [2]), .QB (\$dummy [5]), .D (
             nx424), .CLK (nx648), .S (nx32), .R (nx36)) ;
    mux21_ni ix425 (.Y (nx424), .A0 (\output [2]), .A1 (addResult_2), .S0 (nx658
             )) ;
    dffr ix149 (.Q (nx148), .QB (\$dummy [6]), .D (\input [2]), .CLK (nx662), .R (
         nx654)) ;
    dffsr_ni reg_toOutput_3__dup_1 (.Q (\output [3]), .QB (\$dummy [7]), .D (
             nx434), .CLK (nx648), .S (nx44), .R (nx48)) ;
    mux21_ni ix435 (.Y (nx434), .A0 (\output [3]), .A1 (addResult_3), .S0 (nx658
             )) ;
    dffr ix143 (.Q (nx142), .QB (\$dummy [8]), .D (\input [3]), .CLK (nx662), .R (
         nx654)) ;
    dffsr_ni reg_toOutput_4__dup_1 (.Q (\output [4]), .QB (\$dummy [9]), .D (
             nx444), .CLK (nx648), .S (nx56), .R (nx60)) ;
    mux21_ni ix445 (.Y (nx444), .A0 (\output [4]), .A1 (addResult_4), .S0 (nx658
             )) ;
    dffr ix137 (.Q (nx136), .QB (\$dummy [10]), .D (\input [4]), .CLK (nx662), .R (
         nx654)) ;
    dffsr_ni reg_toOutput_5__dup_1 (.Q (\output [5]), .QB (\$dummy [11]), .D (
             nx454), .CLK (nx650), .S (nx68), .R (nx72)) ;
    mux21_ni ix455 (.Y (nx454), .A0 (\output [5]), .A1 (addResult_5), .S0 (nx658
             )) ;
    dffr ix131 (.Q (nx130), .QB (\$dummy [12]), .D (\input [5]), .CLK (nx662), .R (
         nx654)) ;
    dffsr_ni reg_toOutput_6__dup_1 (.Q (\output [6]), .QB (\$dummy [13]), .D (
             nx464), .CLK (nx650), .S (nx80), .R (nx84)) ;
    mux21_ni ix465 (.Y (nx464), .A0 (\output [6]), .A1 (addResult_6), .S0 (nx658
             )) ;
    dffr ix125 (.Q (nx124), .QB (\$dummy [14]), .D (\input [6]), .CLK (nx662), .R (
         nx656)) ;
    dffsr_ni reg_toOutput_7__dup_1 (.Q (\output [7]), .QB (\$dummy [15]), .D (
             nx474), .CLK (nx650), .S (nx92), .R (nx96)) ;
    mux21_ni ix475 (.Y (nx474), .A0 (\output [7]), .A1 (addResult_7), .S0 (nx660
             )) ;
    dffr ix119 (.Q (nx118), .QB (\$dummy [16]), .D (\input [7]), .CLK (nx632), .R (
         nx656)) ;
    dffsr_ni reg_toOutput_8__dup_1 (.Q (\output [8]), .QB (\$dummy [17]), .D (
             nx484), .CLK (nx650), .S (nx104), .R (nx108)) ;
    mux21_ni ix485 (.Y (nx484), .A0 (\output [8]), .A1 (addResult_8), .S0 (nx660
             )) ;
    dffr ix113 (.Q (nx112), .QB (\$dummy [18]), .D (\input [8]), .CLK (nx632), .R (
         nx656)) ;
    dffsr_ni reg_toOutput_9__dup_1 (.Q (\output [9]), .QB (\$dummy [19]), .D (
             nx494), .CLK (nx650), .S (nx117), .R (nx121)) ;
    mux21_ni ix495 (.Y (nx494), .A0 (\output [9]), .A1 (addResult_9), .S0 (nx660
             )) ;
    dffr ix114 (.Q (nx106), .QB (\$dummy [20]), .D (\input [9]), .CLK (nx632), .R (
         nx656)) ;
    dffsr_ni reg_toOutput_10__dup_1 (.Q (\output [10]), .QB (\$dummy [21]), .D (
             nx504), .CLK (nx652), .S (nx129), .R (nx133)) ;
    mux21_ni ix505 (.Y (nx504), .A0 (\output [10]), .A1 (addResult_10), .S0 (
             nx660)) ;
    dffr ix126 (.Q (nx100), .QB (\$dummy [22]), .D (\input [10]), .CLK (nx632), 
         .R (nx656)) ;
    dffsr_ni reg_toOutput_11__dup_1 (.Q (\output [11]), .QB (\$dummy [23]), .D (
             nx514), .CLK (nx652), .S (nx141), .R (nx145)) ;
    mux21_ni ix515 (.Y (nx514), .A0 (\output [11]), .A1 (addResult_11), .S0 (
             nx660)) ;
    dffr ix138 (.Q (nx94), .QB (\$dummy [24]), .D (\input [11]), .CLK (nx632), .R (
         nx656)) ;
    dffsr_ni reg_toOutput_12__dup_1 (.Q (\output [12]), .QB (\$dummy [25]), .D (
             nx524), .CLK (nx652), .S (nx153), .R (nx157)) ;
    mux21_ni ix525 (.Y (nx524), .A0 (\output [12]), .A1 (addResult_12), .S0 (
             nx660)) ;
    dffr ix150 (.Q (nx88), .QB (\$dummy [26]), .D (\input [12]), .CLK (nx632), .R (
         nx656)) ;
    inv02 ix629 (.Y (nx630), .A (clk)) ;
    inv02 ix631 (.Y (nx632), .A (nx652)) ;
    inv01 ix633 (.Y (nx634), .A (nx533)) ;
    and02 ix9 (.Y (nx8), .A0 (nx664), .A1 (nx160)) ;
    nor02ii ix13 (.Y (nx12), .A0 (nx160), .A1 (nx664)) ;
    and02 ix21 (.Y (nx20), .A0 (nx664), .A1 (nx154)) ;
    nor02ii ix25 (.Y (nx24), .A0 (nx154), .A1 (nx664)) ;
    and02 ix33 (.Y (nx32), .A0 (nx664), .A1 (nx148)) ;
    nor02ii ix37 (.Y (nx36), .A0 (nx148), .A1 (nx664)) ;
    and02 ix45 (.Y (nx44), .A0 (nx664), .A1 (nx142)) ;
    nor02ii ix49 (.Y (nx48), .A0 (nx142), .A1 (nx666)) ;
    and02 ix57 (.Y (nx56), .A0 (nx666), .A1 (nx136)) ;
    nor02ii ix61 (.Y (nx60), .A0 (nx136), .A1 (nx666)) ;
    and02 ix69 (.Y (nx68), .A0 (nx666), .A1 (nx130)) ;
    nor02ii ix73 (.Y (nx72), .A0 (nx130), .A1 (nx666)) ;
    and02 ix81 (.Y (nx80), .A0 (nx666), .A1 (nx124)) ;
    nor02ii ix85 (.Y (nx84), .A0 (nx124), .A1 (nx666)) ;
    and02 ix93 (.Y (nx92), .A0 (nx668), .A1 (nx118)) ;
    nor02ii ix97 (.Y (nx96), .A0 (nx118), .A1 (nx668)) ;
    and02 ix105 (.Y (nx104), .A0 (nx668), .A1 (nx112)) ;
    nor02ii ix109 (.Y (nx108), .A0 (nx112), .A1 (nx668)) ;
    and02 ix118 (.Y (nx117), .A0 (nx668), .A1 (nx106)) ;
    nor02ii ix122 (.Y (nx121), .A0 (nx106), .A1 (nx668)) ;
    and02 ix130 (.Y (nx129), .A0 (nx668), .A1 (nx100)) ;
    nor02ii ix134 (.Y (nx133), .A0 (nx100), .A1 (nx634)) ;
    and02 ix142 (.Y (nx141), .A0 (nx634), .A1 (nx94)) ;
    nor02ii ix146 (.Y (nx145), .A0 (nx94), .A1 (nx634)) ;
    and02 ix154 (.Y (nx153), .A0 (nx634), .A1 (nx88)) ;
    nor02ii ix158 (.Y (nx157), .A0 (nx88), .A1 (nx634)) ;
    inv01 ix647 (.Y (nx648), .A (nx630)) ;
    inv01 ix649 (.Y (nx650), .A (nx630)) ;
    inv01 ix651 (.Y (nx652), .A (nx630)) ;
    buf02 ix653 (.Y (nx654), .A (reset)) ;
    buf02 ix655 (.Y (nx656), .A (reset)) ;
    buf02 ix657 (.Y (nx658), .A (enable)) ;
    buf02 ix659 (.Y (nx660), .A (enable)) ;
    inv02 ix661 (.Y (nx662), .A (clk)) ;
    inv01 ix663 (.Y (nx664), .A (nx533)) ;
    inv01 ix665 (.Y (nx666), .A (nx533)) ;
    inv01 ix667 (.Y (nx668), .A (nx533)) ;
endmodule


module Counter_5 ( enable, reset, clk, load, \output , \input  ) ;

    input enable ;
    input reset ;
    input clk ;
    input load ;
    output [4:0]\output  ;
    input [4:0]\input  ;

    wire addResult_4, addResult_3, addResult_2, addResult_1, addResult_0, one_0, 
         one_4, nx64, NOT_clk, nx8, nx12, nx58, nx20, nx24, nx52, nx32, nx36, 
         nx46, nx44, nx49, nx40, nx57, nx61, nx172, nx182, nx192, nx202, nx212, 
         nx221, nx262, nx268, nx270;
    wire [10:0] \$dummy ;




    my_nadder_5 A1 (.a ({\output [4],\output [3],\output [2],\output [1],
                \output [0]}), .b ({one_4,one_4,one_4,one_4,one_0}), .cin (one_4
                ), .s ({addResult_4,addResult_3,addResult_2,addResult_1,
                addResult_0}), .cout (\$dummy [0])) ;
    fake_gnd ix146 (.Y (one_4)) ;
    fake_vcc ix144 (.Y (one_0)) ;
    dffsr_ni reg_toOutput_0__dup_1 (.Q (\output [0]), .QB (\$dummy [1]), .D (
             nx172), .CLK (clk), .S (nx8), .R (nx12)) ;
    mux21_ni ix173 (.Y (nx172), .A0 (\output [0]), .A1 (addResult_0), .S0 (nx268
             )) ;
    nor02ii ix9 (.Y (nx8), .A0 (nx262), .A1 (nx64)) ;
    nor02_2x ix222 (.Y (nx221), .A0 (nx270), .A1 (load)) ;
    dffr ix65 (.Q (nx64), .QB (\$dummy [2]), .D (\input [0]), .CLK (NOT_clk), .R (
         nx270)) ;
    inv01 ix225 (.Y (NOT_clk), .A (clk)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (nx64), .A1 (nx262)) ;
    dffsr_ni reg_toOutput_1__dup_1 (.Q (\output [1]), .QB (\$dummy [3]), .D (
             nx182), .CLK (clk), .S (nx20), .R (nx24)) ;
    mux21_ni ix183 (.Y (nx182), .A0 (\output [1]), .A1 (addResult_1), .S0 (nx268
             )) ;
    nor02ii ix21 (.Y (nx20), .A0 (nx262), .A1 (nx58)) ;
    dffr ix59 (.Q (nx58), .QB (\$dummy [4]), .D (\input [1]), .CLK (NOT_clk), .R (
         nx270)) ;
    nor02_2x ix25 (.Y (nx24), .A0 (nx58), .A1 (nx262)) ;
    dffsr_ni reg_toOutput_2__dup_1 (.Q (\output [2]), .QB (\$dummy [5]), .D (
             nx192), .CLK (clk), .S (nx32), .R (nx36)) ;
    mux21_ni ix193 (.Y (nx192), .A0 (\output [2]), .A1 (addResult_2), .S0 (nx268
             )) ;
    nor02ii ix33 (.Y (nx32), .A0 (nx262), .A1 (nx52)) ;
    dffr ix53 (.Q (nx52), .QB (\$dummy [6]), .D (\input [2]), .CLK (NOT_clk), .R (
         nx270)) ;
    nor02_2x ix37 (.Y (nx36), .A0 (nx52), .A1 (nx262)) ;
    dffsr_ni reg_toOutput_3__dup_1 (.Q (\output [3]), .QB (\$dummy [7]), .D (
             nx202), .CLK (clk), .S (nx44), .R (nx49)) ;
    mux21_ni ix203 (.Y (nx202), .A0 (\output [3]), .A1 (addResult_3), .S0 (nx268
             )) ;
    nor02ii ix45 (.Y (nx44), .A0 (nx262), .A1 (nx46)) ;
    dffr ix47 (.Q (nx46), .QB (\$dummy [8]), .D (\input [3]), .CLK (NOT_clk), .R (
         nx270)) ;
    nor02_2x ix50 (.Y (nx49), .A0 (nx46), .A1 (nx221)) ;
    dffsr_ni reg_toOutput_4__dup_1 (.Q (\output [4]), .QB (\$dummy [9]), .D (
             nx212), .CLK (clk), .S (nx57), .R (nx61)) ;
    mux21_ni ix213 (.Y (nx212), .A0 (\output [4]), .A1 (addResult_4), .S0 (nx268
             )) ;
    nor02ii ix58 (.Y (nx57), .A0 (nx221), .A1 (nx40)) ;
    dffr ix54 (.Q (nx40), .QB (\$dummy [10]), .D (\input [4]), .CLK (NOT_clk), .R (
         nx270)) ;
    nor02_2x ix62 (.Y (nx61), .A0 (nx40), .A1 (nx221)) ;
    nor02_2x ix261 (.Y (nx262), .A0 (nx270), .A1 (load)) ;
    buf02 ix267 (.Y (nx268), .A (enable)) ;
    buf02 ix269 (.Y (nx270), .A (reset)) ;
endmodule


module Convolution ( current_state, CLK, RST, QImgStat, ACK, LayerInfo, 
                     ImgAddress, OutputImg0, OutputImg1, OutputImg2, OutputImg3, 
                     OutputImg4, outFilter0, outFilter1, ConvOuput ) ;

    input [14:0]current_state ;
    input CLK ;
    input RST ;
    input QImgStat ;
    output ACK ;
    input [15:0]LayerInfo ;
    input [12:0]ImgAddress ;
    input [79:0]OutputImg0 ;
    input [79:0]OutputImg1 ;
    input [79:0]OutputImg2 ;
    input [79:0]OutputImg3 ;
    input [79:0]OutputImg4 ;
    input [399:0]outFilter0 ;
    input [399:0]outFilter1 ;
    output [15:0]ConvOuput ;

    wire FilterToAlu_399, FilterToAlu_398, FilterToAlu_397, FilterToAlu_396, 
         FilterToAlu_395, FilterToAlu_394, FilterToAlu_393, FilterToAlu_392, 
         FilterToAlu_391, FilterToAlu_390, FilterToAlu_389, FilterToAlu_388, 
         FilterToAlu_387, FilterToAlu_386, FilterToAlu_385, FilterToAlu_384, 
         FilterToAlu_383, FilterToAlu_382, FilterToAlu_381, FilterToAlu_380, 
         FilterToAlu_379, FilterToAlu_378, FilterToAlu_377, FilterToAlu_376, 
         FilterToAlu_375, FilterToAlu_374, FilterToAlu_373, FilterToAlu_372, 
         FilterToAlu_371, FilterToAlu_370, FilterToAlu_369, FilterToAlu_368, 
         FilterToAlu_367, FilterToAlu_366, FilterToAlu_365, FilterToAlu_364, 
         FilterToAlu_363, FilterToAlu_362, FilterToAlu_361, FilterToAlu_360, 
         FilterToAlu_359, FilterToAlu_358, FilterToAlu_357, FilterToAlu_356, 
         FilterToAlu_355, FilterToAlu_354, FilterToAlu_353, FilterToAlu_352, 
         FilterToAlu_351, FilterToAlu_350, FilterToAlu_349, FilterToAlu_348, 
         FilterToAlu_347, FilterToAlu_346, FilterToAlu_345, FilterToAlu_344, 
         FilterToAlu_343, FilterToAlu_342, FilterToAlu_341, FilterToAlu_340, 
         FilterToAlu_339, FilterToAlu_338, FilterToAlu_337, FilterToAlu_336, 
         FilterToAlu_335, FilterToAlu_334, FilterToAlu_333, FilterToAlu_332, 
         FilterToAlu_331, FilterToAlu_330, FilterToAlu_329, FilterToAlu_328, 
         FilterToAlu_327, FilterToAlu_326, FilterToAlu_325, FilterToAlu_324, 
         FilterToAlu_323, FilterToAlu_322, FilterToAlu_321, FilterToAlu_320, 
         FilterToAlu_319, FilterToAlu_318, FilterToAlu_317, FilterToAlu_316, 
         FilterToAlu_315, FilterToAlu_314, FilterToAlu_313, FilterToAlu_312, 
         FilterToAlu_311, FilterToAlu_310, FilterToAlu_309, FilterToAlu_308, 
         FilterToAlu_307, FilterToAlu_306, FilterToAlu_305, FilterToAlu_304, 
         FilterToAlu_303, FilterToAlu_302, FilterToAlu_301, FilterToAlu_300, 
         FilterToAlu_299, FilterToAlu_298, FilterToAlu_297, FilterToAlu_296, 
         FilterToAlu_295, FilterToAlu_294, FilterToAlu_293, FilterToAlu_292, 
         FilterToAlu_291, FilterToAlu_290, FilterToAlu_289, FilterToAlu_288, 
         FilterToAlu_287, FilterToAlu_286, FilterToAlu_285, FilterToAlu_284, 
         FilterToAlu_283, FilterToAlu_282, FilterToAlu_281, FilterToAlu_280, 
         FilterToAlu_279, FilterToAlu_278, FilterToAlu_277, FilterToAlu_276, 
         FilterToAlu_275, FilterToAlu_274, FilterToAlu_273, FilterToAlu_272, 
         FilterToAlu_271, FilterToAlu_270, FilterToAlu_269, FilterToAlu_268, 
         FilterToAlu_267, FilterToAlu_266, FilterToAlu_265, FilterToAlu_264, 
         FilterToAlu_263, FilterToAlu_262, FilterToAlu_261, FilterToAlu_260, 
         FilterToAlu_259, FilterToAlu_258, FilterToAlu_257, FilterToAlu_256, 
         FilterToAlu_255, FilterToAlu_254, FilterToAlu_253, FilterToAlu_252, 
         FilterToAlu_251, FilterToAlu_250, FilterToAlu_249, FilterToAlu_248, 
         FilterToAlu_247, FilterToAlu_246, FilterToAlu_245, FilterToAlu_244, 
         FilterToAlu_243, FilterToAlu_242, FilterToAlu_241, FilterToAlu_240, 
         FilterToAlu_239, FilterToAlu_238, FilterToAlu_237, FilterToAlu_236, 
         FilterToAlu_235, FilterToAlu_234, FilterToAlu_233, FilterToAlu_232, 
         FilterToAlu_231, FilterToAlu_230, FilterToAlu_229, FilterToAlu_228, 
         FilterToAlu_227, FilterToAlu_226, FilterToAlu_225, FilterToAlu_224, 
         FilterToAlu_223, FilterToAlu_222, FilterToAlu_221, FilterToAlu_220, 
         FilterToAlu_219, FilterToAlu_218, FilterToAlu_217, FilterToAlu_216, 
         FilterToAlu_215, FilterToAlu_214, FilterToAlu_213, FilterToAlu_212, 
         FilterToAlu_211, FilterToAlu_210, FilterToAlu_209, FilterToAlu_208, 
         FilterToAlu_207, FilterToAlu_206, FilterToAlu_205, FilterToAlu_204, 
         FilterToAlu_203, FilterToAlu_202, FilterToAlu_201, FilterToAlu_200, 
         FilterToAlu_199, FilterToAlu_198, FilterToAlu_197, FilterToAlu_196, 
         FilterToAlu_195, FilterToAlu_194, FilterToAlu_193, FilterToAlu_192, 
         FilterToAlu_191, FilterToAlu_190, FilterToAlu_189, FilterToAlu_188, 
         FilterToAlu_187, FilterToAlu_186, FilterToAlu_185, FilterToAlu_184, 
         FilterToAlu_183, FilterToAlu_182, FilterToAlu_181, FilterToAlu_180, 
         FilterToAlu_179, FilterToAlu_178, FilterToAlu_177, FilterToAlu_176, 
         FilterToAlu_175, FilterToAlu_174, FilterToAlu_173, FilterToAlu_172, 
         FilterToAlu_171, FilterToAlu_170, FilterToAlu_169, FilterToAlu_168, 
         FilterToAlu_167, FilterToAlu_166, FilterToAlu_165, FilterToAlu_164, 
         FilterToAlu_163, FilterToAlu_162, FilterToAlu_161, FilterToAlu_160, 
         FilterToAlu_159, FilterToAlu_158, FilterToAlu_157, FilterToAlu_156, 
         FilterToAlu_155, FilterToAlu_154, FilterToAlu_153, FilterToAlu_152, 
         FilterToAlu_151, FilterToAlu_150, FilterToAlu_149, FilterToAlu_148, 
         FilterToAlu_147, FilterToAlu_146, FilterToAlu_145, FilterToAlu_144, 
         FilterToAlu_143, FilterToAlu_142, FilterToAlu_141, FilterToAlu_140, 
         FilterToAlu_139, FilterToAlu_138, FilterToAlu_137, FilterToAlu_136, 
         FilterToAlu_135, FilterToAlu_134, FilterToAlu_133, FilterToAlu_132, 
         FilterToAlu_131, FilterToAlu_130, FilterToAlu_129, FilterToAlu_128, 
         FilterToAlu_127, FilterToAlu_126, FilterToAlu_125, FilterToAlu_124, 
         FilterToAlu_123, FilterToAlu_122, FilterToAlu_121, FilterToAlu_120, 
         FilterToAlu_119, FilterToAlu_118, FilterToAlu_117, FilterToAlu_116, 
         FilterToAlu_115, FilterToAlu_114, FilterToAlu_113, FilterToAlu_112, 
         FilterToAlu_111, FilterToAlu_110, FilterToAlu_109, FilterToAlu_108, 
         FilterToAlu_107, FilterToAlu_106, FilterToAlu_105, FilterToAlu_104, 
         FilterToAlu_103, FilterToAlu_102, FilterToAlu_101, FilterToAlu_100, 
         FilterToAlu_99, FilterToAlu_98, FilterToAlu_97, FilterToAlu_96, 
         FilterToAlu_95, FilterToAlu_94, FilterToAlu_93, FilterToAlu_92, 
         FilterToAlu_91, FilterToAlu_90, FilterToAlu_89, FilterToAlu_88, 
         FilterToAlu_87, FilterToAlu_86, FilterToAlu_85, FilterToAlu_84, 
         FilterToAlu_83, FilterToAlu_82, FilterToAlu_81, FilterToAlu_80, 
         FilterToAlu_79, FilterToAlu_78, FilterToAlu_77, FilterToAlu_76, 
         FilterToAlu_75, FilterToAlu_74, FilterToAlu_73, FilterToAlu_72, 
         FilterToAlu_71, FilterToAlu_70, FilterToAlu_69, FilterToAlu_68, 
         FilterToAlu_67, FilterToAlu_66, FilterToAlu_65, FilterToAlu_64, 
         FilterToAlu_63, FilterToAlu_62, FilterToAlu_61, FilterToAlu_60, 
         FilterToAlu_59, FilterToAlu_58, FilterToAlu_57, FilterToAlu_56, 
         FilterToAlu_55, FilterToAlu_54, FilterToAlu_53, FilterToAlu_52, 
         FilterToAlu_51, FilterToAlu_50, FilterToAlu_49, FilterToAlu_48, 
         FilterToAlu_47, FilterToAlu_46, FilterToAlu_45, FilterToAlu_44, 
         FilterToAlu_43, FilterToAlu_42, FilterToAlu_41, FilterToAlu_40, 
         FilterToAlu_39, FilterToAlu_38, FilterToAlu_37, FilterToAlu_36, 
         FilterToAlu_35, FilterToAlu_34, FilterToAlu_33, FilterToAlu_32, 
         FilterToAlu_31, FilterToAlu_30, FilterToAlu_29, FilterToAlu_28, 
         FilterToAlu_27, FilterToAlu_26, FilterToAlu_25, FilterToAlu_24, 
         FilterToAlu_23, FilterToAlu_22, FilterToAlu_21, FilterToAlu_20, 
         FilterToAlu_19, FilterToAlu_18, FilterToAlu_17, FilterToAlu_16, 
         FilterToAlu_15, FilterToAlu_14, FilterToAlu_13, FilterToAlu_12, 
         FilterToAlu_11, FilterToAlu_10, FilterToAlu_9, FilterToAlu_8, 
         FilterToAlu_7, FilterToAlu_6, FilterToAlu_5, FilterToAlu_4, 
         FilterToAlu_3, FilterToAlu_2, FilterToAlu_1, FilterToAlu_0, 
         MultiplierOut_792, MultiplierOut_791, MultiplierOut_790, 
         MultiplierOut_789, MultiplierOut_788, MultiplierOut_787, 
         MultiplierOut_786, MultiplierOut_785, MultiplierOut_784, 
         MultiplierOut_783, MultiplierOut_782, MultiplierOut_781, 
         MultiplierOut_780, MultiplierOut_779, MultiplierOut_778, 
         MultiplierOut_777, MultiplierOut_760, MultiplierOut_759, 
         MultiplierOut_758, MultiplierOut_757, MultiplierOut_756, 
         MultiplierOut_755, MultiplierOut_754, MultiplierOut_753, 
         MultiplierOut_752, MultiplierOut_751, MultiplierOut_750, 
         MultiplierOut_749, MultiplierOut_748, MultiplierOut_747, 
         MultiplierOut_746, MultiplierOut_745, MultiplierOut_728, 
         MultiplierOut_727, MultiplierOut_726, MultiplierOut_725, 
         MultiplierOut_724, MultiplierOut_723, MultiplierOut_722, 
         MultiplierOut_721, MultiplierOut_720, MultiplierOut_719, 
         MultiplierOut_718, MultiplierOut_717, MultiplierOut_716, 
         MultiplierOut_715, MultiplierOut_714, MultiplierOut_713, 
         MultiplierOut_696, MultiplierOut_695, MultiplierOut_694, 
         MultiplierOut_693, MultiplierOut_692, MultiplierOut_691, 
         MultiplierOut_690, MultiplierOut_689, MultiplierOut_688, 
         MultiplierOut_687, MultiplierOut_686, MultiplierOut_685, 
         MultiplierOut_684, MultiplierOut_683, MultiplierOut_682, 
         MultiplierOut_681, MultiplierOut_664, MultiplierOut_663, 
         MultiplierOut_662, MultiplierOut_661, MultiplierOut_660, 
         MultiplierOut_659, MultiplierOut_658, MultiplierOut_657, 
         MultiplierOut_656, MultiplierOut_655, MultiplierOut_654, 
         MultiplierOut_653, MultiplierOut_652, MultiplierOut_651, 
         MultiplierOut_650, MultiplierOut_649, MultiplierOut_632, 
         MultiplierOut_631, MultiplierOut_630, MultiplierOut_629, 
         MultiplierOut_628, MultiplierOut_627, MultiplierOut_626, 
         MultiplierOut_625, MultiplierOut_624, MultiplierOut_623, 
         MultiplierOut_622, MultiplierOut_621, MultiplierOut_620, 
         MultiplierOut_619, MultiplierOut_618, MultiplierOut_617, 
         MultiplierOut_600, MultiplierOut_599, MultiplierOut_598, 
         MultiplierOut_597, MultiplierOut_596, MultiplierOut_595, 
         MultiplierOut_594, MultiplierOut_593, MultiplierOut_592, 
         MultiplierOut_591, MultiplierOut_590, MultiplierOut_589, 
         MultiplierOut_588, MultiplierOut_587, MultiplierOut_586, 
         MultiplierOut_585, MultiplierOut_568, MultiplierOut_567, 
         MultiplierOut_566, MultiplierOut_565, MultiplierOut_564, 
         MultiplierOut_563, MultiplierOut_562, MultiplierOut_561, 
         MultiplierOut_560, MultiplierOut_559, MultiplierOut_558, 
         MultiplierOut_557, MultiplierOut_556, MultiplierOut_555, 
         MultiplierOut_554, MultiplierOut_553, MultiplierOut_536, 
         MultiplierOut_535, MultiplierOut_534, MultiplierOut_533, 
         MultiplierOut_532, MultiplierOut_531, MultiplierOut_530, 
         MultiplierOut_529, MultiplierOut_528, MultiplierOut_527, 
         MultiplierOut_526, MultiplierOut_525, MultiplierOut_524, 
         MultiplierOut_523, MultiplierOut_522, MultiplierOut_521, 
         MultiplierOut_504, MultiplierOut_503, MultiplierOut_502, 
         MultiplierOut_501, MultiplierOut_500, MultiplierOut_499, 
         MultiplierOut_498, MultiplierOut_497, MultiplierOut_496, 
         MultiplierOut_495, MultiplierOut_494, MultiplierOut_493, 
         MultiplierOut_492, MultiplierOut_491, MultiplierOut_490, 
         MultiplierOut_489, MultiplierOut_472, MultiplierOut_471, 
         MultiplierOut_470, MultiplierOut_469, MultiplierOut_468, 
         MultiplierOut_467, MultiplierOut_466, MultiplierOut_465, 
         MultiplierOut_464, MultiplierOut_463, MultiplierOut_462, 
         MultiplierOut_461, MultiplierOut_460, MultiplierOut_459, 
         MultiplierOut_458, MultiplierOut_457, MultiplierOut_440, 
         MultiplierOut_439, MultiplierOut_438, MultiplierOut_437, 
         MultiplierOut_436, MultiplierOut_435, MultiplierOut_434, 
         MultiplierOut_433, MultiplierOut_432, MultiplierOut_431, 
         MultiplierOut_430, MultiplierOut_429, MultiplierOut_428, 
         MultiplierOut_427, MultiplierOut_426, MultiplierOut_425, 
         MultiplierOut_408, MultiplierOut_407, MultiplierOut_406, 
         MultiplierOut_405, MultiplierOut_404, MultiplierOut_403, 
         MultiplierOut_402, MultiplierOut_401, MultiplierOut_400, 
         MultiplierOut_399, MultiplierOut_398, MultiplierOut_397, 
         MultiplierOut_396, MultiplierOut_395, MultiplierOut_394, 
         MultiplierOut_393, MultiplierOut_376, MultiplierOut_375, 
         MultiplierOut_374, MultiplierOut_373, MultiplierOut_372, 
         MultiplierOut_371, MultiplierOut_370, MultiplierOut_369, 
         MultiplierOut_368, MultiplierOut_367, MultiplierOut_366, 
         MultiplierOut_365, MultiplierOut_364, MultiplierOut_363, 
         MultiplierOut_362, MultiplierOut_361, MultiplierOut_344, 
         MultiplierOut_343, MultiplierOut_342, MultiplierOut_341, 
         MultiplierOut_340, MultiplierOut_339, MultiplierOut_338, 
         MultiplierOut_337, MultiplierOut_336, MultiplierOut_335, 
         MultiplierOut_334, MultiplierOut_333, MultiplierOut_332, 
         MultiplierOut_331, MultiplierOut_330, MultiplierOut_329, 
         MultiplierOut_312, MultiplierOut_311, MultiplierOut_310, 
         MultiplierOut_309, MultiplierOut_308, MultiplierOut_307, 
         MultiplierOut_306, MultiplierOut_305, MultiplierOut_304, 
         MultiplierOut_303, MultiplierOut_302, MultiplierOut_301, 
         MultiplierOut_300, MultiplierOut_299, MultiplierOut_298, 
         MultiplierOut_297, MultiplierOut_280, MultiplierOut_279, 
         MultiplierOut_278, MultiplierOut_277, MultiplierOut_276, 
         MultiplierOut_275, MultiplierOut_274, MultiplierOut_273, 
         MultiplierOut_272, MultiplierOut_271, MultiplierOut_270, 
         MultiplierOut_269, MultiplierOut_268, MultiplierOut_267, 
         MultiplierOut_266, MultiplierOut_265, MultiplierOut_248, 
         MultiplierOut_247, MultiplierOut_246, MultiplierOut_245, 
         MultiplierOut_244, MultiplierOut_243, MultiplierOut_242, 
         MultiplierOut_241, MultiplierOut_240, MultiplierOut_239, 
         MultiplierOut_238, MultiplierOut_237, MultiplierOut_236, 
         MultiplierOut_235, MultiplierOut_234, MultiplierOut_233, 
         MultiplierOut_216, MultiplierOut_215, MultiplierOut_214, 
         MultiplierOut_213, MultiplierOut_212, MultiplierOut_211, 
         MultiplierOut_210, MultiplierOut_209, MultiplierOut_208, 
         MultiplierOut_207, MultiplierOut_206, MultiplierOut_205, 
         MultiplierOut_204, MultiplierOut_203, MultiplierOut_202, 
         MultiplierOut_201, MultiplierOut_184, MultiplierOut_183, 
         MultiplierOut_182, MultiplierOut_181, MultiplierOut_180, 
         MultiplierOut_179, MultiplierOut_178, MultiplierOut_177, 
         MultiplierOut_176, MultiplierOut_175, MultiplierOut_174, 
         MultiplierOut_173, MultiplierOut_172, MultiplierOut_171, 
         MultiplierOut_170, MultiplierOut_169, MultiplierOut_152, 
         MultiplierOut_151, MultiplierOut_150, MultiplierOut_149, 
         MultiplierOut_148, MultiplierOut_147, MultiplierOut_146, 
         MultiplierOut_145, MultiplierOut_144, MultiplierOut_143, 
         MultiplierOut_142, MultiplierOut_141, MultiplierOut_140, 
         MultiplierOut_139, MultiplierOut_138, MultiplierOut_137, 
         MultiplierOut_120, MultiplierOut_119, MultiplierOut_118, 
         MultiplierOut_117, MultiplierOut_116, MultiplierOut_115, 
         MultiplierOut_114, MultiplierOut_113, MultiplierOut_112, 
         MultiplierOut_111, MultiplierOut_110, MultiplierOut_109, 
         MultiplierOut_108, MultiplierOut_107, MultiplierOut_106, 
         MultiplierOut_105, MultiplierOut_88, MultiplierOut_87, MultiplierOut_86, 
         MultiplierOut_85, MultiplierOut_84, MultiplierOut_83, MultiplierOut_82, 
         MultiplierOut_81, MultiplierOut_80, MultiplierOut_79, MultiplierOut_78, 
         MultiplierOut_77, MultiplierOut_76, MultiplierOut_75, MultiplierOut_74, 
         MultiplierOut_73, MultiplierOut_56, MultiplierOut_55, MultiplierOut_54, 
         MultiplierOut_53, MultiplierOut_52, MultiplierOut_51, MultiplierOut_50, 
         MultiplierOut_49, MultiplierOut_48, MultiplierOut_47, MultiplierOut_46, 
         MultiplierOut_45, MultiplierOut_44, MultiplierOut_43, MultiplierOut_42, 
         MultiplierOut_41, MultiplierOut_24, MultiplierOut_23, MultiplierOut_22, 
         MultiplierOut_21, MultiplierOut_20, MultiplierOut_19, MultiplierOut_18, 
         MultiplierOut_17, MultiplierOut_16, MultiplierOut_15, MultiplierOut_14, 
         MultiplierOut_13, MultiplierOut_12, MultiplierOut_11, MultiplierOut_10, 
         MultiplierOut_9, AddOutputLvL1_191, AddOutputLvL1_190, 
         AddOutputLvL1_189, AddOutputLvL1_188, AddOutputLvL1_187, 
         AddOutputLvL1_186, AddOutputLvL1_185, AddOutputLvL1_184, 
         AddOutputLvL1_183, AddOutputLvL1_182, AddOutputLvL1_181, 
         AddOutputLvL1_180, AddOutputLvL1_179, AddOutputLvL1_178, 
         AddOutputLvL1_177, AddOutputLvL1_176, AddOutputLvL1_175, 
         AddOutputLvL1_174, AddOutputLvL1_173, AddOutputLvL1_172, 
         AddOutputLvL1_171, AddOutputLvL1_170, AddOutputLvL1_169, 
         AddOutputLvL1_168, AddOutputLvL1_167, AddOutputLvL1_166, 
         AddOutputLvL1_165, AddOutputLvL1_164, AddOutputLvL1_163, 
         AddOutputLvL1_162, AddOutputLvL1_161, AddOutputLvL1_160, 
         AddOutputLvL1_159, AddOutputLvL1_158, AddOutputLvL1_157, 
         AddOutputLvL1_156, AddOutputLvL1_155, AddOutputLvL1_154, 
         AddOutputLvL1_153, AddOutputLvL1_152, AddOutputLvL1_151, 
         AddOutputLvL1_150, AddOutputLvL1_149, AddOutputLvL1_148, 
         AddOutputLvL1_147, AddOutputLvL1_146, AddOutputLvL1_145, 
         AddOutputLvL1_144, AddOutputLvL1_143, AddOutputLvL1_142, 
         AddOutputLvL1_141, AddOutputLvL1_140, AddOutputLvL1_139, 
         AddOutputLvL1_138, AddOutputLvL1_137, AddOutputLvL1_136, 
         AddOutputLvL1_135, AddOutputLvL1_134, AddOutputLvL1_133, 
         AddOutputLvL1_132, AddOutputLvL1_131, AddOutputLvL1_130, 
         AddOutputLvL1_129, AddOutputLvL1_128, AddOutputLvL1_127, 
         AddOutputLvL1_126, AddOutputLvL1_125, AddOutputLvL1_124, 
         AddOutputLvL1_123, AddOutputLvL1_122, AddOutputLvL1_121, 
         AddOutputLvL1_120, AddOutputLvL1_119, AddOutputLvL1_118, 
         AddOutputLvL1_117, AddOutputLvL1_116, AddOutputLvL1_115, 
         AddOutputLvL1_114, AddOutputLvL1_113, AddOutputLvL1_112, 
         AddOutputLvL1_111, AddOutputLvL1_110, AddOutputLvL1_109, 
         AddOutputLvL1_108, AddOutputLvL1_107, AddOutputLvL1_106, 
         AddOutputLvL1_105, AddOutputLvL1_104, AddOutputLvL1_103, 
         AddOutputLvL1_102, AddOutputLvL1_101, AddOutputLvL1_100, 
         AddOutputLvL1_99, AddOutputLvL1_98, AddOutputLvL1_97, AddOutputLvL1_96, 
         AddOutputLvL1_95, AddOutputLvL1_94, AddOutputLvL1_93, AddOutputLvL1_92, 
         AddOutputLvL1_91, AddOutputLvL1_90, AddOutputLvL1_89, AddOutputLvL1_88, 
         AddOutputLvL1_87, AddOutputLvL1_86, AddOutputLvL1_85, AddOutputLvL1_84, 
         AddOutputLvL1_83, AddOutputLvL1_82, AddOutputLvL1_81, AddOutputLvL1_80, 
         AddOutputLvL1_79, AddOutputLvL1_78, AddOutputLvL1_77, AddOutputLvL1_76, 
         AddOutputLvL1_75, AddOutputLvL1_74, AddOutputLvL1_73, AddOutputLvL1_72, 
         AddOutputLvL1_71, AddOutputLvL1_70, AddOutputLvL1_69, AddOutputLvL1_68, 
         AddOutputLvL1_67, AddOutputLvL1_66, AddOutputLvL1_65, AddOutputLvL1_64, 
         AddOutputLvL1_63, AddOutputLvL1_62, AddOutputLvL1_61, AddOutputLvL1_60, 
         AddOutputLvL1_59, AddOutputLvL1_58, AddOutputLvL1_57, AddOutputLvL1_56, 
         AddOutputLvL1_55, AddOutputLvL1_54, AddOutputLvL1_53, AddOutputLvL1_52, 
         AddOutputLvL1_51, AddOutputLvL1_50, AddOutputLvL1_49, AddOutputLvL1_48, 
         AddOutputLvL1_47, AddOutputLvL1_46, AddOutputLvL1_45, AddOutputLvL1_44, 
         AddOutputLvL1_43, AddOutputLvL1_42, AddOutputLvL1_41, AddOutputLvL1_40, 
         AddOutputLvL1_39, AddOutputLvL1_38, AddOutputLvL1_37, AddOutputLvL1_36, 
         AddOutputLvL1_35, AddOutputLvL1_34, AddOutputLvL1_33, AddOutputLvL1_32, 
         AddOutputLvL1_31, AddOutputLvL1_30, AddOutputLvL1_29, AddOutputLvL1_28, 
         AddOutputLvL1_27, AddOutputLvL1_26, AddOutputLvL1_25, AddOutputLvL1_24, 
         AddOutputLvL1_23, AddOutputLvL1_22, AddOutputLvL1_21, AddOutputLvL1_20, 
         AddOutputLvL1_19, AddOutputLvL1_18, AddOutputLvL1_17, AddOutputLvL1_16, 
         AddOutputLvL1_15, AddOutputLvL1_14, AddOutputLvL1_13, AddOutputLvL1_12, 
         AddOutputLvL1_11, AddOutputLvL1_10, AddOutputLvL1_9, AddOutputLvL1_8, 
         AddOutputLvL1_7, AddOutputLvL1_6, AddOutputLvL1_5, AddOutputLvL1_4, 
         AddOutputLvL1_3, AddOutputLvL1_2, AddOutputLvL1_1, AddOutputLvL1_0, 
         AddOutputLvL2_95, AddOutputLvL2_94, AddOutputLvL2_93, AddOutputLvL2_92, 
         AddOutputLvL2_91, AddOutputLvL2_90, AddOutputLvL2_89, AddOutputLvL2_88, 
         AddOutputLvL2_87, AddOutputLvL2_86, AddOutputLvL2_85, AddOutputLvL2_84, 
         AddOutputLvL2_83, AddOutputLvL2_82, AddOutputLvL2_81, AddOutputLvL2_80, 
         AddOutputLvL2_79, AddOutputLvL2_78, AddOutputLvL2_77, AddOutputLvL2_76, 
         AddOutputLvL2_75, AddOutputLvL2_74, AddOutputLvL2_73, AddOutputLvL2_72, 
         AddOutputLvL2_71, AddOutputLvL2_70, AddOutputLvL2_69, AddOutputLvL2_68, 
         AddOutputLvL2_67, AddOutputLvL2_66, AddOutputLvL2_65, AddOutputLvL2_64, 
         AddOutputLvL2_63, AddOutputLvL2_62, AddOutputLvL2_61, AddOutputLvL2_60, 
         AddOutputLvL2_59, AddOutputLvL2_58, AddOutputLvL2_57, AddOutputLvL2_56, 
         AddOutputLvL2_55, AddOutputLvL2_54, AddOutputLvL2_53, AddOutputLvL2_52, 
         AddOutputLvL2_51, AddOutputLvL2_50, AddOutputLvL2_49, AddOutputLvL2_48, 
         AddOutputLvL2_47, AddOutputLvL2_46, AddOutputLvL2_45, AddOutputLvL2_44, 
         AddOutputLvL2_43, AddOutputLvL2_42, AddOutputLvL2_41, AddOutputLvL2_40, 
         AddOutputLvL2_39, AddOutputLvL2_38, AddOutputLvL2_37, AddOutputLvL2_36, 
         AddOutputLvL2_35, AddOutputLvL2_34, AddOutputLvL2_33, AddOutputLvL2_32, 
         AddOutputLvL2_31, AddOutputLvL2_30, AddOutputLvL2_29, AddOutputLvL2_28, 
         AddOutputLvL2_27, AddOutputLvL2_26, AddOutputLvL2_25, AddOutputLvL2_24, 
         AddOutputLvL2_23, AddOutputLvL2_22, AddOutputLvL2_21, AddOutputLvL2_20, 
         AddOutputLvL2_19, AddOutputLvL2_18, AddOutputLvL2_17, AddOutputLvL2_16, 
         AddOutputLvL2_15, AddOutputLvL2_14, AddOutputLvL2_13, AddOutputLvL2_12, 
         AddOutputLvL2_11, AddOutputLvL2_10, AddOutputLvL2_9, AddOutputLvL2_8, 
         AddOutputLvL2_7, AddOutputLvL2_6, AddOutputLvL2_5, AddOutputLvL2_4, 
         AddOutputLvL2_3, AddOutputLvL2_2, AddOutputLvL2_1, AddOutputLvL2_0, 
         AddOutputLvL3_47, AddOutputLvL3_46, AddOutputLvL3_45, AddOutputLvL3_44, 
         AddOutputLvL3_43, AddOutputLvL3_42, AddOutputLvL3_41, AddOutputLvL3_40, 
         AddOutputLvL3_39, AddOutputLvL3_38, AddOutputLvL3_37, AddOutputLvL3_36, 
         AddOutputLvL3_35, AddOutputLvL3_34, AddOutputLvL3_33, AddOutputLvL3_32, 
         AddOutputLvL3_31, AddOutputLvL3_30, AddOutputLvL3_29, AddOutputLvL3_28, 
         AddOutputLvL3_27, AddOutputLvL3_26, AddOutputLvL3_25, AddOutputLvL3_24, 
         AddOutputLvL3_23, AddOutputLvL3_22, AddOutputLvL3_21, AddOutputLvL3_20, 
         AddOutputLvL3_19, AddOutputLvL3_18, AddOutputLvL3_17, AddOutputLvL3_16, 
         AddOutputLvL3_15, AddOutputLvL3_14, AddOutputLvL3_13, AddOutputLvL3_12, 
         AddOutputLvL3_11, AddOutputLvL3_10, AddOutputLvL3_9, AddOutputLvL3_8, 
         AddOutputLvL3_7, AddOutputLvL3_6, AddOutputLvL3_5, AddOutputLvL3_4, 
         AddOutputLvL3_3, AddOutputLvL3_2, AddOutputLvL3_1, AddOutputLvL3_0, 
         AddOut33_15, AddOut33_14, AddOut33_13, AddOut33_12, AddOut33_11, 
         AddOut33_10, AddOut33_9, AddOut33_8, AddOut33_7, AddOut33_6, AddOut33_5, 
         AddOut33_4, AddOut33_3, AddOut33_2, AddOut33_1, AddOut33_0, AddOut55_15, 
         AddOut55_14, AddOut55_13, AddOut55_12, AddOut55_11, AddOut55_10, 
         AddOut55_9, AddOut55_8, AddOut55_7, AddOut55_6, AddOut55_5, AddOut55_4, 
         AddOut55_3, AddOut55_2, AddOut55_1, AddOut55_0, Final55_15, Final55_14, 
         Final55_13, Final55_12, Final55_11, Final55_10, Final55_9, Final55_8, 
         Final55_7, Final55_6, Final55_5, Final55_4, Final55_3, Final55_2, 
         Final55_1, Final55_0, CounterOut_2, CounterOut_1, CounterOut_0, 
         SecondInputToMult_143, SecondInputToMult_142, SecondInputToMult_141, 
         SecondInputToMult_140, SecondInputToMult_139, SecondInputToMult_138, 
         SecondInputToMult_137, SecondInputToMult_136, SecondInputToMult_135, 
         SecondInputToMult_134, SecondInputToMult_133, SecondInputToMult_132, 
         SecondInputToMult_131, SecondInputToMult_130, SecondInputToMult_129, 
         SecondInputToMult_128, SecondInputToMult_127, SecondInputToMult_126, 
         SecondInputToMult_125, SecondInputToMult_124, SecondInputToMult_123, 
         SecondInputToMult_122, SecondInputToMult_121, SecondInputToMult_120, 
         SecondInputToMult_119, SecondInputToMult_118, SecondInputToMult_117, 
         SecondInputToMult_116, SecondInputToMult_115, SecondInputToMult_114, 
         SecondInputToMult_113, SecondInputToMult_112, SecondInputToMult_111, 
         SecondInputToMult_110, SecondInputToMult_109, SecondInputToMult_108, 
         SecondInputToMult_107, SecondInputToMult_106, SecondInputToMult_105, 
         SecondInputToMult_104, SecondInputToMult_103, SecondInputToMult_102, 
         SecondInputToMult_101, SecondInputToMult_100, SecondInputToMult_99, 
         SecondInputToMult_98, SecondInputToMult_97, SecondInputToMult_96, 
         SecondInputToMult_95, SecondInputToMult_94, SecondInputToMult_93, 
         SecondInputToMult_92, SecondInputToMult_91, SecondInputToMult_90, 
         SecondInputToMult_89, SecondInputToMult_88, SecondInputToMult_87, 
         SecondInputToMult_86, SecondInputToMult_85, SecondInputToMult_84, 
         SecondInputToMult_83, SecondInputToMult_82, SecondInputToMult_81, 
         SecondInputToMult_80, SecondInputToMult_79, SecondInputToMult_78, 
         SecondInputToMult_77, SecondInputToMult_76, SecondInputToMult_75, 
         SecondInputToMult_74, SecondInputToMult_73, SecondInputToMult_72, 
         SecondInputToMult_71, SecondInputToMult_70, SecondInputToMult_69, 
         SecondInputToMult_68, SecondInputToMult_67, SecondInputToMult_66, 
         SecondInputToMult_65, SecondInputToMult_64, SecondInputToMult_63, 
         SecondInputToMult_62, SecondInputToMult_61, SecondInputToMult_60, 
         SecondInputToMult_59, SecondInputToMult_58, SecondInputToMult_57, 
         SecondInputToMult_56, SecondInputToMult_55, SecondInputToMult_54, 
         SecondInputToMult_53, SecondInputToMult_52, SecondInputToMult_51, 
         SecondInputToMult_50, SecondInputToMult_49, SecondInputToMult_48, 
         CountereEN, CountereRST, GND0, nx6, nx12, nx20, nx32, nx34, nx48, nx68, 
         nx98, nx116, nx134, nx152, nx170, nx188, nx206, nx224, nx510, nx516, 
         nx3552, nx3562, nx7936, nx8052, nx8072, nx8090, nx8108, nx8126, nx8144, 
         nx8162, nx8180, nx8198, nx8216, nx8234, nx8252, nx8270, nx8288, nx8306, 
         nx8324, nx8342, nx8360, nx8378, nx8396, nx8414, nx8432, nx8450, nx8468, 
         nx8486, nx8495, nx8501, nx8511, nx8514, nx8517, nx8520, nx8523, nx8525, 
         nx8528, nx8530, nx8534, nx8536, nx8540, nx8542, nx8546, nx8548, nx8552, 
         nx8554, nx8558, nx8560, nx8564, nx8566, nx8569, nx8571, nx8586, nx8588, 
         nx8590, nx8592, nx8594, nx8596, nx8598, nx8600, nx8602, nx8604, nx8606, 
         nx8608, nx8610, nx8612, nx8614, nx8616, nx8618, nx8620, nx8622, nx8624, 
         nx8626, nx8628, nx8630, nx8632, nx8634, nx8636, nx8638, nx8640, nx8642, 
         nx8644, nx8646, nx8648, nx8650, nx8652, nx8654, nx8656, nx8658, nx8660, 
         nx8662, nx8664, nx8666, nx8668, nx8670, nx8672, nx8674, nx8676, nx8678, 
         nx8680, nx8682, nx8684, nx8686, nx8688, nx8690, nx8692, nx8696, nx8698, 
         nx8700, nx8702, nx8704, nx8706, nx8708, nx8710, nx8712, nx8714, nx8716, 
         nx8718, nx8720, nx8722, nx8724, nx8726, nx8728, nx8730, nx8732, nx8734, 
         nx8736, nx8738, nx8740, nx8742, nx8744, nx8746, nx8748, nx8750, nx8752, 
         nx8754, nx8756, nx8758, nx8760, nx8762, nx8764, nx8766, nx8768, nx8770, 
         nx8772, nx8774, nx8776, nx8778, nx8780, nx8782, nx8784, nx8786, nx8788, 
         nx8790, nx8792, nx8794, nx8796, nx8798, nx8800, nx8802, nx8804, nx8806, 
         nx8808, nx8810, nx8812, nx8814, nx8816, nx8818, nx8820, nx8822, nx8824, 
         nx8826, nx8828, nx8830, nx8832, nx8834, nx8836, nx8838, nx8840, nx8842, 
         nx8844, nx8846, nx8852, nx8854, nx8856, nx8858, nx8860, nx8862, nx8864, 
         nx8866, nx8868, nx8870, nx8872, nx8874, nx8876, nx8878, nx8880, nx8882, 
         nx8884, nx8886, nx8888, nx8890, nx8892, nx8894, nx8896, nx8898, nx8900, 
         nx8902, nx8904, nx8906, nx8908, nx8910, nx8912, nx8914, nx8916, nx8918, 
         nx8920, nx8922, nx8924, nx8926;
    wire [424:0] \$dummy ;




    Multiplier_16 loop3_0_Multip (.A ({FilterToAlu_15,FilterToAlu_14,
                  FilterToAlu_13,FilterToAlu_12,FilterToAlu_11,FilterToAlu_10,
                  FilterToAlu_9,FilterToAlu_8,FilterToAlu_7,FilterToAlu_6,
                  FilterToAlu_5,FilterToAlu_4,FilterToAlu_3,FilterToAlu_2,
                  FilterToAlu_1,FilterToAlu_0}), .B ({OutputImg0[15],
                  OutputImg0[14],OutputImg0[13],OutputImg0[12],OutputImg0[11],
                  OutputImg0[10],OutputImg0[9],OutputImg0[8],OutputImg0[7],
                  OutputImg0[6],OutputImg0[5],OutputImg0[4],OutputImg0[3],
                  OutputImg0[2],OutputImg0[1],OutputImg0[0]}), .F ({\$dummy [0],
                  \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                  \$dummy [6],MultiplierOut_24,MultiplierOut_23,MultiplierOut_22
                  ,MultiplierOut_21,MultiplierOut_20,MultiplierOut_19,
                  MultiplierOut_18,MultiplierOut_17,MultiplierOut_16,
                  MultiplierOut_15,MultiplierOut_14,MultiplierOut_13,
                  MultiplierOut_12,MultiplierOut_11,MultiplierOut_10,
                  MultiplierOut_9,\$dummy [7],\$dummy [8],\$dummy [9],
                  \$dummy [10],\$dummy [11],\$dummy [12],\$dummy [13],
                  \$dummy [14],\$dummy [15]})) ;
    Multiplier_16 loop3_1_Multip (.A ({FilterToAlu_31,FilterToAlu_30,
                  FilterToAlu_29,FilterToAlu_28,FilterToAlu_27,FilterToAlu_26,
                  FilterToAlu_25,FilterToAlu_24,FilterToAlu_23,FilterToAlu_22,
                  FilterToAlu_21,FilterToAlu_20,FilterToAlu_19,FilterToAlu_18,
                  FilterToAlu_17,FilterToAlu_16}), .B ({OutputImg0[31],
                  OutputImg0[30],OutputImg0[29],OutputImg0[28],OutputImg0[27],
                  OutputImg0[26],OutputImg0[25],OutputImg0[24],OutputImg0[23],
                  OutputImg0[22],OutputImg0[21],OutputImg0[20],OutputImg0[19],
                  OutputImg0[18],OutputImg0[17],OutputImg0[16]}), .F ({
                  \$dummy [16],\$dummy [17],\$dummy [18],\$dummy [19],
                  \$dummy [20],\$dummy [21],\$dummy [22],MultiplierOut_56,
                  MultiplierOut_55,MultiplierOut_54,MultiplierOut_53,
                  MultiplierOut_52,MultiplierOut_51,MultiplierOut_50,
                  MultiplierOut_49,MultiplierOut_48,MultiplierOut_47,
                  MultiplierOut_46,MultiplierOut_45,MultiplierOut_44,
                  MultiplierOut_43,MultiplierOut_42,MultiplierOut_41,
                  \$dummy [23],\$dummy [24],\$dummy [25],\$dummy [26],
                  \$dummy [27],\$dummy [28],\$dummy [29],\$dummy [30],
                  \$dummy [31]})) ;
    Multiplier_16 loop3_2_Multip (.A ({FilterToAlu_47,FilterToAlu_46,
                  FilterToAlu_45,FilterToAlu_44,FilterToAlu_43,FilterToAlu_42,
                  FilterToAlu_41,FilterToAlu_40,FilterToAlu_39,FilterToAlu_38,
                  FilterToAlu_37,FilterToAlu_36,FilterToAlu_35,FilterToAlu_34,
                  FilterToAlu_33,FilterToAlu_32}), .B ({OutputImg0[47],
                  OutputImg0[46],OutputImg0[45],OutputImg0[44],OutputImg0[43],
                  OutputImg0[42],OutputImg0[41],OutputImg0[40],OutputImg0[39],
                  OutputImg0[38],OutputImg0[37],OutputImg0[36],OutputImg0[35],
                  OutputImg0[34],OutputImg0[33],OutputImg0[32]}), .F ({
                  \$dummy [32],\$dummy [33],\$dummy [34],\$dummy [35],
                  \$dummy [36],\$dummy [37],\$dummy [38],MultiplierOut_88,
                  MultiplierOut_87,MultiplierOut_86,MultiplierOut_85,
                  MultiplierOut_84,MultiplierOut_83,MultiplierOut_82,
                  MultiplierOut_81,MultiplierOut_80,MultiplierOut_79,
                  MultiplierOut_78,MultiplierOut_77,MultiplierOut_76,
                  MultiplierOut_75,MultiplierOut_74,MultiplierOut_73,
                  \$dummy [39],\$dummy [40],\$dummy [41],\$dummy [42],
                  \$dummy [43],\$dummy [44],\$dummy [45],\$dummy [46],
                  \$dummy [47]})) ;
    Multiplier_16 loop3_3_Multip (.A ({FilterToAlu_63,FilterToAlu_62,
                  FilterToAlu_61,FilterToAlu_60,FilterToAlu_59,FilterToAlu_58,
                  FilterToAlu_57,FilterToAlu_56,FilterToAlu_55,FilterToAlu_54,
                  FilterToAlu_53,FilterToAlu_52,FilterToAlu_51,FilterToAlu_50,
                  FilterToAlu_49,FilterToAlu_48}), .B ({SecondInputToMult_63,
                  SecondInputToMult_62,SecondInputToMult_61,SecondInputToMult_60
                  ,SecondInputToMult_59,SecondInputToMult_58,
                  SecondInputToMult_57,SecondInputToMult_56,SecondInputToMult_55
                  ,SecondInputToMult_54,SecondInputToMult_53,
                  SecondInputToMult_52,SecondInputToMult_51,SecondInputToMult_50
                  ,SecondInputToMult_49,SecondInputToMult_48}), .F ({
                  \$dummy [48],\$dummy [49],\$dummy [50],\$dummy [51],
                  \$dummy [52],\$dummy [53],\$dummy [54],MultiplierOut_120,
                  MultiplierOut_119,MultiplierOut_118,MultiplierOut_117,
                  MultiplierOut_116,MultiplierOut_115,MultiplierOut_114,
                  MultiplierOut_113,MultiplierOut_112,MultiplierOut_111,
                  MultiplierOut_110,MultiplierOut_109,MultiplierOut_108,
                  MultiplierOut_107,MultiplierOut_106,MultiplierOut_105,
                  \$dummy [55],\$dummy [56],\$dummy [57],\$dummy [58],
                  \$dummy [59],\$dummy [60],\$dummy [61],\$dummy [62],
                  \$dummy [63]})) ;
    Multiplier_16 loop3_4_Multip (.A ({FilterToAlu_79,FilterToAlu_78,
                  FilterToAlu_77,FilterToAlu_76,FilterToAlu_75,FilterToAlu_74,
                  FilterToAlu_73,FilterToAlu_72,FilterToAlu_71,FilterToAlu_70,
                  FilterToAlu_69,FilterToAlu_68,FilterToAlu_67,FilterToAlu_66,
                  FilterToAlu_65,FilterToAlu_64}), .B ({SecondInputToMult_79,
                  SecondInputToMult_78,SecondInputToMult_77,SecondInputToMult_76
                  ,SecondInputToMult_75,SecondInputToMult_74,
                  SecondInputToMult_73,SecondInputToMult_72,SecondInputToMult_71
                  ,SecondInputToMult_70,SecondInputToMult_69,
                  SecondInputToMult_68,SecondInputToMult_67,SecondInputToMult_66
                  ,SecondInputToMult_65,SecondInputToMult_64}), .F ({
                  \$dummy [64],\$dummy [65],\$dummy [66],\$dummy [67],
                  \$dummy [68],\$dummy [69],\$dummy [70],MultiplierOut_152,
                  MultiplierOut_151,MultiplierOut_150,MultiplierOut_149,
                  MultiplierOut_148,MultiplierOut_147,MultiplierOut_146,
                  MultiplierOut_145,MultiplierOut_144,MultiplierOut_143,
                  MultiplierOut_142,MultiplierOut_141,MultiplierOut_140,
                  MultiplierOut_139,MultiplierOut_138,MultiplierOut_137,
                  \$dummy [71],\$dummy [72],\$dummy [73],\$dummy [74],
                  \$dummy [75],\$dummy [76],\$dummy [77],\$dummy [78],
                  \$dummy [79]})) ;
    Multiplier_16 loop3_5_Multip (.A ({FilterToAlu_95,FilterToAlu_94,
                  FilterToAlu_93,FilterToAlu_92,FilterToAlu_91,FilterToAlu_90,
                  FilterToAlu_89,FilterToAlu_88,FilterToAlu_87,FilterToAlu_86,
                  FilterToAlu_85,FilterToAlu_84,FilterToAlu_83,FilterToAlu_82,
                  FilterToAlu_81,FilterToAlu_80}), .B ({SecondInputToMult_95,
                  SecondInputToMult_94,SecondInputToMult_93,SecondInputToMult_92
                  ,SecondInputToMult_91,SecondInputToMult_90,
                  SecondInputToMult_89,SecondInputToMult_88,SecondInputToMult_87
                  ,SecondInputToMult_86,SecondInputToMult_85,
                  SecondInputToMult_84,SecondInputToMult_83,SecondInputToMult_82
                  ,SecondInputToMult_81,SecondInputToMult_80}), .F ({
                  \$dummy [80],\$dummy [81],\$dummy [82],\$dummy [83],
                  \$dummy [84],\$dummy [85],\$dummy [86],MultiplierOut_184,
                  MultiplierOut_183,MultiplierOut_182,MultiplierOut_181,
                  MultiplierOut_180,MultiplierOut_179,MultiplierOut_178,
                  MultiplierOut_177,MultiplierOut_176,MultiplierOut_175,
                  MultiplierOut_174,MultiplierOut_173,MultiplierOut_172,
                  MultiplierOut_171,MultiplierOut_170,MultiplierOut_169,
                  \$dummy [87],\$dummy [88],\$dummy [89],\$dummy [90],
                  \$dummy [91],\$dummy [92],\$dummy [93],\$dummy [94],
                  \$dummy [95]})) ;
    Multiplier_16 loop3_6_Multip (.A ({FilterToAlu_111,FilterToAlu_110,
                  FilterToAlu_109,FilterToAlu_108,FilterToAlu_107,
                  FilterToAlu_106,FilterToAlu_105,FilterToAlu_104,
                  FilterToAlu_103,FilterToAlu_102,FilterToAlu_101,
                  FilterToAlu_100,FilterToAlu_99,FilterToAlu_98,FilterToAlu_97,
                  FilterToAlu_96}), .B ({SecondInputToMult_111,
                  SecondInputToMult_110,SecondInputToMult_109,
                  SecondInputToMult_108,SecondInputToMult_107,
                  SecondInputToMult_106,SecondInputToMult_105,
                  SecondInputToMult_104,SecondInputToMult_103,
                  SecondInputToMult_102,SecondInputToMult_101,
                  SecondInputToMult_100,SecondInputToMult_99,
                  SecondInputToMult_98,SecondInputToMult_97,SecondInputToMult_96
                  }), .F ({\$dummy [96],\$dummy [97],\$dummy [98],\$dummy [99],
                  \$dummy [100],\$dummy [101],\$dummy [102],MultiplierOut_216,
                  MultiplierOut_215,MultiplierOut_214,MultiplierOut_213,
                  MultiplierOut_212,MultiplierOut_211,MultiplierOut_210,
                  MultiplierOut_209,MultiplierOut_208,MultiplierOut_207,
                  MultiplierOut_206,MultiplierOut_205,MultiplierOut_204,
                  MultiplierOut_203,MultiplierOut_202,MultiplierOut_201,
                  \$dummy [103],\$dummy [104],\$dummy [105],\$dummy [106],
                  \$dummy [107],\$dummy [108],\$dummy [109],\$dummy [110],
                  \$dummy [111]})) ;
    Multiplier_16 loop3_7_Multip (.A ({FilterToAlu_127,FilterToAlu_126,
                  FilterToAlu_125,FilterToAlu_124,FilterToAlu_123,
                  FilterToAlu_122,FilterToAlu_121,FilterToAlu_120,
                  FilterToAlu_119,FilterToAlu_118,FilterToAlu_117,
                  FilterToAlu_116,FilterToAlu_115,FilterToAlu_114,
                  FilterToAlu_113,FilterToAlu_112}), .B ({SecondInputToMult_127,
                  SecondInputToMult_126,SecondInputToMult_125,
                  SecondInputToMult_124,SecondInputToMult_123,
                  SecondInputToMult_122,SecondInputToMult_121,
                  SecondInputToMult_120,SecondInputToMult_119,
                  SecondInputToMult_118,SecondInputToMult_117,
                  SecondInputToMult_116,SecondInputToMult_115,
                  SecondInputToMult_114,SecondInputToMult_113,
                  SecondInputToMult_112}), .F ({\$dummy [112],\$dummy [113],
                  \$dummy [114],\$dummy [115],\$dummy [116],\$dummy [117],
                  \$dummy [118],MultiplierOut_248,MultiplierOut_247,
                  MultiplierOut_246,MultiplierOut_245,MultiplierOut_244,
                  MultiplierOut_243,MultiplierOut_242,MultiplierOut_241,
                  MultiplierOut_240,MultiplierOut_239,MultiplierOut_238,
                  MultiplierOut_237,MultiplierOut_236,MultiplierOut_235,
                  MultiplierOut_234,MultiplierOut_233,\$dummy [119],
                  \$dummy [120],\$dummy [121],\$dummy [122],\$dummy [123],
                  \$dummy [124],\$dummy [125],\$dummy [126],\$dummy [127]})) ;
    Multiplier_16 loop3_8_Multip (.A ({FilterToAlu_143,FilterToAlu_142,
                  FilterToAlu_141,FilterToAlu_140,FilterToAlu_139,
                  FilterToAlu_138,FilterToAlu_137,FilterToAlu_136,
                  FilterToAlu_135,FilterToAlu_134,FilterToAlu_133,
                  FilterToAlu_132,FilterToAlu_131,FilterToAlu_130,
                  FilterToAlu_129,FilterToAlu_128}), .B ({SecondInputToMult_143,
                  SecondInputToMult_142,SecondInputToMult_141,
                  SecondInputToMult_140,SecondInputToMult_139,
                  SecondInputToMult_138,SecondInputToMult_137,
                  SecondInputToMult_136,SecondInputToMult_135,
                  SecondInputToMult_134,SecondInputToMult_133,
                  SecondInputToMult_132,SecondInputToMult_131,
                  SecondInputToMult_130,SecondInputToMult_129,
                  SecondInputToMult_128}), .F ({\$dummy [128],\$dummy [129],
                  \$dummy [130],\$dummy [131],\$dummy [132],\$dummy [133],
                  \$dummy [134],MultiplierOut_280,MultiplierOut_279,
                  MultiplierOut_278,MultiplierOut_277,MultiplierOut_276,
                  MultiplierOut_275,MultiplierOut_274,MultiplierOut_273,
                  MultiplierOut_272,MultiplierOut_271,MultiplierOut_270,
                  MultiplierOut_269,MultiplierOut_268,MultiplierOut_267,
                  MultiplierOut_266,MultiplierOut_265,\$dummy [135],
                  \$dummy [136],\$dummy [137],\$dummy [138],\$dummy [139],
                  \$dummy [140],\$dummy [141],\$dummy [142],\$dummy [143]})) ;
    Multiplier_16 loop5_9_Multip (.A ({FilterToAlu_159,FilterToAlu_158,
                  FilterToAlu_157,FilterToAlu_156,FilterToAlu_155,
                  FilterToAlu_154,FilterToAlu_153,FilterToAlu_152,
                  FilterToAlu_151,FilterToAlu_150,FilterToAlu_149,
                  FilterToAlu_148,FilterToAlu_147,FilterToAlu_146,
                  FilterToAlu_145,FilterToAlu_144}), .B ({OutputImg1[79],
                  OutputImg1[78],OutputImg1[77],OutputImg1[76],OutputImg1[75],
                  OutputImg1[74],OutputImg1[73],OutputImg1[72],OutputImg1[71],
                  OutputImg1[70],OutputImg1[69],OutputImg1[68],OutputImg1[67],
                  OutputImg1[66],OutputImg1[65],OutputImg1[64]}), .F ({
                  \$dummy [144],\$dummy [145],\$dummy [146],\$dummy [147],
                  \$dummy [148],\$dummy [149],\$dummy [150],MultiplierOut_312,
                  MultiplierOut_311,MultiplierOut_310,MultiplierOut_309,
                  MultiplierOut_308,MultiplierOut_307,MultiplierOut_306,
                  MultiplierOut_305,MultiplierOut_304,MultiplierOut_303,
                  MultiplierOut_302,MultiplierOut_301,MultiplierOut_300,
                  MultiplierOut_299,MultiplierOut_298,MultiplierOut_297,
                  \$dummy [151],\$dummy [152],\$dummy [153],\$dummy [154],
                  \$dummy [155],\$dummy [156],\$dummy [157],\$dummy [158],
                  \$dummy [159]})) ;
    Multiplier_16 loop5_10_Multip (.A ({FilterToAlu_175,FilterToAlu_174,
                  FilterToAlu_173,FilterToAlu_172,FilterToAlu_171,
                  FilterToAlu_170,FilterToAlu_169,FilterToAlu_168,
                  FilterToAlu_167,FilterToAlu_166,FilterToAlu_165,
                  FilterToAlu_164,FilterToAlu_163,FilterToAlu_162,
                  FilterToAlu_161,FilterToAlu_160}), .B ({OutputImg2[15],
                  OutputImg2[14],OutputImg2[13],OutputImg2[12],OutputImg2[11],
                  OutputImg2[10],OutputImg2[9],OutputImg2[8],OutputImg2[7],
                  OutputImg2[6],OutputImg2[5],OutputImg2[4],OutputImg2[3],
                  OutputImg2[2],OutputImg2[1],OutputImg2[0]}), .F ({
                  \$dummy [160],\$dummy [161],\$dummy [162],\$dummy [163],
                  \$dummy [164],\$dummy [165],\$dummy [166],MultiplierOut_344,
                  MultiplierOut_343,MultiplierOut_342,MultiplierOut_341,
                  MultiplierOut_340,MultiplierOut_339,MultiplierOut_338,
                  MultiplierOut_337,MultiplierOut_336,MultiplierOut_335,
                  MultiplierOut_334,MultiplierOut_333,MultiplierOut_332,
                  MultiplierOut_331,MultiplierOut_330,MultiplierOut_329,
                  \$dummy [167],\$dummy [168],\$dummy [169],\$dummy [170],
                  \$dummy [171],\$dummy [172],\$dummy [173],\$dummy [174],
                  \$dummy [175]})) ;
    Multiplier_16 loop5_11_Multip (.A ({FilterToAlu_191,FilterToAlu_190,
                  FilterToAlu_189,FilterToAlu_188,FilterToAlu_187,
                  FilterToAlu_186,FilterToAlu_185,FilterToAlu_184,
                  FilterToAlu_183,FilterToAlu_182,FilterToAlu_181,
                  FilterToAlu_180,FilterToAlu_179,FilterToAlu_178,
                  FilterToAlu_177,FilterToAlu_176}), .B ({OutputImg2[31],
                  OutputImg2[30],OutputImg2[29],OutputImg2[28],OutputImg2[27],
                  OutputImg2[26],OutputImg2[25],OutputImg2[24],OutputImg2[23],
                  OutputImg2[22],OutputImg2[21],OutputImg2[20],OutputImg2[19],
                  OutputImg2[18],OutputImg2[17],OutputImg2[16]}), .F ({
                  \$dummy [176],\$dummy [177],\$dummy [178],\$dummy [179],
                  \$dummy [180],\$dummy [181],\$dummy [182],MultiplierOut_376,
                  MultiplierOut_375,MultiplierOut_374,MultiplierOut_373,
                  MultiplierOut_372,MultiplierOut_371,MultiplierOut_370,
                  MultiplierOut_369,MultiplierOut_368,MultiplierOut_367,
                  MultiplierOut_366,MultiplierOut_365,MultiplierOut_364,
                  MultiplierOut_363,MultiplierOut_362,MultiplierOut_361,
                  \$dummy [183],\$dummy [184],\$dummy [185],\$dummy [186],
                  \$dummy [187],\$dummy [188],\$dummy [189],\$dummy [190],
                  \$dummy [191]})) ;
    Multiplier_16 loop5_12_Multip (.A ({FilterToAlu_207,FilterToAlu_206,
                  FilterToAlu_205,FilterToAlu_204,FilterToAlu_203,
                  FilterToAlu_202,FilterToAlu_201,FilterToAlu_200,
                  FilterToAlu_199,FilterToAlu_198,FilterToAlu_197,
                  FilterToAlu_196,FilterToAlu_195,FilterToAlu_194,
                  FilterToAlu_193,FilterToAlu_192}), .B ({OutputImg2[47],
                  OutputImg2[46],OutputImg2[45],OutputImg2[44],OutputImg2[43],
                  OutputImg2[42],OutputImg2[41],OutputImg2[40],OutputImg2[39],
                  OutputImg2[38],OutputImg2[37],OutputImg2[36],OutputImg2[35],
                  OutputImg2[34],OutputImg2[33],OutputImg2[32]}), .F ({
                  \$dummy [192],\$dummy [193],\$dummy [194],\$dummy [195],
                  \$dummy [196],\$dummy [197],\$dummy [198],MultiplierOut_408,
                  MultiplierOut_407,MultiplierOut_406,MultiplierOut_405,
                  MultiplierOut_404,MultiplierOut_403,MultiplierOut_402,
                  MultiplierOut_401,MultiplierOut_400,MultiplierOut_399,
                  MultiplierOut_398,MultiplierOut_397,MultiplierOut_396,
                  MultiplierOut_395,MultiplierOut_394,MultiplierOut_393,
                  \$dummy [199],\$dummy [200],\$dummy [201],\$dummy [202],
                  \$dummy [203],\$dummy [204],\$dummy [205],\$dummy [206],
                  \$dummy [207]})) ;
    Multiplier_16 loop5_13_Multip (.A ({FilterToAlu_223,FilterToAlu_222,
                  FilterToAlu_221,FilterToAlu_220,FilterToAlu_219,
                  FilterToAlu_218,FilterToAlu_217,FilterToAlu_216,
                  FilterToAlu_215,FilterToAlu_214,FilterToAlu_213,
                  FilterToAlu_212,FilterToAlu_211,FilterToAlu_210,
                  FilterToAlu_209,FilterToAlu_208}), .B ({OutputImg2[63],
                  OutputImg2[62],OutputImg2[61],OutputImg2[60],OutputImg2[59],
                  OutputImg2[58],OutputImg2[57],OutputImg2[56],OutputImg2[55],
                  OutputImg2[54],OutputImg2[53],OutputImg2[52],OutputImg2[51],
                  OutputImg2[50],OutputImg2[49],OutputImg2[48]}), .F ({
                  \$dummy [208],\$dummy [209],\$dummy [210],\$dummy [211],
                  \$dummy [212],\$dummy [213],\$dummy [214],MultiplierOut_440,
                  MultiplierOut_439,MultiplierOut_438,MultiplierOut_437,
                  MultiplierOut_436,MultiplierOut_435,MultiplierOut_434,
                  MultiplierOut_433,MultiplierOut_432,MultiplierOut_431,
                  MultiplierOut_430,MultiplierOut_429,MultiplierOut_428,
                  MultiplierOut_427,MultiplierOut_426,MultiplierOut_425,
                  \$dummy [215],\$dummy [216],\$dummy [217],\$dummy [218],
                  \$dummy [219],\$dummy [220],\$dummy [221],\$dummy [222],
                  \$dummy [223]})) ;
    Multiplier_16 loop5_14_Multip (.A ({FilterToAlu_239,FilterToAlu_238,
                  FilterToAlu_237,FilterToAlu_236,FilterToAlu_235,
                  FilterToAlu_234,FilterToAlu_233,FilterToAlu_232,
                  FilterToAlu_231,FilterToAlu_230,FilterToAlu_229,
                  FilterToAlu_228,FilterToAlu_227,FilterToAlu_226,
                  FilterToAlu_225,FilterToAlu_224}), .B ({OutputImg2[79],
                  OutputImg2[78],OutputImg2[77],OutputImg2[76],OutputImg2[75],
                  OutputImg2[74],OutputImg2[73],OutputImg2[72],OutputImg2[71],
                  OutputImg2[70],OutputImg2[69],OutputImg2[68],OutputImg2[67],
                  OutputImg2[66],OutputImg2[65],OutputImg2[64]}), .F ({
                  \$dummy [224],\$dummy [225],\$dummy [226],\$dummy [227],
                  \$dummy [228],\$dummy [229],\$dummy [230],MultiplierOut_472,
                  MultiplierOut_471,MultiplierOut_470,MultiplierOut_469,
                  MultiplierOut_468,MultiplierOut_467,MultiplierOut_466,
                  MultiplierOut_465,MultiplierOut_464,MultiplierOut_463,
                  MultiplierOut_462,MultiplierOut_461,MultiplierOut_460,
                  MultiplierOut_459,MultiplierOut_458,MultiplierOut_457,
                  \$dummy [231],\$dummy [232],\$dummy [233],\$dummy [234],
                  \$dummy [235],\$dummy [236],\$dummy [237],\$dummy [238],
                  \$dummy [239]})) ;
    Multiplier_16 loop5_15_Multip (.A ({FilterToAlu_255,FilterToAlu_254,
                  FilterToAlu_253,FilterToAlu_252,FilterToAlu_251,
                  FilterToAlu_250,FilterToAlu_249,FilterToAlu_248,
                  FilterToAlu_247,FilterToAlu_246,FilterToAlu_245,
                  FilterToAlu_244,FilterToAlu_243,FilterToAlu_242,
                  FilterToAlu_241,FilterToAlu_240}), .B ({OutputImg3[15],
                  OutputImg3[14],OutputImg3[13],OutputImg3[12],OutputImg3[11],
                  OutputImg3[10],OutputImg3[9],OutputImg3[8],OutputImg3[7],
                  OutputImg3[6],OutputImg3[5],OutputImg3[4],OutputImg3[3],
                  OutputImg3[2],OutputImg3[1],OutputImg3[0]}), .F ({
                  \$dummy [240],\$dummy [241],\$dummy [242],\$dummy [243],
                  \$dummy [244],\$dummy [245],\$dummy [246],MultiplierOut_504,
                  MultiplierOut_503,MultiplierOut_502,MultiplierOut_501,
                  MultiplierOut_500,MultiplierOut_499,MultiplierOut_498,
                  MultiplierOut_497,MultiplierOut_496,MultiplierOut_495,
                  MultiplierOut_494,MultiplierOut_493,MultiplierOut_492,
                  MultiplierOut_491,MultiplierOut_490,MultiplierOut_489,
                  \$dummy [247],\$dummy [248],\$dummy [249],\$dummy [250],
                  \$dummy [251],\$dummy [252],\$dummy [253],\$dummy [254],
                  \$dummy [255]})) ;
    Multiplier_16 loop5_16_Multip (.A ({FilterToAlu_271,FilterToAlu_270,
                  FilterToAlu_269,FilterToAlu_268,FilterToAlu_267,
                  FilterToAlu_266,FilterToAlu_265,FilterToAlu_264,
                  FilterToAlu_263,FilterToAlu_262,FilterToAlu_261,
                  FilterToAlu_260,FilterToAlu_259,FilterToAlu_258,
                  FilterToAlu_257,FilterToAlu_256}), .B ({OutputImg3[31],
                  OutputImg3[30],OutputImg3[29],OutputImg3[28],OutputImg3[27],
                  OutputImg3[26],OutputImg3[25],OutputImg3[24],OutputImg3[23],
                  OutputImg3[22],OutputImg3[21],OutputImg3[20],OutputImg3[19],
                  OutputImg3[18],OutputImg3[17],OutputImg3[16]}), .F ({
                  \$dummy [256],\$dummy [257],\$dummy [258],\$dummy [259],
                  \$dummy [260],\$dummy [261],\$dummy [262],MultiplierOut_536,
                  MultiplierOut_535,MultiplierOut_534,MultiplierOut_533,
                  MultiplierOut_532,MultiplierOut_531,MultiplierOut_530,
                  MultiplierOut_529,MultiplierOut_528,MultiplierOut_527,
                  MultiplierOut_526,MultiplierOut_525,MultiplierOut_524,
                  MultiplierOut_523,MultiplierOut_522,MultiplierOut_521,
                  \$dummy [263],\$dummy [264],\$dummy [265],\$dummy [266],
                  \$dummy [267],\$dummy [268],\$dummy [269],\$dummy [270],
                  \$dummy [271]})) ;
    Multiplier_16 loop5_17_Multip (.A ({FilterToAlu_287,FilterToAlu_286,
                  FilterToAlu_285,FilterToAlu_284,FilterToAlu_283,
                  FilterToAlu_282,FilterToAlu_281,FilterToAlu_280,
                  FilterToAlu_279,FilterToAlu_278,FilterToAlu_277,
                  FilterToAlu_276,FilterToAlu_275,FilterToAlu_274,
                  FilterToAlu_273,FilterToAlu_272}), .B ({OutputImg3[47],
                  OutputImg3[46],OutputImg3[45],OutputImg3[44],OutputImg3[43],
                  OutputImg3[42],OutputImg3[41],OutputImg3[40],OutputImg3[39],
                  OutputImg3[38],OutputImg3[37],OutputImg3[36],OutputImg3[35],
                  OutputImg3[34],OutputImg3[33],OutputImg3[32]}), .F ({
                  \$dummy [272],\$dummy [273],\$dummy [274],\$dummy [275],
                  \$dummy [276],\$dummy [277],\$dummy [278],MultiplierOut_568,
                  MultiplierOut_567,MultiplierOut_566,MultiplierOut_565,
                  MultiplierOut_564,MultiplierOut_563,MultiplierOut_562,
                  MultiplierOut_561,MultiplierOut_560,MultiplierOut_559,
                  MultiplierOut_558,MultiplierOut_557,MultiplierOut_556,
                  MultiplierOut_555,MultiplierOut_554,MultiplierOut_553,
                  \$dummy [279],\$dummy [280],\$dummy [281],\$dummy [282],
                  \$dummy [283],\$dummy [284],\$dummy [285],\$dummy [286],
                  \$dummy [287]})) ;
    Multiplier_16 loop5_18_Multip (.A ({FilterToAlu_303,FilterToAlu_302,
                  FilterToAlu_301,FilterToAlu_300,FilterToAlu_299,
                  FilterToAlu_298,FilterToAlu_297,FilterToAlu_296,
                  FilterToAlu_295,FilterToAlu_294,FilterToAlu_293,
                  FilterToAlu_292,FilterToAlu_291,FilterToAlu_290,
                  FilterToAlu_289,FilterToAlu_288}), .B ({OutputImg3[63],
                  OutputImg3[62],OutputImg3[61],OutputImg3[60],OutputImg3[59],
                  OutputImg3[58],OutputImg3[57],OutputImg3[56],OutputImg3[55],
                  OutputImg3[54],OutputImg3[53],OutputImg3[52],OutputImg3[51],
                  OutputImg3[50],OutputImg3[49],OutputImg3[48]}), .F ({
                  \$dummy [288],\$dummy [289],\$dummy [290],\$dummy [291],
                  \$dummy [292],\$dummy [293],\$dummy [294],MultiplierOut_600,
                  MultiplierOut_599,MultiplierOut_598,MultiplierOut_597,
                  MultiplierOut_596,MultiplierOut_595,MultiplierOut_594,
                  MultiplierOut_593,MultiplierOut_592,MultiplierOut_591,
                  MultiplierOut_590,MultiplierOut_589,MultiplierOut_588,
                  MultiplierOut_587,MultiplierOut_586,MultiplierOut_585,
                  \$dummy [295],\$dummy [296],\$dummy [297],\$dummy [298],
                  \$dummy [299],\$dummy [300],\$dummy [301],\$dummy [302],
                  \$dummy [303]})) ;
    Multiplier_16 loop5_19_Multip (.A ({FilterToAlu_319,FilterToAlu_318,
                  FilterToAlu_317,FilterToAlu_316,FilterToAlu_315,
                  FilterToAlu_314,FilterToAlu_313,FilterToAlu_312,
                  FilterToAlu_311,FilterToAlu_310,FilterToAlu_309,
                  FilterToAlu_308,FilterToAlu_307,FilterToAlu_306,
                  FilterToAlu_305,FilterToAlu_304}), .B ({OutputImg3[79],
                  OutputImg3[78],OutputImg3[77],OutputImg3[76],OutputImg3[75],
                  OutputImg3[74],OutputImg3[73],OutputImg3[72],OutputImg3[71],
                  OutputImg3[70],OutputImg3[69],OutputImg3[68],OutputImg3[67],
                  OutputImg3[66],OutputImg3[65],OutputImg3[64]}), .F ({
                  \$dummy [304],\$dummy [305],\$dummy [306],\$dummy [307],
                  \$dummy [308],\$dummy [309],\$dummy [310],MultiplierOut_632,
                  MultiplierOut_631,MultiplierOut_630,MultiplierOut_629,
                  MultiplierOut_628,MultiplierOut_627,MultiplierOut_626,
                  MultiplierOut_625,MultiplierOut_624,MultiplierOut_623,
                  MultiplierOut_622,MultiplierOut_621,MultiplierOut_620,
                  MultiplierOut_619,MultiplierOut_618,MultiplierOut_617,
                  \$dummy [311],\$dummy [312],\$dummy [313],\$dummy [314],
                  \$dummy [315],\$dummy [316],\$dummy [317],\$dummy [318],
                  \$dummy [319]})) ;
    Multiplier_16 loop5_20_Multip (.A ({FilterToAlu_335,FilterToAlu_334,
                  FilterToAlu_333,FilterToAlu_332,FilterToAlu_331,
                  FilterToAlu_330,FilterToAlu_329,FilterToAlu_328,
                  FilterToAlu_327,FilterToAlu_326,FilterToAlu_325,
                  FilterToAlu_324,FilterToAlu_323,FilterToAlu_322,
                  FilterToAlu_321,FilterToAlu_320}), .B ({OutputImg4[15],
                  OutputImg4[14],OutputImg4[13],OutputImg4[12],OutputImg4[11],
                  OutputImg4[10],OutputImg4[9],OutputImg4[8],OutputImg4[7],
                  OutputImg4[6],OutputImg4[5],OutputImg4[4],OutputImg4[3],
                  OutputImg4[2],OutputImg4[1],OutputImg4[0]}), .F ({
                  \$dummy [320],\$dummy [321],\$dummy [322],\$dummy [323],
                  \$dummy [324],\$dummy [325],\$dummy [326],MultiplierOut_664,
                  MultiplierOut_663,MultiplierOut_662,MultiplierOut_661,
                  MultiplierOut_660,MultiplierOut_659,MultiplierOut_658,
                  MultiplierOut_657,MultiplierOut_656,MultiplierOut_655,
                  MultiplierOut_654,MultiplierOut_653,MultiplierOut_652,
                  MultiplierOut_651,MultiplierOut_650,MultiplierOut_649,
                  \$dummy [327],\$dummy [328],\$dummy [329],\$dummy [330],
                  \$dummy [331],\$dummy [332],\$dummy [333],\$dummy [334],
                  \$dummy [335]})) ;
    Multiplier_16 loop5_21_Multip (.A ({FilterToAlu_351,FilterToAlu_350,
                  FilterToAlu_349,FilterToAlu_348,FilterToAlu_347,
                  FilterToAlu_346,FilterToAlu_345,FilterToAlu_344,
                  FilterToAlu_343,FilterToAlu_342,FilterToAlu_341,
                  FilterToAlu_340,FilterToAlu_339,FilterToAlu_338,
                  FilterToAlu_337,FilterToAlu_336}), .B ({OutputImg4[31],
                  OutputImg4[30],OutputImg4[29],OutputImg4[28],OutputImg4[27],
                  OutputImg4[26],OutputImg4[25],OutputImg4[24],OutputImg4[23],
                  OutputImg4[22],OutputImg4[21],OutputImg4[20],OutputImg4[19],
                  OutputImg4[18],OutputImg4[17],OutputImg4[16]}), .F ({
                  \$dummy [336],\$dummy [337],\$dummy [338],\$dummy [339],
                  \$dummy [340],\$dummy [341],\$dummy [342],MultiplierOut_696,
                  MultiplierOut_695,MultiplierOut_694,MultiplierOut_693,
                  MultiplierOut_692,MultiplierOut_691,MultiplierOut_690,
                  MultiplierOut_689,MultiplierOut_688,MultiplierOut_687,
                  MultiplierOut_686,MultiplierOut_685,MultiplierOut_684,
                  MultiplierOut_683,MultiplierOut_682,MultiplierOut_681,
                  \$dummy [343],\$dummy [344],\$dummy [345],\$dummy [346],
                  \$dummy [347],\$dummy [348],\$dummy [349],\$dummy [350],
                  \$dummy [351]})) ;
    Multiplier_16 loop5_22_Multip (.A ({FilterToAlu_367,FilterToAlu_366,
                  FilterToAlu_365,FilterToAlu_364,FilterToAlu_363,
                  FilterToAlu_362,FilterToAlu_361,FilterToAlu_360,
                  FilterToAlu_359,FilterToAlu_358,FilterToAlu_357,
                  FilterToAlu_356,FilterToAlu_355,FilterToAlu_354,
                  FilterToAlu_353,FilterToAlu_352}), .B ({OutputImg4[47],
                  OutputImg4[46],OutputImg4[45],OutputImg4[44],OutputImg4[43],
                  OutputImg4[42],OutputImg4[41],OutputImg4[40],OutputImg4[39],
                  OutputImg4[38],OutputImg4[37],OutputImg4[36],OutputImg4[35],
                  OutputImg4[34],OutputImg4[33],OutputImg4[32]}), .F ({
                  \$dummy [352],\$dummy [353],\$dummy [354],\$dummy [355],
                  \$dummy [356],\$dummy [357],\$dummy [358],MultiplierOut_728,
                  MultiplierOut_727,MultiplierOut_726,MultiplierOut_725,
                  MultiplierOut_724,MultiplierOut_723,MultiplierOut_722,
                  MultiplierOut_721,MultiplierOut_720,MultiplierOut_719,
                  MultiplierOut_718,MultiplierOut_717,MultiplierOut_716,
                  MultiplierOut_715,MultiplierOut_714,MultiplierOut_713,
                  \$dummy [359],\$dummy [360],\$dummy [361],\$dummy [362],
                  \$dummy [363],\$dummy [364],\$dummy [365],\$dummy [366],
                  \$dummy [367]})) ;
    Multiplier_16 loop5_23_Multip (.A ({FilterToAlu_383,FilterToAlu_382,
                  FilterToAlu_381,FilterToAlu_380,FilterToAlu_379,
                  FilterToAlu_378,FilterToAlu_377,FilterToAlu_376,
                  FilterToAlu_375,FilterToAlu_374,FilterToAlu_373,
                  FilterToAlu_372,FilterToAlu_371,FilterToAlu_370,
                  FilterToAlu_369,FilterToAlu_368}), .B ({OutputImg4[63],
                  OutputImg4[62],OutputImg4[61],OutputImg4[60],OutputImg4[59],
                  OutputImg4[58],OutputImg4[57],OutputImg4[56],OutputImg4[55],
                  OutputImg4[54],OutputImg4[53],OutputImg4[52],OutputImg4[51],
                  OutputImg4[50],OutputImg4[49],OutputImg4[48]}), .F ({
                  \$dummy [368],\$dummy [369],\$dummy [370],\$dummy [371],
                  \$dummy [372],\$dummy [373],\$dummy [374],MultiplierOut_760,
                  MultiplierOut_759,MultiplierOut_758,MultiplierOut_757,
                  MultiplierOut_756,MultiplierOut_755,MultiplierOut_754,
                  MultiplierOut_753,MultiplierOut_752,MultiplierOut_751,
                  MultiplierOut_750,MultiplierOut_749,MultiplierOut_748,
                  MultiplierOut_747,MultiplierOut_746,MultiplierOut_745,
                  \$dummy [375],\$dummy [376],\$dummy [377],\$dummy [378],
                  \$dummy [379],\$dummy [380],\$dummy [381],\$dummy [382],
                  \$dummy [383]})) ;
    Multiplier_16 loop5_24_Multip (.A ({FilterToAlu_399,FilterToAlu_398,
                  FilterToAlu_397,FilterToAlu_396,FilterToAlu_395,
                  FilterToAlu_394,FilterToAlu_393,FilterToAlu_392,
                  FilterToAlu_391,FilterToAlu_390,FilterToAlu_389,
                  FilterToAlu_388,FilterToAlu_387,FilterToAlu_386,
                  FilterToAlu_385,FilterToAlu_384}), .B ({OutputImg4[79],
                  OutputImg4[78],OutputImg4[77],OutputImg4[76],OutputImg4[75],
                  OutputImg4[74],OutputImg4[73],OutputImg4[72],OutputImg4[71],
                  OutputImg4[70],OutputImg4[69],OutputImg4[68],OutputImg4[67],
                  OutputImg4[66],OutputImg4[65],OutputImg4[64]}), .F ({
                  \$dummy [384],\$dummy [385],\$dummy [386],\$dummy [387],
                  \$dummy [388],\$dummy [389],\$dummy [390],MultiplierOut_792,
                  MultiplierOut_791,MultiplierOut_790,MultiplierOut_789,
                  MultiplierOut_788,MultiplierOut_787,MultiplierOut_786,
                  MultiplierOut_785,MultiplierOut_784,MultiplierOut_783,
                  MultiplierOut_782,MultiplierOut_781,MultiplierOut_780,
                  MultiplierOut_779,MultiplierOut_778,MultiplierOut_777,
                  \$dummy [391],\$dummy [392],\$dummy [393],\$dummy [394],
                  \$dummy [395],\$dummy [396],\$dummy [397],\$dummy [398],
                  \$dummy [399]})) ;
    my_nadder_16 adder1 (.a ({MultiplierOut_24,MultiplierOut_23,MultiplierOut_22
                 ,MultiplierOut_21,MultiplierOut_20,MultiplierOut_19,
                 MultiplierOut_18,MultiplierOut_17,MultiplierOut_16,
                 MultiplierOut_15,MultiplierOut_14,MultiplierOut_13,
                 MultiplierOut_12,MultiplierOut_11,MultiplierOut_10,
                 MultiplierOut_9}), .b ({MultiplierOut_56,MultiplierOut_55,
                 MultiplierOut_54,MultiplierOut_53,MultiplierOut_52,
                 MultiplierOut_51,MultiplierOut_50,MultiplierOut_49,
                 MultiplierOut_48,MultiplierOut_47,MultiplierOut_46,
                 MultiplierOut_45,MultiplierOut_44,MultiplierOut_43,
                 MultiplierOut_42,MultiplierOut_41}), .cin (GND0), .s ({
                 AddOutputLvL1_15,AddOutputLvL1_14,AddOutputLvL1_13,
                 AddOutputLvL1_12,AddOutputLvL1_11,AddOutputLvL1_10,
                 AddOutputLvL1_9,AddOutputLvL1_8,AddOutputLvL1_7,AddOutputLvL1_6
                 ,AddOutputLvL1_5,AddOutputLvL1_4,AddOutputLvL1_3,
                 AddOutputLvL1_2,AddOutputLvL1_1,AddOutputLvL1_0}), .cout (
                 \$dummy [400])) ;
    my_nadder_16 adder2 (.a ({MultiplierOut_88,MultiplierOut_87,MultiplierOut_86
                 ,MultiplierOut_85,MultiplierOut_84,MultiplierOut_83,
                 MultiplierOut_82,MultiplierOut_81,MultiplierOut_80,
                 MultiplierOut_79,MultiplierOut_78,MultiplierOut_77,
                 MultiplierOut_76,MultiplierOut_75,MultiplierOut_74,
                 MultiplierOut_73}), .b ({MultiplierOut_120,MultiplierOut_119,
                 MultiplierOut_118,MultiplierOut_117,MultiplierOut_116,
                 MultiplierOut_115,MultiplierOut_114,MultiplierOut_113,
                 MultiplierOut_112,MultiplierOut_111,MultiplierOut_110,
                 MultiplierOut_109,MultiplierOut_108,MultiplierOut_107,
                 MultiplierOut_106,MultiplierOut_105}), .cin (GND0), .s ({
                 AddOutputLvL1_31,AddOutputLvL1_30,AddOutputLvL1_29,
                 AddOutputLvL1_28,AddOutputLvL1_27,AddOutputLvL1_26,
                 AddOutputLvL1_25,AddOutputLvL1_24,AddOutputLvL1_23,
                 AddOutputLvL1_22,AddOutputLvL1_21,AddOutputLvL1_20,
                 AddOutputLvL1_19,AddOutputLvL1_18,AddOutputLvL1_17,
                 AddOutputLvL1_16}), .cout (\$dummy [401])) ;
    my_nadder_16 adder3 (.a ({MultiplierOut_152,MultiplierOut_151,
                 MultiplierOut_150,MultiplierOut_149,MultiplierOut_148,
                 MultiplierOut_147,MultiplierOut_146,MultiplierOut_145,
                 MultiplierOut_144,MultiplierOut_143,MultiplierOut_142,
                 MultiplierOut_141,MultiplierOut_140,MultiplierOut_139,
                 MultiplierOut_138,MultiplierOut_137}), .b ({MultiplierOut_184,
                 MultiplierOut_183,MultiplierOut_182,MultiplierOut_181,
                 MultiplierOut_180,MultiplierOut_179,MultiplierOut_178,
                 MultiplierOut_177,MultiplierOut_176,MultiplierOut_175,
                 MultiplierOut_174,MultiplierOut_173,MultiplierOut_172,
                 MultiplierOut_171,MultiplierOut_170,MultiplierOut_169}), .cin (
                 GND0), .s ({AddOutputLvL1_47,AddOutputLvL1_46,AddOutputLvL1_45,
                 AddOutputLvL1_44,AddOutputLvL1_43,AddOutputLvL1_42,
                 AddOutputLvL1_41,AddOutputLvL1_40,AddOutputLvL1_39,
                 AddOutputLvL1_38,AddOutputLvL1_37,AddOutputLvL1_36,
                 AddOutputLvL1_35,AddOutputLvL1_34,AddOutputLvL1_33,
                 AddOutputLvL1_32}), .cout (\$dummy [402])) ;
    my_nadder_16 adder4 (.a ({MultiplierOut_216,MultiplierOut_215,
                 MultiplierOut_214,MultiplierOut_213,MultiplierOut_212,
                 MultiplierOut_211,MultiplierOut_210,MultiplierOut_209,
                 MultiplierOut_208,MultiplierOut_207,MultiplierOut_206,
                 MultiplierOut_205,MultiplierOut_204,MultiplierOut_203,
                 MultiplierOut_202,MultiplierOut_201}), .b ({MultiplierOut_248,
                 MultiplierOut_247,MultiplierOut_246,MultiplierOut_245,
                 MultiplierOut_244,MultiplierOut_243,MultiplierOut_242,
                 MultiplierOut_241,MultiplierOut_240,MultiplierOut_239,
                 MultiplierOut_238,MultiplierOut_237,MultiplierOut_236,
                 MultiplierOut_235,MultiplierOut_234,MultiplierOut_233}), .cin (
                 GND0), .s ({AddOutputLvL1_63,AddOutputLvL1_62,AddOutputLvL1_61,
                 AddOutputLvL1_60,AddOutputLvL1_59,AddOutputLvL1_58,
                 AddOutputLvL1_57,AddOutputLvL1_56,AddOutputLvL1_55,
                 AddOutputLvL1_54,AddOutputLvL1_53,AddOutputLvL1_52,
                 AddOutputLvL1_51,AddOutputLvL1_50,AddOutputLvL1_49,
                 AddOutputLvL1_48}), .cout (\$dummy [403])) ;
    my_nadder_16 adder12 (.a ({AddOutputLvL1_15,AddOutputLvL1_14,
                 AddOutputLvL1_13,AddOutputLvL1_12,AddOutputLvL1_11,
                 AddOutputLvL1_10,AddOutputLvL1_9,AddOutputLvL1_8,
                 AddOutputLvL1_7,AddOutputLvL1_6,AddOutputLvL1_5,AddOutputLvL1_4
                 ,AddOutputLvL1_3,AddOutputLvL1_2,AddOutputLvL1_1,
                 AddOutputLvL1_0}), .b ({AddOutputLvL1_31,AddOutputLvL1_30,
                 AddOutputLvL1_29,AddOutputLvL1_28,AddOutputLvL1_27,
                 AddOutputLvL1_26,AddOutputLvL1_25,AddOutputLvL1_24,
                 AddOutputLvL1_23,AddOutputLvL1_22,AddOutputLvL1_21,
                 AddOutputLvL1_20,AddOutputLvL1_19,AddOutputLvL1_18,
                 AddOutputLvL1_17,AddOutputLvL1_16}), .cin (GND0), .s ({
                 AddOutputLvL2_15,AddOutputLvL2_14,AddOutputLvL2_13,
                 AddOutputLvL2_12,AddOutputLvL2_11,AddOutputLvL2_10,
                 AddOutputLvL2_9,AddOutputLvL2_8,AddOutputLvL2_7,AddOutputLvL2_6
                 ,AddOutputLvL2_5,AddOutputLvL2_4,AddOutputLvL2_3,
                 AddOutputLvL2_2,AddOutputLvL2_1,AddOutputLvL2_0}), .cout (
                 \$dummy [404])) ;
    my_nadder_16 adder13 (.a ({AddOutputLvL1_47,AddOutputLvL1_46,
                 AddOutputLvL1_45,AddOutputLvL1_44,AddOutputLvL1_43,
                 AddOutputLvL1_42,AddOutputLvL1_41,AddOutputLvL1_40,
                 AddOutputLvL1_39,AddOutputLvL1_38,AddOutputLvL1_37,
                 AddOutputLvL1_36,AddOutputLvL1_35,AddOutputLvL1_34,
                 AddOutputLvL1_33,AddOutputLvL1_32}), .b ({AddOutputLvL1_63,
                 AddOutputLvL1_62,AddOutputLvL1_61,AddOutputLvL1_60,
                 AddOutputLvL1_59,AddOutputLvL1_58,AddOutputLvL1_57,
                 AddOutputLvL1_56,AddOutputLvL1_55,AddOutputLvL1_54,
                 AddOutputLvL1_53,AddOutputLvL1_52,AddOutputLvL1_51,
                 AddOutputLvL1_50,AddOutputLvL1_49,AddOutputLvL1_48}), .cin (
                 GND0), .s ({AddOutputLvL2_31,AddOutputLvL2_30,AddOutputLvL2_29,
                 AddOutputLvL2_28,AddOutputLvL2_27,AddOutputLvL2_26,
                 AddOutputLvL2_25,AddOutputLvL2_24,AddOutputLvL2_23,
                 AddOutputLvL2_22,AddOutputLvL2_21,AddOutputLvL2_20,
                 AddOutputLvL2_19,AddOutputLvL2_18,AddOutputLvL2_17,
                 AddOutputLvL2_16}), .cout (\$dummy [405])) ;
    my_nadder_16 adder18 (.a ({AddOutputLvL2_15,AddOutputLvL2_14,
                 AddOutputLvL2_13,AddOutputLvL2_12,AddOutputLvL2_11,
                 AddOutputLvL2_10,AddOutputLvL2_9,AddOutputLvL2_8,
                 AddOutputLvL2_7,AddOutputLvL2_6,AddOutputLvL2_5,AddOutputLvL2_4
                 ,AddOutputLvL2_3,AddOutputLvL2_2,AddOutputLvL2_1,
                 AddOutputLvL2_0}), .b ({AddOutputLvL2_31,AddOutputLvL2_30,
                 AddOutputLvL2_29,AddOutputLvL2_28,AddOutputLvL2_27,
                 AddOutputLvL2_26,AddOutputLvL2_25,AddOutputLvL2_24,
                 AddOutputLvL2_23,AddOutputLvL2_22,AddOutputLvL2_21,
                 AddOutputLvL2_20,AddOutputLvL2_19,AddOutputLvL2_18,
                 AddOutputLvL2_17,AddOutputLvL2_16}), .cin (GND0), .s ({
                 AddOutputLvL3_15,AddOutputLvL3_14,AddOutputLvL3_13,
                 AddOutputLvL3_12,AddOutputLvL3_11,AddOutputLvL3_10,
                 AddOutputLvL3_9,AddOutputLvL3_8,AddOutputLvL3_7,AddOutputLvL3_6
                 ,AddOutputLvL3_5,AddOutputLvL3_4,AddOutputLvL3_3,
                 AddOutputLvL3_2,AddOutputLvL3_1,AddOutputLvL3_0}), .cout (
                 \$dummy [406])) ;
    my_nadder_16 adder21 (.a ({AddOutputLvL3_15,AddOutputLvL3_14,
                 AddOutputLvL3_13,AddOutputLvL3_12,AddOutputLvL3_11,
                 AddOutputLvL3_10,AddOutputLvL3_9,AddOutputLvL3_8,
                 AddOutputLvL3_7,AddOutputLvL3_6,AddOutputLvL3_5,AddOutputLvL3_4
                 ,AddOutputLvL3_3,AddOutputLvL3_2,AddOutputLvL3_1,
                 AddOutputLvL3_0}), .b ({MultiplierOut_280,MultiplierOut_279,
                 MultiplierOut_278,MultiplierOut_277,MultiplierOut_276,
                 MultiplierOut_275,MultiplierOut_274,MultiplierOut_273,
                 MultiplierOut_272,MultiplierOut_271,MultiplierOut_270,
                 MultiplierOut_269,MultiplierOut_268,MultiplierOut_267,
                 MultiplierOut_266,MultiplierOut_265}), .cin (GND0), .s ({
                 AddOut33_15,AddOut33_14,AddOut33_13,AddOut33_12,AddOut33_11,
                 AddOut33_10,AddOut33_9,AddOut33_8,AddOut33_7,AddOut33_6,
                 AddOut33_5,AddOut33_4,AddOut33_3,AddOut33_2,AddOut33_1,
                 AddOut33_0}), .cout (\$dummy [407])) ;
    my_nadder_16 adder5 (.a ({MultiplierOut_312,MultiplierOut_311,
                 MultiplierOut_310,MultiplierOut_309,MultiplierOut_308,
                 MultiplierOut_307,MultiplierOut_306,MultiplierOut_305,
                 MultiplierOut_304,MultiplierOut_303,MultiplierOut_302,
                 MultiplierOut_301,MultiplierOut_300,MultiplierOut_299,
                 MultiplierOut_298,MultiplierOut_297}), .b ({MultiplierOut_344,
                 MultiplierOut_343,MultiplierOut_342,MultiplierOut_341,
                 MultiplierOut_340,MultiplierOut_339,MultiplierOut_338,
                 MultiplierOut_337,MultiplierOut_336,MultiplierOut_335,
                 MultiplierOut_334,MultiplierOut_333,MultiplierOut_332,
                 MultiplierOut_331,MultiplierOut_330,MultiplierOut_329}), .cin (
                 GND0), .s ({AddOutputLvL1_79,AddOutputLvL1_78,AddOutputLvL1_77,
                 AddOutputLvL1_76,AddOutputLvL1_75,AddOutputLvL1_74,
                 AddOutputLvL1_73,AddOutputLvL1_72,AddOutputLvL1_71,
                 AddOutputLvL1_70,AddOutputLvL1_69,AddOutputLvL1_68,
                 AddOutputLvL1_67,AddOutputLvL1_66,AddOutputLvL1_65,
                 AddOutputLvL1_64}), .cout (\$dummy [408])) ;
    my_nadder_16 adder6 (.a ({MultiplierOut_376,MultiplierOut_375,
                 MultiplierOut_374,MultiplierOut_373,MultiplierOut_372,
                 MultiplierOut_371,MultiplierOut_370,MultiplierOut_369,
                 MultiplierOut_368,MultiplierOut_367,MultiplierOut_366,
                 MultiplierOut_365,MultiplierOut_364,MultiplierOut_363,
                 MultiplierOut_362,MultiplierOut_361}), .b ({MultiplierOut_408,
                 MultiplierOut_407,MultiplierOut_406,MultiplierOut_405,
                 MultiplierOut_404,MultiplierOut_403,MultiplierOut_402,
                 MultiplierOut_401,MultiplierOut_400,MultiplierOut_399,
                 MultiplierOut_398,MultiplierOut_397,MultiplierOut_396,
                 MultiplierOut_395,MultiplierOut_394,MultiplierOut_393}), .cin (
                 GND0), .s ({AddOutputLvL1_95,AddOutputLvL1_94,AddOutputLvL1_93,
                 AddOutputLvL1_92,AddOutputLvL1_91,AddOutputLvL1_90,
                 AddOutputLvL1_89,AddOutputLvL1_88,AddOutputLvL1_87,
                 AddOutputLvL1_86,AddOutputLvL1_85,AddOutputLvL1_84,
                 AddOutputLvL1_83,AddOutputLvL1_82,AddOutputLvL1_81,
                 AddOutputLvL1_80}), .cout (\$dummy [409])) ;
    my_nadder_16 adder7 (.a ({MultiplierOut_440,MultiplierOut_439,
                 MultiplierOut_438,MultiplierOut_437,MultiplierOut_436,
                 MultiplierOut_435,MultiplierOut_434,MultiplierOut_433,
                 MultiplierOut_432,MultiplierOut_431,MultiplierOut_430,
                 MultiplierOut_429,MultiplierOut_428,MultiplierOut_427,
                 MultiplierOut_426,MultiplierOut_425}), .b ({MultiplierOut_472,
                 MultiplierOut_471,MultiplierOut_470,MultiplierOut_469,
                 MultiplierOut_468,MultiplierOut_467,MultiplierOut_466,
                 MultiplierOut_465,MultiplierOut_464,MultiplierOut_463,
                 MultiplierOut_462,MultiplierOut_461,MultiplierOut_460,
                 MultiplierOut_459,MultiplierOut_458,MultiplierOut_457}), .cin (
                 GND0), .s ({AddOutputLvL1_111,AddOutputLvL1_110,
                 AddOutputLvL1_109,AddOutputLvL1_108,AddOutputLvL1_107,
                 AddOutputLvL1_106,AddOutputLvL1_105,AddOutputLvL1_104,
                 AddOutputLvL1_103,AddOutputLvL1_102,AddOutputLvL1_101,
                 AddOutputLvL1_100,AddOutputLvL1_99,AddOutputLvL1_98,
                 AddOutputLvL1_97,AddOutputLvL1_96}), .cout (\$dummy [410])) ;
    my_nadder_16 adder8 (.a ({MultiplierOut_504,MultiplierOut_503,
                 MultiplierOut_502,MultiplierOut_501,MultiplierOut_500,
                 MultiplierOut_499,MultiplierOut_498,MultiplierOut_497,
                 MultiplierOut_496,MultiplierOut_495,MultiplierOut_494,
                 MultiplierOut_493,MultiplierOut_492,MultiplierOut_491,
                 MultiplierOut_490,MultiplierOut_489}), .b ({MultiplierOut_536,
                 MultiplierOut_535,MultiplierOut_534,MultiplierOut_533,
                 MultiplierOut_532,MultiplierOut_531,MultiplierOut_530,
                 MultiplierOut_529,MultiplierOut_528,MultiplierOut_527,
                 MultiplierOut_526,MultiplierOut_525,MultiplierOut_524,
                 MultiplierOut_523,MultiplierOut_522,MultiplierOut_521}), .cin (
                 GND0), .s ({AddOutputLvL1_127,AddOutputLvL1_126,
                 AddOutputLvL1_125,AddOutputLvL1_124,AddOutputLvL1_123,
                 AddOutputLvL1_122,AddOutputLvL1_121,AddOutputLvL1_120,
                 AddOutputLvL1_119,AddOutputLvL1_118,AddOutputLvL1_117,
                 AddOutputLvL1_116,AddOutputLvL1_115,AddOutputLvL1_114,
                 AddOutputLvL1_113,AddOutputLvL1_112}), .cout (\$dummy [411])) ;
    my_nadder_16 adder9 (.a ({MultiplierOut_568,MultiplierOut_567,
                 MultiplierOut_566,MultiplierOut_565,MultiplierOut_564,
                 MultiplierOut_563,MultiplierOut_562,MultiplierOut_561,
                 MultiplierOut_560,MultiplierOut_559,MultiplierOut_558,
                 MultiplierOut_557,MultiplierOut_556,MultiplierOut_555,
                 MultiplierOut_554,MultiplierOut_553}), .b ({MultiplierOut_600,
                 MultiplierOut_599,MultiplierOut_598,MultiplierOut_597,
                 MultiplierOut_596,MultiplierOut_595,MultiplierOut_594,
                 MultiplierOut_593,MultiplierOut_592,MultiplierOut_591,
                 MultiplierOut_590,MultiplierOut_589,MultiplierOut_588,
                 MultiplierOut_587,MultiplierOut_586,MultiplierOut_585}), .cin (
                 GND0), .s ({AddOutputLvL1_143,AddOutputLvL1_142,
                 AddOutputLvL1_141,AddOutputLvL1_140,AddOutputLvL1_139,
                 AddOutputLvL1_138,AddOutputLvL1_137,AddOutputLvL1_136,
                 AddOutputLvL1_135,AddOutputLvL1_134,AddOutputLvL1_133,
                 AddOutputLvL1_132,AddOutputLvL1_131,AddOutputLvL1_130,
                 AddOutputLvL1_129,AddOutputLvL1_128}), .cout (\$dummy [412])) ;
    my_nadder_16 adder10 (.a ({MultiplierOut_632,MultiplierOut_631,
                 MultiplierOut_630,MultiplierOut_629,MultiplierOut_628,
                 MultiplierOut_627,MultiplierOut_626,MultiplierOut_625,
                 MultiplierOut_624,MultiplierOut_623,MultiplierOut_622,
                 MultiplierOut_621,MultiplierOut_620,MultiplierOut_619,
                 MultiplierOut_618,MultiplierOut_617}), .b ({MultiplierOut_664,
                 MultiplierOut_663,MultiplierOut_662,MultiplierOut_661,
                 MultiplierOut_660,MultiplierOut_659,MultiplierOut_658,
                 MultiplierOut_657,MultiplierOut_656,MultiplierOut_655,
                 MultiplierOut_654,MultiplierOut_653,MultiplierOut_652,
                 MultiplierOut_651,MultiplierOut_650,MultiplierOut_649}), .cin (
                 GND0), .s ({AddOutputLvL1_159,AddOutputLvL1_158,
                 AddOutputLvL1_157,AddOutputLvL1_156,AddOutputLvL1_155,
                 AddOutputLvL1_154,AddOutputLvL1_153,AddOutputLvL1_152,
                 AddOutputLvL1_151,AddOutputLvL1_150,AddOutputLvL1_149,
                 AddOutputLvL1_148,AddOutputLvL1_147,AddOutputLvL1_146,
                 AddOutputLvL1_145,AddOutputLvL1_144}), .cout (\$dummy [413])) ;
    my_nadder_16 adder11 (.a ({MultiplierOut_696,MultiplierOut_695,
                 MultiplierOut_694,MultiplierOut_693,MultiplierOut_692,
                 MultiplierOut_691,MultiplierOut_690,MultiplierOut_689,
                 MultiplierOut_688,MultiplierOut_687,MultiplierOut_686,
                 MultiplierOut_685,MultiplierOut_684,MultiplierOut_683,
                 MultiplierOut_682,MultiplierOut_681}), .b ({MultiplierOut_728,
                 MultiplierOut_727,MultiplierOut_726,MultiplierOut_725,
                 MultiplierOut_724,MultiplierOut_723,MultiplierOut_722,
                 MultiplierOut_721,MultiplierOut_720,MultiplierOut_719,
                 MultiplierOut_718,MultiplierOut_717,MultiplierOut_716,
                 MultiplierOut_715,MultiplierOut_714,MultiplierOut_713}), .cin (
                 GND0), .s ({AddOutputLvL1_175,AddOutputLvL1_174,
                 AddOutputLvL1_173,AddOutputLvL1_172,AddOutputLvL1_171,
                 AddOutputLvL1_170,AddOutputLvL1_169,AddOutputLvL1_168,
                 AddOutputLvL1_167,AddOutputLvL1_166,AddOutputLvL1_165,
                 AddOutputLvL1_164,AddOutputLvL1_163,AddOutputLvL1_162,
                 AddOutputLvL1_161,AddOutputLvL1_160}), .cout (\$dummy [414])) ;
    my_nadder_16 adder0 (.a ({MultiplierOut_760,MultiplierOut_759,
                 MultiplierOut_758,MultiplierOut_757,MultiplierOut_756,
                 MultiplierOut_755,MultiplierOut_754,MultiplierOut_753,
                 MultiplierOut_752,MultiplierOut_751,MultiplierOut_750,
                 MultiplierOut_749,MultiplierOut_748,MultiplierOut_747,
                 MultiplierOut_746,MultiplierOut_745}), .b ({MultiplierOut_792,
                 MultiplierOut_791,MultiplierOut_790,MultiplierOut_789,
                 MultiplierOut_788,MultiplierOut_787,MultiplierOut_786,
                 MultiplierOut_785,MultiplierOut_784,MultiplierOut_783,
                 MultiplierOut_782,MultiplierOut_781,MultiplierOut_780,
                 MultiplierOut_779,MultiplierOut_778,MultiplierOut_777}), .cin (
                 GND0), .s ({AddOutputLvL1_191,AddOutputLvL1_190,
                 AddOutputLvL1_189,AddOutputLvL1_188,AddOutputLvL1_187,
                 AddOutputLvL1_186,AddOutputLvL1_185,AddOutputLvL1_184,
                 AddOutputLvL1_183,AddOutputLvL1_182,AddOutputLvL1_181,
                 AddOutputLvL1_180,AddOutputLvL1_179,AddOutputLvL1_178,
                 AddOutputLvL1_177,AddOutputLvL1_176}), .cout (\$dummy [415])) ;
    my_nadder_16 adder14 (.a ({AddOutputLvL1_79,AddOutputLvL1_78,
                 AddOutputLvL1_77,AddOutputLvL1_76,AddOutputLvL1_75,
                 AddOutputLvL1_74,AddOutputLvL1_73,AddOutputLvL1_72,
                 AddOutputLvL1_71,AddOutputLvL1_70,AddOutputLvL1_69,
                 AddOutputLvL1_68,AddOutputLvL1_67,AddOutputLvL1_66,
                 AddOutputLvL1_65,AddOutputLvL1_64}), .b ({AddOutputLvL1_95,
                 AddOutputLvL1_94,AddOutputLvL1_93,AddOutputLvL1_92,
                 AddOutputLvL1_91,AddOutputLvL1_90,AddOutputLvL1_89,
                 AddOutputLvL1_88,AddOutputLvL1_87,AddOutputLvL1_86,
                 AddOutputLvL1_85,AddOutputLvL1_84,AddOutputLvL1_83,
                 AddOutputLvL1_82,AddOutputLvL1_81,AddOutputLvL1_80}), .cin (
                 GND0), .s ({AddOutputLvL2_47,AddOutputLvL2_46,AddOutputLvL2_45,
                 AddOutputLvL2_44,AddOutputLvL2_43,AddOutputLvL2_42,
                 AddOutputLvL2_41,AddOutputLvL2_40,AddOutputLvL2_39,
                 AddOutputLvL2_38,AddOutputLvL2_37,AddOutputLvL2_36,
                 AddOutputLvL2_35,AddOutputLvL2_34,AddOutputLvL2_33,
                 AddOutputLvL2_32}), .cout (\$dummy [416])) ;
    my_nadder_16 adder15 (.a ({AddOutputLvL1_111,AddOutputLvL1_110,
                 AddOutputLvL1_109,AddOutputLvL1_108,AddOutputLvL1_107,
                 AddOutputLvL1_106,AddOutputLvL1_105,AddOutputLvL1_104,
                 AddOutputLvL1_103,AddOutputLvL1_102,AddOutputLvL1_101,
                 AddOutputLvL1_100,AddOutputLvL1_99,AddOutputLvL1_98,
                 AddOutputLvL1_97,AddOutputLvL1_96}), .b ({AddOutputLvL1_127,
                 AddOutputLvL1_126,AddOutputLvL1_125,AddOutputLvL1_124,
                 AddOutputLvL1_123,AddOutputLvL1_122,AddOutputLvL1_121,
                 AddOutputLvL1_120,AddOutputLvL1_119,AddOutputLvL1_118,
                 AddOutputLvL1_117,AddOutputLvL1_116,AddOutputLvL1_115,
                 AddOutputLvL1_114,AddOutputLvL1_113,AddOutputLvL1_112}), .cin (
                 GND0), .s ({AddOutputLvL2_63,AddOutputLvL2_62,AddOutputLvL2_61,
                 AddOutputLvL2_60,AddOutputLvL2_59,AddOutputLvL2_58,
                 AddOutputLvL2_57,AddOutputLvL2_56,AddOutputLvL2_55,
                 AddOutputLvL2_54,AddOutputLvL2_53,AddOutputLvL2_52,
                 AddOutputLvL2_51,AddOutputLvL2_50,AddOutputLvL2_49,
                 AddOutputLvL2_48}), .cout (\$dummy [417])) ;
    my_nadder_16 adder16 (.a ({AddOutputLvL1_143,AddOutputLvL1_142,
                 AddOutputLvL1_141,AddOutputLvL1_140,AddOutputLvL1_139,
                 AddOutputLvL1_138,AddOutputLvL1_137,AddOutputLvL1_136,
                 AddOutputLvL1_135,AddOutputLvL1_134,AddOutputLvL1_133,
                 AddOutputLvL1_132,AddOutputLvL1_131,AddOutputLvL1_130,
                 AddOutputLvL1_129,AddOutputLvL1_128}), .b ({AddOutputLvL1_159,
                 AddOutputLvL1_158,AddOutputLvL1_157,AddOutputLvL1_156,
                 AddOutputLvL1_155,AddOutputLvL1_154,AddOutputLvL1_153,
                 AddOutputLvL1_152,AddOutputLvL1_151,AddOutputLvL1_150,
                 AddOutputLvL1_149,AddOutputLvL1_148,AddOutputLvL1_147,
                 AddOutputLvL1_146,AddOutputLvL1_145,AddOutputLvL1_144}), .cin (
                 GND0), .s ({AddOutputLvL2_79,AddOutputLvL2_78,AddOutputLvL2_77,
                 AddOutputLvL2_76,AddOutputLvL2_75,AddOutputLvL2_74,
                 AddOutputLvL2_73,AddOutputLvL2_72,AddOutputLvL2_71,
                 AddOutputLvL2_70,AddOutputLvL2_69,AddOutputLvL2_68,
                 AddOutputLvL2_67,AddOutputLvL2_66,AddOutputLvL2_65,
                 AddOutputLvL2_64}), .cout (\$dummy [418])) ;
    my_nadder_16 adder17 (.a ({AddOutputLvL1_175,AddOutputLvL1_174,
                 AddOutputLvL1_173,AddOutputLvL1_172,AddOutputLvL1_171,
                 AddOutputLvL1_170,AddOutputLvL1_169,AddOutputLvL1_168,
                 AddOutputLvL1_167,AddOutputLvL1_166,AddOutputLvL1_165,
                 AddOutputLvL1_164,AddOutputLvL1_163,AddOutputLvL1_162,
                 AddOutputLvL1_161,AddOutputLvL1_160}), .b ({AddOutputLvL1_191,
                 AddOutputLvL1_190,AddOutputLvL1_189,AddOutputLvL1_188,
                 AddOutputLvL1_187,AddOutputLvL1_186,AddOutputLvL1_185,
                 AddOutputLvL1_184,AddOutputLvL1_183,AddOutputLvL1_182,
                 AddOutputLvL1_181,AddOutputLvL1_180,AddOutputLvL1_179,
                 AddOutputLvL1_178,AddOutputLvL1_177,AddOutputLvL1_176}), .cin (
                 GND0), .s ({AddOutputLvL2_95,AddOutputLvL2_94,AddOutputLvL2_93,
                 AddOutputLvL2_92,AddOutputLvL2_91,AddOutputLvL2_90,
                 AddOutputLvL2_89,AddOutputLvL2_88,AddOutputLvL2_87,
                 AddOutputLvL2_86,AddOutputLvL2_85,AddOutputLvL2_84,
                 AddOutputLvL2_83,AddOutputLvL2_82,AddOutputLvL2_81,
                 AddOutputLvL2_80}), .cout (\$dummy [419])) ;
    my_nadder_16 adder19 (.a ({AddOutputLvL2_47,AddOutputLvL2_46,
                 AddOutputLvL2_45,AddOutputLvL2_44,AddOutputLvL2_43,
                 AddOutputLvL2_42,AddOutputLvL2_41,AddOutputLvL2_40,
                 AddOutputLvL2_39,AddOutputLvL2_38,AddOutputLvL2_37,
                 AddOutputLvL2_36,AddOutputLvL2_35,AddOutputLvL2_34,
                 AddOutputLvL2_33,AddOutputLvL2_32}), .b ({AddOutputLvL2_63,
                 AddOutputLvL2_62,AddOutputLvL2_61,AddOutputLvL2_60,
                 AddOutputLvL2_59,AddOutputLvL2_58,AddOutputLvL2_57,
                 AddOutputLvL2_56,AddOutputLvL2_55,AddOutputLvL2_54,
                 AddOutputLvL2_53,AddOutputLvL2_52,AddOutputLvL2_51,
                 AddOutputLvL2_50,AddOutputLvL2_49,AddOutputLvL2_48}), .cin (
                 GND0), .s ({AddOutputLvL3_31,AddOutputLvL3_30,AddOutputLvL3_29,
                 AddOutputLvL3_28,AddOutputLvL3_27,AddOutputLvL3_26,
                 AddOutputLvL3_25,AddOutputLvL3_24,AddOutputLvL3_23,
                 AddOutputLvL3_22,AddOutputLvL3_21,AddOutputLvL3_20,
                 AddOutputLvL3_19,AddOutputLvL3_18,AddOutputLvL3_17,
                 AddOutputLvL3_16}), .cout (\$dummy [420])) ;
    my_nadder_16 adder20 (.a ({AddOutputLvL2_79,AddOutputLvL2_78,
                 AddOutputLvL2_77,AddOutputLvL2_76,AddOutputLvL2_75,
                 AddOutputLvL2_74,AddOutputLvL2_73,AddOutputLvL2_72,
                 AddOutputLvL2_71,AddOutputLvL2_70,AddOutputLvL2_69,
                 AddOutputLvL2_68,AddOutputLvL2_67,AddOutputLvL2_66,
                 AddOutputLvL2_65,AddOutputLvL2_64}), .b ({AddOutputLvL2_95,
                 AddOutputLvL2_94,AddOutputLvL2_93,AddOutputLvL2_92,
                 AddOutputLvL2_91,AddOutputLvL2_90,AddOutputLvL2_89,
                 AddOutputLvL2_88,AddOutputLvL2_87,AddOutputLvL2_86,
                 AddOutputLvL2_85,AddOutputLvL2_84,AddOutputLvL2_83,
                 AddOutputLvL2_82,AddOutputLvL2_81,AddOutputLvL2_80}), .cin (
                 GND0), .s ({AddOutputLvL3_47,AddOutputLvL3_46,AddOutputLvL3_45,
                 AddOutputLvL3_44,AddOutputLvL3_43,AddOutputLvL3_42,
                 AddOutputLvL3_41,AddOutputLvL3_40,AddOutputLvL3_39,
                 AddOutputLvL3_38,AddOutputLvL3_37,AddOutputLvL3_36,
                 AddOutputLvL3_35,AddOutputLvL3_34,AddOutputLvL3_33,
                 AddOutputLvL3_32}), .cout (\$dummy [421])) ;
    my_nadder_16 adder22 (.a ({AddOutputLvL3_31,AddOutputLvL3_30,
                 AddOutputLvL3_29,AddOutputLvL3_28,AddOutputLvL3_27,
                 AddOutputLvL3_26,AddOutputLvL3_25,AddOutputLvL3_24,
                 AddOutputLvL3_23,AddOutputLvL3_22,AddOutputLvL3_21,
                 AddOutputLvL3_20,AddOutputLvL3_19,AddOutputLvL3_18,
                 AddOutputLvL3_17,AddOutputLvL3_16}), .b ({AddOutputLvL3_47,
                 AddOutputLvL3_46,AddOutputLvL3_45,AddOutputLvL3_44,
                 AddOutputLvL3_43,AddOutputLvL3_42,AddOutputLvL3_41,
                 AddOutputLvL3_40,AddOutputLvL3_39,AddOutputLvL3_38,
                 AddOutputLvL3_37,AddOutputLvL3_36,AddOutputLvL3_35,
                 AddOutputLvL3_34,AddOutputLvL3_33,AddOutputLvL3_32}), .cin (
                 GND0), .s ({AddOut55_15,AddOut55_14,AddOut55_13,AddOut55_12,
                 AddOut55_11,AddOut55_10,AddOut55_9,AddOut55_8,AddOut55_7,
                 AddOut55_6,AddOut55_5,AddOut55_4,AddOut55_3,AddOut55_2,
                 AddOut55_1,AddOut55_0}), .cout (\$dummy [422])) ;
    my_nadder_16 adder23 (.a ({AddOut55_15,AddOut55_14,AddOut55_13,AddOut55_12,
                 AddOut55_11,AddOut55_10,AddOut55_9,AddOut55_8,AddOut55_7,
                 AddOut55_6,AddOut55_5,AddOut55_4,AddOut55_3,AddOut55_2,
                 AddOut55_1,AddOut55_0}), .b ({AddOut33_15,AddOut33_14,
                 AddOut33_13,AddOut33_12,AddOut33_11,AddOut33_10,AddOut33_9,
                 AddOut33_8,AddOut33_7,AddOut33_6,AddOut33_5,AddOut33_4,
                 AddOut33_3,AddOut33_2,AddOut33_1,AddOut33_0}), .cin (GND0), .s (
                 {Final55_15,Final55_14,Final55_13,Final55_12,Final55_11,
                 Final55_10,Final55_9,Final55_8,Final55_7,Final55_6,Final55_5,
                 Final55_4,Final55_3,Final55_2,Final55_1,Final55_0}), .cout (
                 \$dummy [423])) ;
    Counter_3 EndCounter (.enable (CountereEN), .reset (CountereRST), .clk (CLK)
              , .load (GND0), .\output  ({CounterOut_2,CounterOut_1,CounterOut_0
              }), .\input  ({GND0,GND0,GND0})) ;
    fake_gnd ix6941 (.Y (GND0)) ;
    or02 ix3555 (.Y (CountereRST), .A0 (nx3552), .A1 (RST)) ;
    nor03_2x ix3553 (.Y (nx3552), .A0 (CounterOut_0), .A1 (nx7936), .A2 (
             CounterOut_1)) ;
    inv01 ix7937 (.Y (nx7936), .A (CounterOut_2)) ;
    nor02ii ix3571 (.Y (CountereEN), .A0 (ACK), .A1 (current_state[7])) ;
    dffs_ni reg_ACKC_dup_1 (.Q (ACK), .QB (\$dummy [424]), .D (GND0), .CLK (CLK)
            , .S (nx3562)) ;
    and03 ix3563 (.Y (nx3562), .A0 (CounterOut_0), .A1 (nx7936), .A2 (
          CounterOut_1)) ;
    mux21_ni ix3425 (.Y (SecondInputToMult_48), .A0 (OutputImg1[0]), .A1 (
             OutputImg0[48]), .S0 (nx8858)) ;
    mux21_ni ix3433 (.Y (SecondInputToMult_49), .A0 (OutputImg1[1]), .A1 (
             OutputImg0[49]), .S0 (nx8858)) ;
    mux21_ni ix3441 (.Y (SecondInputToMult_50), .A0 (OutputImg1[2]), .A1 (
             OutputImg0[50]), .S0 (nx8858)) ;
    mux21_ni ix3449 (.Y (SecondInputToMult_51), .A0 (OutputImg1[3]), .A1 (
             OutputImg0[51]), .S0 (nx8858)) ;
    mux21_ni ix3457 (.Y (SecondInputToMult_52), .A0 (OutputImg1[4]), .A1 (
             OutputImg0[52]), .S0 (nx8858)) ;
    mux21_ni ix3465 (.Y (SecondInputToMult_53), .A0 (OutputImg1[5]), .A1 (
             OutputImg0[53]), .S0 (nx8858)) ;
    mux21_ni ix3473 (.Y (SecondInputToMult_54), .A0 (OutputImg1[6]), .A1 (
             OutputImg0[54]), .S0 (nx8858)) ;
    mux21_ni ix3481 (.Y (SecondInputToMult_55), .A0 (OutputImg1[7]), .A1 (
             OutputImg0[55]), .S0 (nx8860)) ;
    mux21_ni ix3489 (.Y (SecondInputToMult_56), .A0 (OutputImg1[8]), .A1 (
             OutputImg0[56]), .S0 (nx8860)) ;
    mux21_ni ix3497 (.Y (SecondInputToMult_57), .A0 (OutputImg1[9]), .A1 (
             OutputImg0[57]), .S0 (nx8860)) ;
    mux21_ni ix3505 (.Y (SecondInputToMult_58), .A0 (OutputImg1[10]), .A1 (
             OutputImg0[58]), .S0 (nx8860)) ;
    mux21_ni ix3513 (.Y (SecondInputToMult_59), .A0 (OutputImg1[11]), .A1 (
             OutputImg0[59]), .S0 (nx8860)) ;
    mux21_ni ix3521 (.Y (SecondInputToMult_60), .A0 (OutputImg1[12]), .A1 (
             OutputImg0[60]), .S0 (nx8860)) ;
    mux21_ni ix3529 (.Y (SecondInputToMult_61), .A0 (OutputImg1[13]), .A1 (
             OutputImg0[61]), .S0 (nx8860)) ;
    mux21_ni ix3537 (.Y (SecondInputToMult_62), .A0 (OutputImg1[14]), .A1 (
             OutputImg0[62]), .S0 (nx8862)) ;
    mux21_ni ix3545 (.Y (SecondInputToMult_63), .A0 (OutputImg1[15]), .A1 (
             OutputImg0[63]), .S0 (nx8862)) ;
    mux21_ni ix3297 (.Y (SecondInputToMult_64), .A0 (OutputImg1[16]), .A1 (
             OutputImg0[64]), .S0 (nx8862)) ;
    mux21_ni ix3305 (.Y (SecondInputToMult_65), .A0 (OutputImg1[17]), .A1 (
             OutputImg0[65]), .S0 (nx8862)) ;
    mux21_ni ix3313 (.Y (SecondInputToMult_66), .A0 (OutputImg1[18]), .A1 (
             OutputImg0[66]), .S0 (nx8862)) ;
    mux21_ni ix3321 (.Y (SecondInputToMult_67), .A0 (OutputImg1[19]), .A1 (
             OutputImg0[67]), .S0 (nx8862)) ;
    mux21_ni ix3329 (.Y (SecondInputToMult_68), .A0 (OutputImg1[20]), .A1 (
             OutputImg0[68]), .S0 (nx8862)) ;
    mux21_ni ix3337 (.Y (SecondInputToMult_69), .A0 (OutputImg1[21]), .A1 (
             OutputImg0[69]), .S0 (nx8864)) ;
    mux21_ni ix3345 (.Y (SecondInputToMult_70), .A0 (OutputImg1[22]), .A1 (
             OutputImg0[70]), .S0 (nx8864)) ;
    mux21_ni ix3353 (.Y (SecondInputToMult_71), .A0 (OutputImg1[23]), .A1 (
             OutputImg0[71]), .S0 (nx8864)) ;
    mux21_ni ix3361 (.Y (SecondInputToMult_72), .A0 (OutputImg1[24]), .A1 (
             OutputImg0[72]), .S0 (nx8864)) ;
    mux21_ni ix3369 (.Y (SecondInputToMult_73), .A0 (OutputImg1[25]), .A1 (
             OutputImg0[73]), .S0 (nx8864)) ;
    mux21_ni ix3377 (.Y (SecondInputToMult_74), .A0 (OutputImg1[26]), .A1 (
             OutputImg0[74]), .S0 (nx8864)) ;
    mux21_ni ix3385 (.Y (SecondInputToMult_75), .A0 (OutputImg1[27]), .A1 (
             OutputImg0[75]), .S0 (nx8864)) ;
    mux21_ni ix3393 (.Y (SecondInputToMult_76), .A0 (OutputImg1[28]), .A1 (
             OutputImg0[76]), .S0 (nx8866)) ;
    mux21_ni ix3401 (.Y (SecondInputToMult_77), .A0 (OutputImg1[29]), .A1 (
             OutputImg0[77]), .S0 (nx8866)) ;
    mux21_ni ix3409 (.Y (SecondInputToMult_78), .A0 (OutputImg1[30]), .A1 (
             OutputImg0[78]), .S0 (nx8866)) ;
    mux21_ni ix3417 (.Y (SecondInputToMult_79), .A0 (OutputImg1[31]), .A1 (
             OutputImg0[79]), .S0 (nx8866)) ;
    mux21_ni ix3169 (.Y (SecondInputToMult_80), .A0 (OutputImg1[32]), .A1 (
             OutputImg1[0]), .S0 (nx8866)) ;
    mux21_ni ix3177 (.Y (SecondInputToMult_81), .A0 (OutputImg1[33]), .A1 (
             OutputImg1[1]), .S0 (nx8866)) ;
    mux21_ni ix3185 (.Y (SecondInputToMult_82), .A0 (OutputImg1[34]), .A1 (
             OutputImg1[2]), .S0 (nx8866)) ;
    mux21_ni ix3193 (.Y (SecondInputToMult_83), .A0 (OutputImg1[35]), .A1 (
             OutputImg1[3]), .S0 (nx8868)) ;
    mux21_ni ix3201 (.Y (SecondInputToMult_84), .A0 (OutputImg1[36]), .A1 (
             OutputImg1[4]), .S0 (nx8868)) ;
    mux21_ni ix3209 (.Y (SecondInputToMult_85), .A0 (OutputImg1[37]), .A1 (
             OutputImg1[5]), .S0 (nx8868)) ;
    mux21_ni ix3217 (.Y (SecondInputToMult_86), .A0 (OutputImg1[38]), .A1 (
             OutputImg1[6]), .S0 (nx8868)) ;
    mux21_ni ix3225 (.Y (SecondInputToMult_87), .A0 (OutputImg1[39]), .A1 (
             OutputImg1[7]), .S0 (nx8868)) ;
    mux21_ni ix3233 (.Y (SecondInputToMult_88), .A0 (OutputImg1[40]), .A1 (
             OutputImg1[8]), .S0 (nx8868)) ;
    mux21_ni ix3241 (.Y (SecondInputToMult_89), .A0 (OutputImg1[41]), .A1 (
             OutputImg1[9]), .S0 (nx8868)) ;
    mux21_ni ix3249 (.Y (SecondInputToMult_90), .A0 (OutputImg1[42]), .A1 (
             OutputImg1[10]), .S0 (nx8870)) ;
    mux21_ni ix3257 (.Y (SecondInputToMult_91), .A0 (OutputImg1[43]), .A1 (
             OutputImg1[11]), .S0 (nx8870)) ;
    mux21_ni ix3265 (.Y (SecondInputToMult_92), .A0 (OutputImg1[44]), .A1 (
             OutputImg1[12]), .S0 (nx8870)) ;
    mux21_ni ix3273 (.Y (SecondInputToMult_93), .A0 (OutputImg1[45]), .A1 (
             OutputImg1[13]), .S0 (nx8870)) ;
    mux21_ni ix3281 (.Y (SecondInputToMult_94), .A0 (OutputImg1[46]), .A1 (
             OutputImg1[14]), .S0 (nx8870)) ;
    mux21_ni ix3289 (.Y (SecondInputToMult_95), .A0 (OutputImg1[47]), .A1 (
             OutputImg1[15]), .S0 (nx8870)) ;
    mux21_ni ix3041 (.Y (SecondInputToMult_96), .A0 (OutputImg2[0]), .A1 (
             OutputImg1[16]), .S0 (nx8870)) ;
    mux21_ni ix3049 (.Y (SecondInputToMult_97), .A0 (OutputImg2[1]), .A1 (
             OutputImg1[17]), .S0 (nx8872)) ;
    mux21_ni ix3057 (.Y (SecondInputToMult_98), .A0 (OutputImg2[2]), .A1 (
             OutputImg1[18]), .S0 (nx8872)) ;
    mux21_ni ix3065 (.Y (SecondInputToMult_99), .A0 (OutputImg2[3]), .A1 (
             OutputImg1[19]), .S0 (nx8872)) ;
    mux21_ni ix3073 (.Y (SecondInputToMult_100), .A0 (OutputImg2[4]), .A1 (
             OutputImg1[20]), .S0 (nx8872)) ;
    mux21_ni ix3081 (.Y (SecondInputToMult_101), .A0 (OutputImg2[5]), .A1 (
             OutputImg1[21]), .S0 (nx8872)) ;
    mux21_ni ix3089 (.Y (SecondInputToMult_102), .A0 (OutputImg2[6]), .A1 (
             OutputImg1[22]), .S0 (nx8872)) ;
    mux21_ni ix3097 (.Y (SecondInputToMult_103), .A0 (OutputImg2[7]), .A1 (
             OutputImg1[23]), .S0 (nx8872)) ;
    mux21_ni ix3105 (.Y (SecondInputToMult_104), .A0 (OutputImg2[8]), .A1 (
             OutputImg1[24]), .S0 (nx8874)) ;
    mux21_ni ix3113 (.Y (SecondInputToMult_105), .A0 (OutputImg2[9]), .A1 (
             OutputImg1[25]), .S0 (nx8874)) ;
    mux21_ni ix3121 (.Y (SecondInputToMult_106), .A0 (OutputImg2[10]), .A1 (
             OutputImg1[26]), .S0 (nx8874)) ;
    mux21_ni ix3129 (.Y (SecondInputToMult_107), .A0 (OutputImg2[11]), .A1 (
             OutputImg1[27]), .S0 (nx8874)) ;
    mux21_ni ix3137 (.Y (SecondInputToMult_108), .A0 (OutputImg2[12]), .A1 (
             OutputImg1[28]), .S0 (nx8874)) ;
    mux21_ni ix3145 (.Y (SecondInputToMult_109), .A0 (OutputImg2[13]), .A1 (
             OutputImg1[29]), .S0 (nx8874)) ;
    mux21_ni ix3153 (.Y (SecondInputToMult_110), .A0 (OutputImg2[14]), .A1 (
             OutputImg1[30]), .S0 (nx8874)) ;
    mux21_ni ix3161 (.Y (SecondInputToMult_111), .A0 (OutputImg2[15]), .A1 (
             OutputImg1[31]), .S0 (nx8876)) ;
    mux21_ni ix2913 (.Y (SecondInputToMult_112), .A0 (OutputImg2[16]), .A1 (
             OutputImg1[32]), .S0 (nx8876)) ;
    mux21_ni ix2921 (.Y (SecondInputToMult_113), .A0 (OutputImg2[17]), .A1 (
             OutputImg1[33]), .S0 (nx8876)) ;
    mux21_ni ix2929 (.Y (SecondInputToMult_114), .A0 (OutputImg2[18]), .A1 (
             OutputImg1[34]), .S0 (nx8876)) ;
    mux21_ni ix2937 (.Y (SecondInputToMult_115), .A0 (OutputImg2[19]), .A1 (
             OutputImg1[35]), .S0 (nx8876)) ;
    mux21_ni ix2945 (.Y (SecondInputToMult_116), .A0 (OutputImg2[20]), .A1 (
             OutputImg1[36]), .S0 (nx8876)) ;
    mux21_ni ix2953 (.Y (SecondInputToMult_117), .A0 (OutputImg2[21]), .A1 (
             OutputImg1[37]), .S0 (nx8876)) ;
    mux21_ni ix2961 (.Y (SecondInputToMult_118), .A0 (OutputImg2[22]), .A1 (
             OutputImg1[38]), .S0 (nx8878)) ;
    mux21_ni ix2969 (.Y (SecondInputToMult_119), .A0 (OutputImg2[23]), .A1 (
             OutputImg1[39]), .S0 (nx8878)) ;
    mux21_ni ix2977 (.Y (SecondInputToMult_120), .A0 (OutputImg2[24]), .A1 (
             OutputImg1[40]), .S0 (nx8878)) ;
    mux21_ni ix2985 (.Y (SecondInputToMult_121), .A0 (OutputImg2[25]), .A1 (
             OutputImg1[41]), .S0 (nx8878)) ;
    mux21_ni ix2993 (.Y (SecondInputToMult_122), .A0 (OutputImg2[26]), .A1 (
             OutputImg1[42]), .S0 (nx8878)) ;
    mux21_ni ix3001 (.Y (SecondInputToMult_123), .A0 (OutputImg2[27]), .A1 (
             OutputImg1[43]), .S0 (nx8878)) ;
    mux21_ni ix3009 (.Y (SecondInputToMult_124), .A0 (OutputImg2[28]), .A1 (
             OutputImg1[44]), .S0 (nx8878)) ;
    mux21_ni ix3017 (.Y (SecondInputToMult_125), .A0 (OutputImg2[29]), .A1 (
             OutputImg1[45]), .S0 (nx8880)) ;
    mux21_ni ix3025 (.Y (SecondInputToMult_126), .A0 (OutputImg2[30]), .A1 (
             OutputImg1[46]), .S0 (nx8880)) ;
    mux21_ni ix3033 (.Y (SecondInputToMult_127), .A0 (OutputImg2[31]), .A1 (
             OutputImg1[47]), .S0 (nx8880)) ;
    mux21_ni ix2785 (.Y (SecondInputToMult_128), .A0 (OutputImg2[32]), .A1 (
             OutputImg1[48]), .S0 (nx8880)) ;
    mux21_ni ix2793 (.Y (SecondInputToMult_129), .A0 (OutputImg2[33]), .A1 (
             OutputImg1[49]), .S0 (nx8880)) ;
    mux21_ni ix2801 (.Y (SecondInputToMult_130), .A0 (OutputImg2[34]), .A1 (
             OutputImg1[50]), .S0 (nx8880)) ;
    mux21_ni ix2809 (.Y (SecondInputToMult_131), .A0 (OutputImg2[35]), .A1 (
             OutputImg1[51]), .S0 (nx8880)) ;
    mux21_ni ix2817 (.Y (SecondInputToMult_132), .A0 (OutputImg2[36]), .A1 (
             OutputImg1[52]), .S0 (nx8882)) ;
    mux21_ni ix2825 (.Y (SecondInputToMult_133), .A0 (OutputImg2[37]), .A1 (
             OutputImg1[53]), .S0 (nx8882)) ;
    mux21_ni ix2833 (.Y (SecondInputToMult_134), .A0 (OutputImg2[38]), .A1 (
             OutputImg1[54]), .S0 (nx8882)) ;
    mux21_ni ix2841 (.Y (SecondInputToMult_135), .A0 (OutputImg2[39]), .A1 (
             OutputImg1[55]), .S0 (nx8882)) ;
    mux21_ni ix2849 (.Y (SecondInputToMult_136), .A0 (OutputImg2[40]), .A1 (
             OutputImg1[56]), .S0 (nx8882)) ;
    mux21_ni ix2857 (.Y (SecondInputToMult_137), .A0 (OutputImg2[41]), .A1 (
             OutputImg1[57]), .S0 (nx8882)) ;
    mux21_ni ix2865 (.Y (SecondInputToMult_138), .A0 (OutputImg2[42]), .A1 (
             OutputImg1[58]), .S0 (nx8882)) ;
    mux21_ni ix2873 (.Y (SecondInputToMult_139), .A0 (OutputImg2[43]), .A1 (
             OutputImg1[59]), .S0 (nx8884)) ;
    mux21_ni ix2881 (.Y (SecondInputToMult_140), .A0 (OutputImg2[44]), .A1 (
             OutputImg1[60]), .S0 (nx8884)) ;
    mux21_ni ix2889 (.Y (SecondInputToMult_141), .A0 (OutputImg2[45]), .A1 (
             OutputImg1[61]), .S0 (nx8884)) ;
    mux21_ni ix2897 (.Y (SecondInputToMult_142), .A0 (OutputImg2[46]), .A1 (
             OutputImg1[62]), .S0 (nx8884)) ;
    mux21_ni ix2905 (.Y (SecondInputToMult_143), .A0 (OutputImg2[47]), .A1 (
             OutputImg1[63]), .S0 (nx8884)) ;
    ao22 ix2681 (.Y (FilterToAlu_0), .A0 (outFilter0[0]), .A1 (nx8586), .B0 (
         outFilter1[0]), .B1 (nx8696)) ;
    nor02_2x ix511 (.Y (nx510), .A0 (nx8896), .A1 (nx8852)) ;
    ao22 ix2687 (.Y (FilterToAlu_1), .A0 (outFilter0[1]), .A1 (nx8586), .B0 (
         outFilter1[1]), .B1 (nx8696)) ;
    ao22 ix2693 (.Y (FilterToAlu_2), .A0 (outFilter0[2]), .A1 (nx8586), .B0 (
         outFilter1[2]), .B1 (nx8696)) ;
    ao22 ix2699 (.Y (FilterToAlu_3), .A0 (outFilter0[3]), .A1 (nx8586), .B0 (
         outFilter1[3]), .B1 (nx8696)) ;
    ao22 ix2705 (.Y (FilterToAlu_4), .A0 (outFilter0[4]), .A1 (nx8586), .B0 (
         outFilter1[4]), .B1 (nx8696)) ;
    ao22 ix2711 (.Y (FilterToAlu_5), .A0 (outFilter0[5]), .A1 (nx8586), .B0 (
         outFilter1[5]), .B1 (nx8696)) ;
    ao22 ix2717 (.Y (FilterToAlu_6), .A0 (outFilter0[6]), .A1 (nx8586), .B0 (
         outFilter1[6]), .B1 (nx8696)) ;
    ao22 ix2723 (.Y (FilterToAlu_7), .A0 (outFilter0[7]), .A1 (nx8588), .B0 (
         outFilter1[7]), .B1 (nx8698)) ;
    ao22 ix2729 (.Y (FilterToAlu_8), .A0 (outFilter0[8]), .A1 (nx8588), .B0 (
         outFilter1[8]), .B1 (nx8698)) ;
    nand02 ix505 (.Y (FilterToAlu_9), .A0 (nx8052), .A1 (nx8924)) ;
    mux21 ix8053 (.Y (nx8052), .A0 (outFilter0[9]), .A1 (outFilter1[9]), .S0 (
          nx8896)) ;
    ao22 ix2735 (.Y (FilterToAlu_10), .A0 (outFilter0[10]), .A1 (nx8588), .B0 (
         outFilter1[10]), .B1 (nx8698)) ;
    ao22 ix2741 (.Y (FilterToAlu_11), .A0 (outFilter0[11]), .A1 (nx8588), .B0 (
         outFilter1[11]), .B1 (nx8698)) ;
    ao22 ix2747 (.Y (FilterToAlu_12), .A0 (outFilter0[12]), .A1 (nx8588), .B0 (
         outFilter1[12]), .B1 (nx8698)) ;
    ao22 ix2753 (.Y (FilterToAlu_13), .A0 (outFilter0[13]), .A1 (nx8588), .B0 (
         outFilter1[13]), .B1 (nx8698)) ;
    ao22 ix2759 (.Y (FilterToAlu_14), .A0 (outFilter0[14]), .A1 (nx8588), .B0 (
         outFilter1[14]), .B1 (nx8698)) ;
    ao22 ix2765 (.Y (FilterToAlu_15), .A0 (outFilter0[15]), .A1 (nx8590), .B0 (
         outFilter1[15]), .B1 (nx8700)) ;
    ao22 ix2591 (.Y (FilterToAlu_16), .A0 (outFilter0[16]), .A1 (nx8590), .B0 (
         outFilter1[16]), .B1 (nx8700)) ;
    ao22 ix2597 (.Y (FilterToAlu_17), .A0 (outFilter0[17]), .A1 (nx8590), .B0 (
         outFilter1[17]), .B1 (nx8700)) ;
    ao22 ix2603 (.Y (FilterToAlu_18), .A0 (outFilter0[18]), .A1 (nx8590), .B0 (
         outFilter1[18]), .B1 (nx8700)) ;
    ao22 ix2609 (.Y (FilterToAlu_19), .A0 (outFilter0[19]), .A1 (nx8590), .B0 (
         outFilter1[19]), .B1 (nx8700)) ;
    ao22 ix2615 (.Y (FilterToAlu_20), .A0 (outFilter0[20]), .A1 (nx8590), .B0 (
         outFilter1[20]), .B1 (nx8700)) ;
    ao22 ix2621 (.Y (FilterToAlu_21), .A0 (outFilter0[21]), .A1 (nx8590), .B0 (
         outFilter1[21]), .B1 (nx8700)) ;
    ao22 ix2627 (.Y (FilterToAlu_22), .A0 (outFilter0[22]), .A1 (nx8592), .B0 (
         outFilter1[22]), .B1 (nx8702)) ;
    ao22 ix2633 (.Y (FilterToAlu_23), .A0 (outFilter0[23]), .A1 (nx8592), .B0 (
         outFilter1[23]), .B1 (nx8702)) ;
    ao22 ix2639 (.Y (FilterToAlu_24), .A0 (outFilter0[24]), .A1 (nx8592), .B0 (
         outFilter1[24]), .B1 (nx8702)) ;
    nand02 ix495 (.Y (FilterToAlu_25), .A0 (nx8072), .A1 (nx8924)) ;
    mux21 ix8073 (.Y (nx8072), .A0 (outFilter0[25]), .A1 (outFilter1[25]), .S0 (
          nx8896)) ;
    ao22 ix2645 (.Y (FilterToAlu_26), .A0 (outFilter0[26]), .A1 (nx8592), .B0 (
         outFilter1[26]), .B1 (nx8702)) ;
    ao22 ix2651 (.Y (FilterToAlu_27), .A0 (outFilter0[27]), .A1 (nx8592), .B0 (
         outFilter1[27]), .B1 (nx8702)) ;
    ao22 ix2657 (.Y (FilterToAlu_28), .A0 (outFilter0[28]), .A1 (nx8592), .B0 (
         outFilter1[28]), .B1 (nx8702)) ;
    ao22 ix2663 (.Y (FilterToAlu_29), .A0 (outFilter0[29]), .A1 (nx8592), .B0 (
         outFilter1[29]), .B1 (nx8702)) ;
    ao22 ix2669 (.Y (FilterToAlu_30), .A0 (outFilter0[30]), .A1 (nx8594), .B0 (
         outFilter1[30]), .B1 (nx8704)) ;
    ao22 ix2675 (.Y (FilterToAlu_31), .A0 (outFilter0[31]), .A1 (nx8594), .B0 (
         outFilter1[31]), .B1 (nx8704)) ;
    ao22 ix2501 (.Y (FilterToAlu_32), .A0 (outFilter0[32]), .A1 (nx8594), .B0 (
         outFilter1[32]), .B1 (nx8704)) ;
    ao22 ix2507 (.Y (FilterToAlu_33), .A0 (outFilter0[33]), .A1 (nx8594), .B0 (
         outFilter1[33]), .B1 (nx8704)) ;
    ao22 ix2513 (.Y (FilterToAlu_34), .A0 (outFilter0[34]), .A1 (nx8594), .B0 (
         outFilter1[34]), .B1 (nx8704)) ;
    ao22 ix2519 (.Y (FilterToAlu_35), .A0 (outFilter0[35]), .A1 (nx8594), .B0 (
         outFilter1[35]), .B1 (nx8704)) ;
    ao22 ix2525 (.Y (FilterToAlu_36), .A0 (outFilter0[36]), .A1 (nx8594), .B0 (
         outFilter1[36]), .B1 (nx8704)) ;
    ao22 ix2531 (.Y (FilterToAlu_37), .A0 (outFilter0[37]), .A1 (nx8596), .B0 (
         outFilter1[37]), .B1 (nx8706)) ;
    ao22 ix2537 (.Y (FilterToAlu_38), .A0 (outFilter0[38]), .A1 (nx8596), .B0 (
         outFilter1[38]), .B1 (nx8706)) ;
    ao22 ix2543 (.Y (FilterToAlu_39), .A0 (outFilter0[39]), .A1 (nx8596), .B0 (
         outFilter1[39]), .B1 (nx8706)) ;
    ao22 ix2549 (.Y (FilterToAlu_40), .A0 (outFilter0[40]), .A1 (nx8596), .B0 (
         outFilter1[40]), .B1 (nx8706)) ;
    nand02 ix485 (.Y (FilterToAlu_41), .A0 (nx8090), .A1 (nx8924)) ;
    mux21 ix8091 (.Y (nx8090), .A0 (outFilter0[41]), .A1 (outFilter1[41]), .S0 (
          nx8896)) ;
    ao22 ix2555 (.Y (FilterToAlu_42), .A0 (outFilter0[42]), .A1 (nx8596), .B0 (
         outFilter1[42]), .B1 (nx8706)) ;
    ao22 ix2561 (.Y (FilterToAlu_43), .A0 (outFilter0[43]), .A1 (nx8596), .B0 (
         outFilter1[43]), .B1 (nx8706)) ;
    ao22 ix2567 (.Y (FilterToAlu_44), .A0 (outFilter0[44]), .A1 (nx8596), .B0 (
         outFilter1[44]), .B1 (nx8706)) ;
    ao22 ix2573 (.Y (FilterToAlu_45), .A0 (outFilter0[45]), .A1 (nx8598), .B0 (
         outFilter1[45]), .B1 (nx8708)) ;
    ao22 ix2579 (.Y (FilterToAlu_46), .A0 (outFilter0[46]), .A1 (nx8598), .B0 (
         outFilter1[46]), .B1 (nx8708)) ;
    ao22 ix2585 (.Y (FilterToAlu_47), .A0 (outFilter0[47]), .A1 (nx8598), .B0 (
         outFilter1[47]), .B1 (nx8708)) ;
    ao22 ix2411 (.Y (FilterToAlu_48), .A0 (outFilter0[48]), .A1 (nx8598), .B0 (
         outFilter1[48]), .B1 (nx8708)) ;
    ao22 ix2417 (.Y (FilterToAlu_49), .A0 (outFilter0[49]), .A1 (nx8598), .B0 (
         outFilter1[49]), .B1 (nx8708)) ;
    ao22 ix2423 (.Y (FilterToAlu_50), .A0 (outFilter0[50]), .A1 (nx8598), .B0 (
         outFilter1[50]), .B1 (nx8708)) ;
    ao22 ix2429 (.Y (FilterToAlu_51), .A0 (outFilter0[51]), .A1 (nx8598), .B0 (
         outFilter1[51]), .B1 (nx8708)) ;
    ao22 ix2435 (.Y (FilterToAlu_52), .A0 (outFilter0[52]), .A1 (nx8600), .B0 (
         outFilter1[52]), .B1 (nx8710)) ;
    ao22 ix2441 (.Y (FilterToAlu_53), .A0 (outFilter0[53]), .A1 (nx8600), .B0 (
         outFilter1[53]), .B1 (nx8710)) ;
    ao22 ix2447 (.Y (FilterToAlu_54), .A0 (outFilter0[54]), .A1 (nx8600), .B0 (
         outFilter1[54]), .B1 (nx8710)) ;
    ao22 ix2453 (.Y (FilterToAlu_55), .A0 (outFilter0[55]), .A1 (nx8600), .B0 (
         outFilter1[55]), .B1 (nx8710)) ;
    ao22 ix2459 (.Y (FilterToAlu_56), .A0 (outFilter0[56]), .A1 (nx8600), .B0 (
         outFilter1[56]), .B1 (nx8710)) ;
    nand02 ix475 (.Y (FilterToAlu_57), .A0 (nx8108), .A1 (nx8924)) ;
    mux21 ix8109 (.Y (nx8108), .A0 (outFilter0[57]), .A1 (outFilter1[57]), .S0 (
          nx8896)) ;
    ao22 ix2465 (.Y (FilterToAlu_58), .A0 (outFilter0[58]), .A1 (nx8600), .B0 (
         outFilter1[58]), .B1 (nx8710)) ;
    ao22 ix2471 (.Y (FilterToAlu_59), .A0 (outFilter0[59]), .A1 (nx8600), .B0 (
         outFilter1[59]), .B1 (nx8710)) ;
    ao22 ix2477 (.Y (FilterToAlu_60), .A0 (outFilter0[60]), .A1 (nx8602), .B0 (
         outFilter1[60]), .B1 (nx8712)) ;
    ao22 ix2483 (.Y (FilterToAlu_61), .A0 (outFilter0[61]), .A1 (nx8602), .B0 (
         outFilter1[61]), .B1 (nx8712)) ;
    ao22 ix2489 (.Y (FilterToAlu_62), .A0 (outFilter0[62]), .A1 (nx8602), .B0 (
         outFilter1[62]), .B1 (nx8712)) ;
    ao22 ix2495 (.Y (FilterToAlu_63), .A0 (outFilter0[63]), .A1 (nx8602), .B0 (
         outFilter1[63]), .B1 (nx8712)) ;
    ao22 ix2321 (.Y (FilterToAlu_64), .A0 (outFilter0[64]), .A1 (nx8602), .B0 (
         outFilter1[64]), .B1 (nx8712)) ;
    ao22 ix2327 (.Y (FilterToAlu_65), .A0 (outFilter0[65]), .A1 (nx8602), .B0 (
         outFilter1[65]), .B1 (nx8712)) ;
    ao22 ix2333 (.Y (FilterToAlu_66), .A0 (outFilter0[66]), .A1 (nx8602), .B0 (
         outFilter1[66]), .B1 (nx8712)) ;
    ao22 ix2339 (.Y (FilterToAlu_67), .A0 (outFilter0[67]), .A1 (nx8604), .B0 (
         outFilter1[67]), .B1 (nx8714)) ;
    ao22 ix2345 (.Y (FilterToAlu_68), .A0 (outFilter0[68]), .A1 (nx8604), .B0 (
         outFilter1[68]), .B1 (nx8714)) ;
    ao22 ix2351 (.Y (FilterToAlu_69), .A0 (outFilter0[69]), .A1 (nx8604), .B0 (
         outFilter1[69]), .B1 (nx8714)) ;
    ao22 ix2357 (.Y (FilterToAlu_70), .A0 (outFilter0[70]), .A1 (nx8604), .B0 (
         outFilter1[70]), .B1 (nx8714)) ;
    ao22 ix2363 (.Y (FilterToAlu_71), .A0 (outFilter0[71]), .A1 (nx8604), .B0 (
         outFilter1[71]), .B1 (nx8714)) ;
    ao22 ix2369 (.Y (FilterToAlu_72), .A0 (outFilter0[72]), .A1 (nx8604), .B0 (
         outFilter1[72]), .B1 (nx8714)) ;
    nand02 ix465 (.Y (FilterToAlu_73), .A0 (nx8126), .A1 (nx8924)) ;
    mux21 ix8127 (.Y (nx8126), .A0 (outFilter0[73]), .A1 (outFilter1[73]), .S0 (
          nx8896)) ;
    ao22 ix2375 (.Y (FilterToAlu_74), .A0 (outFilter0[74]), .A1 (nx8604), .B0 (
         outFilter1[74]), .B1 (nx8714)) ;
    ao22 ix2381 (.Y (FilterToAlu_75), .A0 (outFilter0[75]), .A1 (nx8606), .B0 (
         outFilter1[75]), .B1 (nx8716)) ;
    ao22 ix2387 (.Y (FilterToAlu_76), .A0 (outFilter0[76]), .A1 (nx8606), .B0 (
         outFilter1[76]), .B1 (nx8716)) ;
    ao22 ix2393 (.Y (FilterToAlu_77), .A0 (outFilter0[77]), .A1 (nx8606), .B0 (
         outFilter1[77]), .B1 (nx8716)) ;
    ao22 ix2399 (.Y (FilterToAlu_78), .A0 (outFilter0[78]), .A1 (nx8606), .B0 (
         outFilter1[78]), .B1 (nx8716)) ;
    ao22 ix2405 (.Y (FilterToAlu_79), .A0 (outFilter0[79]), .A1 (nx8606), .B0 (
         outFilter1[79]), .B1 (nx8716)) ;
    ao22 ix2231 (.Y (FilterToAlu_80), .A0 (outFilter0[80]), .A1 (nx8606), .B0 (
         outFilter1[80]), .B1 (nx8716)) ;
    ao22 ix2237 (.Y (FilterToAlu_81), .A0 (outFilter0[81]), .A1 (nx8606), .B0 (
         outFilter1[81]), .B1 (nx8716)) ;
    ao22 ix2243 (.Y (FilterToAlu_82), .A0 (outFilter0[82]), .A1 (nx8608), .B0 (
         outFilter1[82]), .B1 (nx8718)) ;
    ao22 ix2249 (.Y (FilterToAlu_83), .A0 (outFilter0[83]), .A1 (nx8608), .B0 (
         outFilter1[83]), .B1 (nx8718)) ;
    ao22 ix2255 (.Y (FilterToAlu_84), .A0 (outFilter0[84]), .A1 (nx8608), .B0 (
         outFilter1[84]), .B1 (nx8718)) ;
    ao22 ix2261 (.Y (FilterToAlu_85), .A0 (outFilter0[85]), .A1 (nx8608), .B0 (
         outFilter1[85]), .B1 (nx8718)) ;
    ao22 ix2267 (.Y (FilterToAlu_86), .A0 (outFilter0[86]), .A1 (nx8608), .B0 (
         outFilter1[86]), .B1 (nx8718)) ;
    ao22 ix2273 (.Y (FilterToAlu_87), .A0 (outFilter0[87]), .A1 (nx8608), .B0 (
         outFilter1[87]), .B1 (nx8718)) ;
    ao22 ix2279 (.Y (FilterToAlu_88), .A0 (outFilter0[88]), .A1 (nx8608), .B0 (
         outFilter1[88]), .B1 (nx8718)) ;
    nand02 ix455 (.Y (FilterToAlu_89), .A0 (nx8144), .A1 (nx8924)) ;
    mux21 ix8145 (.Y (nx8144), .A0 (outFilter0[89]), .A1 (outFilter1[89]), .S0 (
          nx8896)) ;
    ao22 ix2285 (.Y (FilterToAlu_90), .A0 (outFilter0[90]), .A1 (nx8610), .B0 (
         outFilter1[90]), .B1 (nx8720)) ;
    ao22 ix2291 (.Y (FilterToAlu_91), .A0 (outFilter0[91]), .A1 (nx8610), .B0 (
         outFilter1[91]), .B1 (nx8720)) ;
    ao22 ix2297 (.Y (FilterToAlu_92), .A0 (outFilter0[92]), .A1 (nx8610), .B0 (
         outFilter1[92]), .B1 (nx8720)) ;
    ao22 ix2303 (.Y (FilterToAlu_93), .A0 (outFilter0[93]), .A1 (nx8610), .B0 (
         outFilter1[93]), .B1 (nx8720)) ;
    ao22 ix2309 (.Y (FilterToAlu_94), .A0 (outFilter0[94]), .A1 (nx8610), .B0 (
         outFilter1[94]), .B1 (nx8720)) ;
    ao22 ix2315 (.Y (FilterToAlu_95), .A0 (outFilter0[95]), .A1 (nx8610), .B0 (
         outFilter1[95]), .B1 (nx8720)) ;
    ao22 ix2141 (.Y (FilterToAlu_96), .A0 (outFilter0[96]), .A1 (nx8610), .B0 (
         outFilter1[96]), .B1 (nx8720)) ;
    ao22 ix2147 (.Y (FilterToAlu_97), .A0 (outFilter0[97]), .A1 (nx8612), .B0 (
         outFilter1[97]), .B1 (nx8722)) ;
    ao22 ix2153 (.Y (FilterToAlu_98), .A0 (outFilter0[98]), .A1 (nx8612), .B0 (
         outFilter1[98]), .B1 (nx8722)) ;
    ao22 ix2159 (.Y (FilterToAlu_99), .A0 (outFilter0[99]), .A1 (nx8612), .B0 (
         outFilter1[99]), .B1 (nx8722)) ;
    ao22 ix2165 (.Y (FilterToAlu_100), .A0 (outFilter0[100]), .A1 (nx8612), .B0 (
         outFilter1[100]), .B1 (nx8722)) ;
    ao22 ix2171 (.Y (FilterToAlu_101), .A0 (outFilter0[101]), .A1 (nx8612), .B0 (
         outFilter1[101]), .B1 (nx8722)) ;
    ao22 ix2177 (.Y (FilterToAlu_102), .A0 (outFilter0[102]), .A1 (nx8612), .B0 (
         outFilter1[102]), .B1 (nx8722)) ;
    ao22 ix2183 (.Y (FilterToAlu_103), .A0 (outFilter0[103]), .A1 (nx8612), .B0 (
         outFilter1[103]), .B1 (nx8722)) ;
    ao22 ix2189 (.Y (FilterToAlu_104), .A0 (outFilter0[104]), .A1 (nx8614), .B0 (
         outFilter1[104]), .B1 (nx8724)) ;
    nand02 ix445 (.Y (FilterToAlu_105), .A0 (nx8162), .A1 (nx8924)) ;
    mux21 ix8163 (.Y (nx8162), .A0 (outFilter0[105]), .A1 (outFilter1[105]), .S0 (
          nx8898)) ;
    ao22 ix2195 (.Y (FilterToAlu_106), .A0 (outFilter0[106]), .A1 (nx8614), .B0 (
         outFilter1[106]), .B1 (nx8724)) ;
    ao22 ix2201 (.Y (FilterToAlu_107), .A0 (outFilter0[107]), .A1 (nx8614), .B0 (
         outFilter1[107]), .B1 (nx8724)) ;
    ao22 ix2207 (.Y (FilterToAlu_108), .A0 (outFilter0[108]), .A1 (nx8614), .B0 (
         outFilter1[108]), .B1 (nx8724)) ;
    ao22 ix2213 (.Y (FilterToAlu_109), .A0 (outFilter0[109]), .A1 (nx8614), .B0 (
         outFilter1[109]), .B1 (nx8724)) ;
    ao22 ix2219 (.Y (FilterToAlu_110), .A0 (outFilter0[110]), .A1 (nx8614), .B0 (
         outFilter1[110]), .B1 (nx8724)) ;
    ao22 ix2225 (.Y (FilterToAlu_111), .A0 (outFilter0[111]), .A1 (nx8614), .B0 (
         outFilter1[111]), .B1 (nx8724)) ;
    ao22 ix2051 (.Y (FilterToAlu_112), .A0 (outFilter0[112]), .A1 (nx8616), .B0 (
         outFilter1[112]), .B1 (nx8726)) ;
    ao22 ix2057 (.Y (FilterToAlu_113), .A0 (outFilter0[113]), .A1 (nx8616), .B0 (
         outFilter1[113]), .B1 (nx8726)) ;
    ao22 ix2063 (.Y (FilterToAlu_114), .A0 (outFilter0[114]), .A1 (nx8616), .B0 (
         outFilter1[114]), .B1 (nx8726)) ;
    ao22 ix2069 (.Y (FilterToAlu_115), .A0 (outFilter0[115]), .A1 (nx8616), .B0 (
         outFilter1[115]), .B1 (nx8726)) ;
    ao22 ix2075 (.Y (FilterToAlu_116), .A0 (outFilter0[116]), .A1 (nx8616), .B0 (
         outFilter1[116]), .B1 (nx8726)) ;
    ao22 ix2081 (.Y (FilterToAlu_117), .A0 (outFilter0[117]), .A1 (nx8616), .B0 (
         outFilter1[117]), .B1 (nx8726)) ;
    ao22 ix2087 (.Y (FilterToAlu_118), .A0 (outFilter0[118]), .A1 (nx8616), .B0 (
         outFilter1[118]), .B1 (nx8726)) ;
    ao22 ix2093 (.Y (FilterToAlu_119), .A0 (outFilter0[119]), .A1 (nx8618), .B0 (
         outFilter1[119]), .B1 (nx8728)) ;
    ao22 ix2099 (.Y (FilterToAlu_120), .A0 (outFilter0[120]), .A1 (nx8618), .B0 (
         outFilter1[120]), .B1 (nx8728)) ;
    nand02 ix435 (.Y (FilterToAlu_121), .A0 (nx8180), .A1 (nx8806)) ;
    mux21 ix8181 (.Y (nx8180), .A0 (outFilter0[121]), .A1 (outFilter1[121]), .S0 (
          nx8898)) ;
    ao22 ix2105 (.Y (FilterToAlu_122), .A0 (outFilter0[122]), .A1 (nx8618), .B0 (
         outFilter1[122]), .B1 (nx8728)) ;
    ao22 ix2111 (.Y (FilterToAlu_123), .A0 (outFilter0[123]), .A1 (nx8618), .B0 (
         outFilter1[123]), .B1 (nx8728)) ;
    ao22 ix2117 (.Y (FilterToAlu_124), .A0 (outFilter0[124]), .A1 (nx8618), .B0 (
         outFilter1[124]), .B1 (nx8728)) ;
    ao22 ix2123 (.Y (FilterToAlu_125), .A0 (outFilter0[125]), .A1 (nx8618), .B0 (
         outFilter1[125]), .B1 (nx8728)) ;
    ao22 ix2129 (.Y (FilterToAlu_126), .A0 (outFilter0[126]), .A1 (nx8618), .B0 (
         outFilter1[126]), .B1 (nx8728)) ;
    ao22 ix2135 (.Y (FilterToAlu_127), .A0 (outFilter0[127]), .A1 (nx8620), .B0 (
         outFilter1[127]), .B1 (nx8730)) ;
    ao22 ix1961 (.Y (FilterToAlu_128), .A0 (outFilter0[128]), .A1 (nx8620), .B0 (
         outFilter1[128]), .B1 (nx8730)) ;
    ao22 ix1967 (.Y (FilterToAlu_129), .A0 (outFilter0[129]), .A1 (nx8620), .B0 (
         outFilter1[129]), .B1 (nx8730)) ;
    ao22 ix1973 (.Y (FilterToAlu_130), .A0 (outFilter0[130]), .A1 (nx8620), .B0 (
         outFilter1[130]), .B1 (nx8730)) ;
    ao22 ix1979 (.Y (FilterToAlu_131), .A0 (outFilter0[131]), .A1 (nx8620), .B0 (
         outFilter1[131]), .B1 (nx8730)) ;
    ao22 ix1985 (.Y (FilterToAlu_132), .A0 (outFilter0[132]), .A1 (nx8620), .B0 (
         outFilter1[132]), .B1 (nx8730)) ;
    ao22 ix1991 (.Y (FilterToAlu_133), .A0 (outFilter0[133]), .A1 (nx8620), .B0 (
         outFilter1[133]), .B1 (nx8730)) ;
    ao22 ix1997 (.Y (FilterToAlu_134), .A0 (outFilter0[134]), .A1 (nx8622), .B0 (
         outFilter1[134]), .B1 (nx8732)) ;
    ao22 ix2003 (.Y (FilterToAlu_135), .A0 (outFilter0[135]), .A1 (nx8622), .B0 (
         outFilter1[135]), .B1 (nx8732)) ;
    ao22 ix2009 (.Y (FilterToAlu_136), .A0 (outFilter0[136]), .A1 (nx8622), .B0 (
         outFilter1[136]), .B1 (nx8732)) ;
    nand02 ix425 (.Y (FilterToAlu_137), .A0 (nx8198), .A1 (nx8806)) ;
    mux21 ix8199 (.Y (nx8198), .A0 (outFilter0[137]), .A1 (outFilter1[137]), .S0 (
          nx8898)) ;
    ao22 ix2015 (.Y (FilterToAlu_138), .A0 (outFilter0[138]), .A1 (nx8622), .B0 (
         outFilter1[138]), .B1 (nx8732)) ;
    ao22 ix2021 (.Y (FilterToAlu_139), .A0 (outFilter0[139]), .A1 (nx8622), .B0 (
         outFilter1[139]), .B1 (nx8732)) ;
    ao22 ix2027 (.Y (FilterToAlu_140), .A0 (outFilter0[140]), .A1 (nx8622), .B0 (
         outFilter1[140]), .B1 (nx8732)) ;
    ao22 ix2033 (.Y (FilterToAlu_141), .A0 (outFilter0[141]), .A1 (nx8622), .B0 (
         outFilter1[141]), .B1 (nx8732)) ;
    ao22 ix2039 (.Y (FilterToAlu_142), .A0 (outFilter0[142]), .A1 (nx8624), .B0 (
         outFilter1[142]), .B1 (nx8734)) ;
    ao22 ix2045 (.Y (FilterToAlu_143), .A0 (outFilter0[143]), .A1 (nx8624), .B0 (
         outFilter1[143]), .B1 (nx8734)) ;
    ao22 ix1871 (.Y (FilterToAlu_144), .A0 (outFilter0[144]), .A1 (nx8624), .B0 (
         outFilter1[144]), .B1 (nx8734)) ;
    ao22 ix1877 (.Y (FilterToAlu_145), .A0 (outFilter0[145]), .A1 (nx8624), .B0 (
         outFilter1[145]), .B1 (nx8734)) ;
    ao22 ix1883 (.Y (FilterToAlu_146), .A0 (outFilter0[146]), .A1 (nx8624), .B0 (
         outFilter1[146]), .B1 (nx8734)) ;
    ao22 ix1889 (.Y (FilterToAlu_147), .A0 (outFilter0[147]), .A1 (nx8624), .B0 (
         outFilter1[147]), .B1 (nx8734)) ;
    ao22 ix1895 (.Y (FilterToAlu_148), .A0 (outFilter0[148]), .A1 (nx8624), .B0 (
         outFilter1[148]), .B1 (nx8734)) ;
    ao22 ix1901 (.Y (FilterToAlu_149), .A0 (outFilter0[149]), .A1 (nx8626), .B0 (
         outFilter1[149]), .B1 (nx8736)) ;
    ao22 ix1907 (.Y (FilterToAlu_150), .A0 (outFilter0[150]), .A1 (nx8626), .B0 (
         outFilter1[150]), .B1 (nx8736)) ;
    ao22 ix1913 (.Y (FilterToAlu_151), .A0 (outFilter0[151]), .A1 (nx8626), .B0 (
         outFilter1[151]), .B1 (nx8736)) ;
    ao22 ix1919 (.Y (FilterToAlu_152), .A0 (outFilter0[152]), .A1 (nx8626), .B0 (
         outFilter1[152]), .B1 (nx8736)) ;
    nand02 ix415 (.Y (FilterToAlu_153), .A0 (nx8216), .A1 (nx8806)) ;
    mux21 ix8217 (.Y (nx8216), .A0 (outFilter0[153]), .A1 (outFilter1[153]), .S0 (
          nx8898)) ;
    ao22 ix1925 (.Y (FilterToAlu_154), .A0 (outFilter0[154]), .A1 (nx8626), .B0 (
         outFilter1[154]), .B1 (nx8736)) ;
    ao22 ix1931 (.Y (FilterToAlu_155), .A0 (outFilter0[155]), .A1 (nx8626), .B0 (
         outFilter1[155]), .B1 (nx8736)) ;
    ao22 ix1937 (.Y (FilterToAlu_156), .A0 (outFilter0[156]), .A1 (nx8626), .B0 (
         outFilter1[156]), .B1 (nx8736)) ;
    ao22 ix1943 (.Y (FilterToAlu_157), .A0 (outFilter0[157]), .A1 (nx8628), .B0 (
         outFilter1[157]), .B1 (nx8738)) ;
    ao22 ix1949 (.Y (FilterToAlu_158), .A0 (outFilter0[158]), .A1 (nx8628), .B0 (
         outFilter1[158]), .B1 (nx8738)) ;
    ao22 ix1955 (.Y (FilterToAlu_159), .A0 (outFilter0[159]), .A1 (nx8628), .B0 (
         outFilter1[159]), .B1 (nx8738)) ;
    ao22 ix1781 (.Y (FilterToAlu_160), .A0 (outFilter0[160]), .A1 (nx8628), .B0 (
         outFilter1[160]), .B1 (nx8738)) ;
    ao22 ix1787 (.Y (FilterToAlu_161), .A0 (outFilter0[161]), .A1 (nx8628), .B0 (
         outFilter1[161]), .B1 (nx8738)) ;
    ao22 ix1793 (.Y (FilterToAlu_162), .A0 (outFilter0[162]), .A1 (nx8628), .B0 (
         outFilter1[162]), .B1 (nx8738)) ;
    ao22 ix1799 (.Y (FilterToAlu_163), .A0 (outFilter0[163]), .A1 (nx8628), .B0 (
         outFilter1[163]), .B1 (nx8738)) ;
    ao22 ix1805 (.Y (FilterToAlu_164), .A0 (outFilter0[164]), .A1 (nx8630), .B0 (
         outFilter1[164]), .B1 (nx8740)) ;
    ao22 ix1811 (.Y (FilterToAlu_165), .A0 (outFilter0[165]), .A1 (nx8630), .B0 (
         outFilter1[165]), .B1 (nx8740)) ;
    ao22 ix1817 (.Y (FilterToAlu_166), .A0 (outFilter0[166]), .A1 (nx8630), .B0 (
         outFilter1[166]), .B1 (nx8740)) ;
    ao22 ix1823 (.Y (FilterToAlu_167), .A0 (outFilter0[167]), .A1 (nx8630), .B0 (
         outFilter1[167]), .B1 (nx8740)) ;
    ao22 ix1829 (.Y (FilterToAlu_168), .A0 (outFilter0[168]), .A1 (nx8630), .B0 (
         outFilter1[168]), .B1 (nx8740)) ;
    nand02 ix405 (.Y (FilterToAlu_169), .A0 (nx8234), .A1 (nx8806)) ;
    mux21 ix8235 (.Y (nx8234), .A0 (outFilter0[169]), .A1 (outFilter1[169]), .S0 (
          nx8898)) ;
    ao22 ix1835 (.Y (FilterToAlu_170), .A0 (outFilter0[170]), .A1 (nx8630), .B0 (
         outFilter1[170]), .B1 (nx8740)) ;
    ao22 ix1841 (.Y (FilterToAlu_171), .A0 (outFilter0[171]), .A1 (nx8630), .B0 (
         outFilter1[171]), .B1 (nx8740)) ;
    ao22 ix1847 (.Y (FilterToAlu_172), .A0 (outFilter0[172]), .A1 (nx8632), .B0 (
         outFilter1[172]), .B1 (nx8742)) ;
    ao22 ix1853 (.Y (FilterToAlu_173), .A0 (outFilter0[173]), .A1 (nx8632), .B0 (
         outFilter1[173]), .B1 (nx8742)) ;
    ao22 ix1859 (.Y (FilterToAlu_174), .A0 (outFilter0[174]), .A1 (nx8632), .B0 (
         outFilter1[174]), .B1 (nx8742)) ;
    ao22 ix1865 (.Y (FilterToAlu_175), .A0 (outFilter0[175]), .A1 (nx8632), .B0 (
         outFilter1[175]), .B1 (nx8742)) ;
    ao22 ix1691 (.Y (FilterToAlu_176), .A0 (outFilter0[176]), .A1 (nx8632), .B0 (
         outFilter1[176]), .B1 (nx8742)) ;
    ao22 ix1697 (.Y (FilterToAlu_177), .A0 (outFilter0[177]), .A1 (nx8632), .B0 (
         outFilter1[177]), .B1 (nx8742)) ;
    ao22 ix1703 (.Y (FilterToAlu_178), .A0 (outFilter0[178]), .A1 (nx8632), .B0 (
         outFilter1[178]), .B1 (nx8742)) ;
    ao22 ix1709 (.Y (FilterToAlu_179), .A0 (outFilter0[179]), .A1 (nx8634), .B0 (
         outFilter1[179]), .B1 (nx8744)) ;
    ao22 ix1715 (.Y (FilterToAlu_180), .A0 (outFilter0[180]), .A1 (nx8634), .B0 (
         outFilter1[180]), .B1 (nx8744)) ;
    ao22 ix1721 (.Y (FilterToAlu_181), .A0 (outFilter0[181]), .A1 (nx8634), .B0 (
         outFilter1[181]), .B1 (nx8744)) ;
    ao22 ix1727 (.Y (FilterToAlu_182), .A0 (outFilter0[182]), .A1 (nx8634), .B0 (
         outFilter1[182]), .B1 (nx8744)) ;
    ao22 ix1733 (.Y (FilterToAlu_183), .A0 (outFilter0[183]), .A1 (nx8634), .B0 (
         outFilter1[183]), .B1 (nx8744)) ;
    ao22 ix1739 (.Y (FilterToAlu_184), .A0 (outFilter0[184]), .A1 (nx8634), .B0 (
         outFilter1[184]), .B1 (nx8744)) ;
    nand02 ix395 (.Y (FilterToAlu_185), .A0 (nx8252), .A1 (nx8806)) ;
    mux21 ix8253 (.Y (nx8252), .A0 (outFilter0[185]), .A1 (outFilter1[185]), .S0 (
          nx8898)) ;
    ao22 ix1745 (.Y (FilterToAlu_186), .A0 (outFilter0[186]), .A1 (nx8634), .B0 (
         outFilter1[186]), .B1 (nx8744)) ;
    ao22 ix1751 (.Y (FilterToAlu_187), .A0 (outFilter0[187]), .A1 (nx8636), .B0 (
         outFilter1[187]), .B1 (nx8746)) ;
    ao22 ix1757 (.Y (FilterToAlu_188), .A0 (outFilter0[188]), .A1 (nx8636), .B0 (
         outFilter1[188]), .B1 (nx8746)) ;
    ao22 ix1763 (.Y (FilterToAlu_189), .A0 (outFilter0[189]), .A1 (nx8636), .B0 (
         outFilter1[189]), .B1 (nx8746)) ;
    ao22 ix1769 (.Y (FilterToAlu_190), .A0 (outFilter0[190]), .A1 (nx8636), .B0 (
         outFilter1[190]), .B1 (nx8746)) ;
    ao22 ix1775 (.Y (FilterToAlu_191), .A0 (outFilter0[191]), .A1 (nx8636), .B0 (
         outFilter1[191]), .B1 (nx8746)) ;
    ao22 ix1601 (.Y (FilterToAlu_192), .A0 (outFilter0[192]), .A1 (nx8636), .B0 (
         outFilter1[192]), .B1 (nx8746)) ;
    ao22 ix1607 (.Y (FilterToAlu_193), .A0 (outFilter0[193]), .A1 (nx8636), .B0 (
         outFilter1[193]), .B1 (nx8746)) ;
    ao22 ix1613 (.Y (FilterToAlu_194), .A0 (outFilter0[194]), .A1 (nx8638), .B0 (
         outFilter1[194]), .B1 (nx8748)) ;
    ao22 ix1619 (.Y (FilterToAlu_195), .A0 (outFilter0[195]), .A1 (nx8638), .B0 (
         outFilter1[195]), .B1 (nx8748)) ;
    ao22 ix1625 (.Y (FilterToAlu_196), .A0 (outFilter0[196]), .A1 (nx8638), .B0 (
         outFilter1[196]), .B1 (nx8748)) ;
    ao22 ix1631 (.Y (FilterToAlu_197), .A0 (outFilter0[197]), .A1 (nx8638), .B0 (
         outFilter1[197]), .B1 (nx8748)) ;
    ao22 ix1637 (.Y (FilterToAlu_198), .A0 (outFilter0[198]), .A1 (nx8638), .B0 (
         outFilter1[198]), .B1 (nx8748)) ;
    ao22 ix1643 (.Y (FilterToAlu_199), .A0 (outFilter0[199]), .A1 (nx8638), .B0 (
         outFilter1[199]), .B1 (nx8748)) ;
    ao22 ix1649 (.Y (FilterToAlu_200), .A0 (outFilter0[200]), .A1 (nx8638), .B0 (
         outFilter1[200]), .B1 (nx8748)) ;
    nand02 ix385 (.Y (FilterToAlu_201), .A0 (nx8270), .A1 (nx8806)) ;
    mux21 ix8271 (.Y (nx8270), .A0 (outFilter0[201]), .A1 (outFilter1[201]), .S0 (
          nx8898)) ;
    ao22 ix1655 (.Y (FilterToAlu_202), .A0 (outFilter0[202]), .A1 (nx8640), .B0 (
         outFilter1[202]), .B1 (nx8750)) ;
    ao22 ix1661 (.Y (FilterToAlu_203), .A0 (outFilter0[203]), .A1 (nx8640), .B0 (
         outFilter1[203]), .B1 (nx8750)) ;
    ao22 ix1667 (.Y (FilterToAlu_204), .A0 (outFilter0[204]), .A1 (nx8640), .B0 (
         outFilter1[204]), .B1 (nx8750)) ;
    ao22 ix1673 (.Y (FilterToAlu_205), .A0 (outFilter0[205]), .A1 (nx8640), .B0 (
         outFilter1[205]), .B1 (nx8750)) ;
    ao22 ix1679 (.Y (FilterToAlu_206), .A0 (outFilter0[206]), .A1 (nx8640), .B0 (
         outFilter1[206]), .B1 (nx8750)) ;
    ao22 ix1685 (.Y (FilterToAlu_207), .A0 (outFilter0[207]), .A1 (nx8640), .B0 (
         outFilter1[207]), .B1 (nx8750)) ;
    ao22 ix1511 (.Y (FilterToAlu_208), .A0 (outFilter0[208]), .A1 (nx8640), .B0 (
         outFilter1[208]), .B1 (nx8750)) ;
    ao22 ix1517 (.Y (FilterToAlu_209), .A0 (outFilter0[209]), .A1 (nx8642), .B0 (
         outFilter1[209]), .B1 (nx8752)) ;
    ao22 ix1523 (.Y (FilterToAlu_210), .A0 (outFilter0[210]), .A1 (nx8642), .B0 (
         outFilter1[210]), .B1 (nx8752)) ;
    ao22 ix1529 (.Y (FilterToAlu_211), .A0 (outFilter0[211]), .A1 (nx8642), .B0 (
         outFilter1[211]), .B1 (nx8752)) ;
    ao22 ix1535 (.Y (FilterToAlu_212), .A0 (outFilter0[212]), .A1 (nx8642), .B0 (
         outFilter1[212]), .B1 (nx8752)) ;
    ao22 ix1541 (.Y (FilterToAlu_213), .A0 (outFilter0[213]), .A1 (nx8642), .B0 (
         outFilter1[213]), .B1 (nx8752)) ;
    ao22 ix1547 (.Y (FilterToAlu_214), .A0 (outFilter0[214]), .A1 (nx8642), .B0 (
         outFilter1[214]), .B1 (nx8752)) ;
    ao22 ix1553 (.Y (FilterToAlu_215), .A0 (outFilter0[215]), .A1 (nx8642), .B0 (
         outFilter1[215]), .B1 (nx8752)) ;
    ao22 ix1559 (.Y (FilterToAlu_216), .A0 (outFilter0[216]), .A1 (nx8644), .B0 (
         outFilter1[216]), .B1 (nx8754)) ;
    nand02 ix375 (.Y (FilterToAlu_217), .A0 (nx8288), .A1 (nx8806)) ;
    mux21 ix8289 (.Y (nx8288), .A0 (outFilter0[217]), .A1 (outFilter1[217]), .S0 (
          nx8900)) ;
    ao22 ix1565 (.Y (FilterToAlu_218), .A0 (outFilter0[218]), .A1 (nx8644), .B0 (
         outFilter1[218]), .B1 (nx8754)) ;
    ao22 ix1571 (.Y (FilterToAlu_219), .A0 (outFilter0[219]), .A1 (nx8644), .B0 (
         outFilter1[219]), .B1 (nx8754)) ;
    ao22 ix1577 (.Y (FilterToAlu_220), .A0 (outFilter0[220]), .A1 (nx8644), .B0 (
         outFilter1[220]), .B1 (nx8754)) ;
    ao22 ix1583 (.Y (FilterToAlu_221), .A0 (outFilter0[221]), .A1 (nx8644), .B0 (
         outFilter1[221]), .B1 (nx8754)) ;
    ao22 ix1589 (.Y (FilterToAlu_222), .A0 (outFilter0[222]), .A1 (nx8644), .B0 (
         outFilter1[222]), .B1 (nx8754)) ;
    ao22 ix1595 (.Y (FilterToAlu_223), .A0 (outFilter0[223]), .A1 (nx8644), .B0 (
         outFilter1[223]), .B1 (nx8754)) ;
    ao22 ix1421 (.Y (FilterToAlu_224), .A0 (outFilter0[224]), .A1 (nx8646), .B0 (
         outFilter1[224]), .B1 (nx8756)) ;
    ao22 ix1427 (.Y (FilterToAlu_225), .A0 (outFilter0[225]), .A1 (nx8646), .B0 (
         outFilter1[225]), .B1 (nx8756)) ;
    ao22 ix1433 (.Y (FilterToAlu_226), .A0 (outFilter0[226]), .A1 (nx8646), .B0 (
         outFilter1[226]), .B1 (nx8756)) ;
    ao22 ix1439 (.Y (FilterToAlu_227), .A0 (outFilter0[227]), .A1 (nx8646), .B0 (
         outFilter1[227]), .B1 (nx8756)) ;
    ao22 ix1445 (.Y (FilterToAlu_228), .A0 (outFilter0[228]), .A1 (nx8646), .B0 (
         outFilter1[228]), .B1 (nx8756)) ;
    ao22 ix1451 (.Y (FilterToAlu_229), .A0 (outFilter0[229]), .A1 (nx8646), .B0 (
         outFilter1[229]), .B1 (nx8756)) ;
    ao22 ix1457 (.Y (FilterToAlu_230), .A0 (outFilter0[230]), .A1 (nx8646), .B0 (
         outFilter1[230]), .B1 (nx8756)) ;
    ao22 ix1463 (.Y (FilterToAlu_231), .A0 (outFilter0[231]), .A1 (nx8648), .B0 (
         outFilter1[231]), .B1 (nx8758)) ;
    ao22 ix1469 (.Y (FilterToAlu_232), .A0 (outFilter0[232]), .A1 (nx8648), .B0 (
         outFilter1[232]), .B1 (nx8758)) ;
    nand02 ix365 (.Y (FilterToAlu_233), .A0 (nx8306), .A1 (nx8808)) ;
    mux21 ix8307 (.Y (nx8306), .A0 (outFilter0[233]), .A1 (outFilter1[233]), .S0 (
          nx8900)) ;
    ao22 ix1475 (.Y (FilterToAlu_234), .A0 (outFilter0[234]), .A1 (nx8648), .B0 (
         outFilter1[234]), .B1 (nx8758)) ;
    ao22 ix1481 (.Y (FilterToAlu_235), .A0 (outFilter0[235]), .A1 (nx8648), .B0 (
         outFilter1[235]), .B1 (nx8758)) ;
    ao22 ix1487 (.Y (FilterToAlu_236), .A0 (outFilter0[236]), .A1 (nx8648), .B0 (
         outFilter1[236]), .B1 (nx8758)) ;
    ao22 ix1493 (.Y (FilterToAlu_237), .A0 (outFilter0[237]), .A1 (nx8648), .B0 (
         outFilter1[237]), .B1 (nx8758)) ;
    ao22 ix1499 (.Y (FilterToAlu_238), .A0 (outFilter0[238]), .A1 (nx8648), .B0 (
         outFilter1[238]), .B1 (nx8758)) ;
    ao22 ix1505 (.Y (FilterToAlu_239), .A0 (outFilter0[239]), .A1 (nx8650), .B0 (
         outFilter1[239]), .B1 (nx8760)) ;
    ao22 ix1331 (.Y (FilterToAlu_240), .A0 (outFilter0[240]), .A1 (nx8650), .B0 (
         outFilter1[240]), .B1 (nx8760)) ;
    ao22 ix1337 (.Y (FilterToAlu_241), .A0 (outFilter0[241]), .A1 (nx8650), .B0 (
         outFilter1[241]), .B1 (nx8760)) ;
    ao22 ix1343 (.Y (FilterToAlu_242), .A0 (outFilter0[242]), .A1 (nx8650), .B0 (
         outFilter1[242]), .B1 (nx8760)) ;
    ao22 ix1349 (.Y (FilterToAlu_243), .A0 (outFilter0[243]), .A1 (nx8650), .B0 (
         outFilter1[243]), .B1 (nx8760)) ;
    ao22 ix1355 (.Y (FilterToAlu_244), .A0 (outFilter0[244]), .A1 (nx8650), .B0 (
         outFilter1[244]), .B1 (nx8760)) ;
    ao22 ix1361 (.Y (FilterToAlu_245), .A0 (outFilter0[245]), .A1 (nx8650), .B0 (
         outFilter1[245]), .B1 (nx8760)) ;
    ao22 ix1367 (.Y (FilterToAlu_246), .A0 (outFilter0[246]), .A1 (nx8652), .B0 (
         outFilter1[246]), .B1 (nx8762)) ;
    ao22 ix1373 (.Y (FilterToAlu_247), .A0 (outFilter0[247]), .A1 (nx8652), .B0 (
         outFilter1[247]), .B1 (nx8762)) ;
    ao22 ix1379 (.Y (FilterToAlu_248), .A0 (outFilter0[248]), .A1 (nx8652), .B0 (
         outFilter1[248]), .B1 (nx8762)) ;
    nand02 ix355 (.Y (FilterToAlu_249), .A0 (nx8324), .A1 (nx8808)) ;
    mux21 ix8325 (.Y (nx8324), .A0 (outFilter0[249]), .A1 (outFilter1[249]), .S0 (
          nx8900)) ;
    ao22 ix1385 (.Y (FilterToAlu_250), .A0 (outFilter0[250]), .A1 (nx8652), .B0 (
         outFilter1[250]), .B1 (nx8762)) ;
    ao22 ix1391 (.Y (FilterToAlu_251), .A0 (outFilter0[251]), .A1 (nx8652), .B0 (
         outFilter1[251]), .B1 (nx8762)) ;
    ao22 ix1397 (.Y (FilterToAlu_252), .A0 (outFilter0[252]), .A1 (nx8652), .B0 (
         outFilter1[252]), .B1 (nx8762)) ;
    ao22 ix1403 (.Y (FilterToAlu_253), .A0 (outFilter0[253]), .A1 (nx8652), .B0 (
         outFilter1[253]), .B1 (nx8762)) ;
    ao22 ix1409 (.Y (FilterToAlu_254), .A0 (outFilter0[254]), .A1 (nx8654), .B0 (
         outFilter1[254]), .B1 (nx8764)) ;
    ao22 ix1415 (.Y (FilterToAlu_255), .A0 (outFilter0[255]), .A1 (nx8654), .B0 (
         outFilter1[255]), .B1 (nx8764)) ;
    ao22 ix1241 (.Y (FilterToAlu_256), .A0 (outFilter0[256]), .A1 (nx8654), .B0 (
         outFilter1[256]), .B1 (nx8764)) ;
    ao22 ix1247 (.Y (FilterToAlu_257), .A0 (outFilter0[257]), .A1 (nx8654), .B0 (
         outFilter1[257]), .B1 (nx8764)) ;
    ao22 ix1253 (.Y (FilterToAlu_258), .A0 (outFilter0[258]), .A1 (nx8654), .B0 (
         outFilter1[258]), .B1 (nx8764)) ;
    ao22 ix1259 (.Y (FilterToAlu_259), .A0 (outFilter0[259]), .A1 (nx8654), .B0 (
         outFilter1[259]), .B1 (nx8764)) ;
    ao22 ix1265 (.Y (FilterToAlu_260), .A0 (outFilter0[260]), .A1 (nx8654), .B0 (
         outFilter1[260]), .B1 (nx8764)) ;
    ao22 ix1271 (.Y (FilterToAlu_261), .A0 (outFilter0[261]), .A1 (nx8656), .B0 (
         outFilter1[261]), .B1 (nx8766)) ;
    ao22 ix1277 (.Y (FilterToAlu_262), .A0 (outFilter0[262]), .A1 (nx8656), .B0 (
         outFilter1[262]), .B1 (nx8766)) ;
    ao22 ix1283 (.Y (FilterToAlu_263), .A0 (outFilter0[263]), .A1 (nx8656), .B0 (
         outFilter1[263]), .B1 (nx8766)) ;
    ao22 ix1289 (.Y (FilterToAlu_264), .A0 (outFilter0[264]), .A1 (nx8656), .B0 (
         outFilter1[264]), .B1 (nx8766)) ;
    nand02 ix345 (.Y (FilterToAlu_265), .A0 (nx8342), .A1 (nx8808)) ;
    mux21 ix8343 (.Y (nx8342), .A0 (outFilter0[265]), .A1 (outFilter1[265]), .S0 (
          nx8900)) ;
    ao22 ix1295 (.Y (FilterToAlu_266), .A0 (outFilter0[266]), .A1 (nx8656), .B0 (
         outFilter1[266]), .B1 (nx8766)) ;
    ao22 ix1301 (.Y (FilterToAlu_267), .A0 (outFilter0[267]), .A1 (nx8656), .B0 (
         outFilter1[267]), .B1 (nx8766)) ;
    ao22 ix1307 (.Y (FilterToAlu_268), .A0 (outFilter0[268]), .A1 (nx8656), .B0 (
         outFilter1[268]), .B1 (nx8766)) ;
    ao22 ix1313 (.Y (FilterToAlu_269), .A0 (outFilter0[269]), .A1 (nx8658), .B0 (
         outFilter1[269]), .B1 (nx8768)) ;
    ao22 ix1319 (.Y (FilterToAlu_270), .A0 (outFilter0[270]), .A1 (nx8658), .B0 (
         outFilter1[270]), .B1 (nx8768)) ;
    ao22 ix1325 (.Y (FilterToAlu_271), .A0 (outFilter0[271]), .A1 (nx8658), .B0 (
         outFilter1[271]), .B1 (nx8768)) ;
    ao22 ix1151 (.Y (FilterToAlu_272), .A0 (outFilter0[272]), .A1 (nx8658), .B0 (
         outFilter1[272]), .B1 (nx8768)) ;
    ao22 ix1157 (.Y (FilterToAlu_273), .A0 (outFilter0[273]), .A1 (nx8658), .B0 (
         outFilter1[273]), .B1 (nx8768)) ;
    ao22 ix1163 (.Y (FilterToAlu_274), .A0 (outFilter0[274]), .A1 (nx8658), .B0 (
         outFilter1[274]), .B1 (nx8768)) ;
    ao22 ix1169 (.Y (FilterToAlu_275), .A0 (outFilter0[275]), .A1 (nx8658), .B0 (
         outFilter1[275]), .B1 (nx8768)) ;
    ao22 ix1175 (.Y (FilterToAlu_276), .A0 (outFilter0[276]), .A1 (nx8660), .B0 (
         outFilter1[276]), .B1 (nx8770)) ;
    ao22 ix1181 (.Y (FilterToAlu_277), .A0 (outFilter0[277]), .A1 (nx8660), .B0 (
         outFilter1[277]), .B1 (nx8770)) ;
    ao22 ix1187 (.Y (FilterToAlu_278), .A0 (outFilter0[278]), .A1 (nx8660), .B0 (
         outFilter1[278]), .B1 (nx8770)) ;
    ao22 ix1193 (.Y (FilterToAlu_279), .A0 (outFilter0[279]), .A1 (nx8660), .B0 (
         outFilter1[279]), .B1 (nx8770)) ;
    ao22 ix1199 (.Y (FilterToAlu_280), .A0 (outFilter0[280]), .A1 (nx8660), .B0 (
         outFilter1[280]), .B1 (nx8770)) ;
    nand02 ix335 (.Y (FilterToAlu_281), .A0 (nx8360), .A1 (nx8808)) ;
    mux21 ix8361 (.Y (nx8360), .A0 (outFilter0[281]), .A1 (outFilter1[281]), .S0 (
          nx8900)) ;
    ao22 ix1205 (.Y (FilterToAlu_282), .A0 (outFilter0[282]), .A1 (nx8660), .B0 (
         outFilter1[282]), .B1 (nx8770)) ;
    ao22 ix1211 (.Y (FilterToAlu_283), .A0 (outFilter0[283]), .A1 (nx8660), .B0 (
         outFilter1[283]), .B1 (nx8770)) ;
    ao22 ix1217 (.Y (FilterToAlu_284), .A0 (outFilter0[284]), .A1 (nx8662), .B0 (
         outFilter1[284]), .B1 (nx8772)) ;
    ao22 ix1223 (.Y (FilterToAlu_285), .A0 (outFilter0[285]), .A1 (nx8662), .B0 (
         outFilter1[285]), .B1 (nx8772)) ;
    ao22 ix1229 (.Y (FilterToAlu_286), .A0 (outFilter0[286]), .A1 (nx8662), .B0 (
         outFilter1[286]), .B1 (nx8772)) ;
    ao22 ix1235 (.Y (FilterToAlu_287), .A0 (outFilter0[287]), .A1 (nx8662), .B0 (
         outFilter1[287]), .B1 (nx8772)) ;
    ao22 ix1061 (.Y (FilterToAlu_288), .A0 (outFilter0[288]), .A1 (nx8662), .B0 (
         outFilter1[288]), .B1 (nx8772)) ;
    ao22 ix1067 (.Y (FilterToAlu_289), .A0 (outFilter0[289]), .A1 (nx8662), .B0 (
         outFilter1[289]), .B1 (nx8772)) ;
    ao22 ix1073 (.Y (FilterToAlu_290), .A0 (outFilter0[290]), .A1 (nx8662), .B0 (
         outFilter1[290]), .B1 (nx8772)) ;
    ao22 ix1079 (.Y (FilterToAlu_291), .A0 (outFilter0[291]), .A1 (nx8664), .B0 (
         outFilter1[291]), .B1 (nx8774)) ;
    ao22 ix1085 (.Y (FilterToAlu_292), .A0 (outFilter0[292]), .A1 (nx8664), .B0 (
         outFilter1[292]), .B1 (nx8774)) ;
    ao22 ix1091 (.Y (FilterToAlu_293), .A0 (outFilter0[293]), .A1 (nx8664), .B0 (
         outFilter1[293]), .B1 (nx8774)) ;
    ao22 ix1097 (.Y (FilterToAlu_294), .A0 (outFilter0[294]), .A1 (nx8664), .B0 (
         outFilter1[294]), .B1 (nx8774)) ;
    ao22 ix1103 (.Y (FilterToAlu_295), .A0 (outFilter0[295]), .A1 (nx8664), .B0 (
         outFilter1[295]), .B1 (nx8774)) ;
    ao22 ix1109 (.Y (FilterToAlu_296), .A0 (outFilter0[296]), .A1 (nx8664), .B0 (
         outFilter1[296]), .B1 (nx8774)) ;
    nand02 ix325 (.Y (FilterToAlu_297), .A0 (nx8378), .A1 (nx8808)) ;
    mux21 ix8379 (.Y (nx8378), .A0 (outFilter0[297]), .A1 (outFilter1[297]), .S0 (
          nx8900)) ;
    ao22 ix1115 (.Y (FilterToAlu_298), .A0 (outFilter0[298]), .A1 (nx8664), .B0 (
         outFilter1[298]), .B1 (nx8774)) ;
    ao22 ix1121 (.Y (FilterToAlu_299), .A0 (outFilter0[299]), .A1 (nx8666), .B0 (
         outFilter1[299]), .B1 (nx8776)) ;
    ao22 ix1127 (.Y (FilterToAlu_300), .A0 (outFilter0[300]), .A1 (nx8666), .B0 (
         outFilter1[300]), .B1 (nx8776)) ;
    ao22 ix1133 (.Y (FilterToAlu_301), .A0 (outFilter0[301]), .A1 (nx8666), .B0 (
         outFilter1[301]), .B1 (nx8776)) ;
    ao22 ix1139 (.Y (FilterToAlu_302), .A0 (outFilter0[302]), .A1 (nx8666), .B0 (
         outFilter1[302]), .B1 (nx8776)) ;
    ao22 ix1145 (.Y (FilterToAlu_303), .A0 (outFilter0[303]), .A1 (nx8666), .B0 (
         outFilter1[303]), .B1 (nx8776)) ;
    ao22 ix971 (.Y (FilterToAlu_304), .A0 (outFilter0[304]), .A1 (nx8666), .B0 (
         outFilter1[304]), .B1 (nx8776)) ;
    ao22 ix977 (.Y (FilterToAlu_305), .A0 (outFilter0[305]), .A1 (nx8666), .B0 (
         outFilter1[305]), .B1 (nx8776)) ;
    ao22 ix983 (.Y (FilterToAlu_306), .A0 (outFilter0[306]), .A1 (nx8668), .B0 (
         outFilter1[306]), .B1 (nx8778)) ;
    ao22 ix989 (.Y (FilterToAlu_307), .A0 (outFilter0[307]), .A1 (nx8668), .B0 (
         outFilter1[307]), .B1 (nx8778)) ;
    ao22 ix995 (.Y (FilterToAlu_308), .A0 (outFilter0[308]), .A1 (nx8668), .B0 (
         outFilter1[308]), .B1 (nx8778)) ;
    ao22 ix1001 (.Y (FilterToAlu_309), .A0 (outFilter0[309]), .A1 (nx8668), .B0 (
         outFilter1[309]), .B1 (nx8778)) ;
    ao22 ix1007 (.Y (FilterToAlu_310), .A0 (outFilter0[310]), .A1 (nx8668), .B0 (
         outFilter1[310]), .B1 (nx8778)) ;
    ao22 ix1013 (.Y (FilterToAlu_311), .A0 (outFilter0[311]), .A1 (nx8668), .B0 (
         outFilter1[311]), .B1 (nx8778)) ;
    ao22 ix1019 (.Y (FilterToAlu_312), .A0 (outFilter0[312]), .A1 (nx8668), .B0 (
         outFilter1[312]), .B1 (nx8778)) ;
    nand02 ix315 (.Y (FilterToAlu_313), .A0 (nx8396), .A1 (nx8808)) ;
    mux21 ix8397 (.Y (nx8396), .A0 (outFilter0[313]), .A1 (outFilter1[313]), .S0 (
          nx8900)) ;
    ao22 ix1025 (.Y (FilterToAlu_314), .A0 (outFilter0[314]), .A1 (nx8670), .B0 (
         outFilter1[314]), .B1 (nx8780)) ;
    ao22 ix1031 (.Y (FilterToAlu_315), .A0 (outFilter0[315]), .A1 (nx8670), .B0 (
         outFilter1[315]), .B1 (nx8780)) ;
    ao22 ix1037 (.Y (FilterToAlu_316), .A0 (outFilter0[316]), .A1 (nx8670), .B0 (
         outFilter1[316]), .B1 (nx8780)) ;
    ao22 ix1043 (.Y (FilterToAlu_317), .A0 (outFilter0[317]), .A1 (nx8670), .B0 (
         outFilter1[317]), .B1 (nx8780)) ;
    ao22 ix1049 (.Y (FilterToAlu_318), .A0 (outFilter0[318]), .A1 (nx8670), .B0 (
         outFilter1[318]), .B1 (nx8780)) ;
    ao22 ix1055 (.Y (FilterToAlu_319), .A0 (outFilter0[319]), .A1 (nx8670), .B0 (
         outFilter1[319]), .B1 (nx8780)) ;
    ao22 ix881 (.Y (FilterToAlu_320), .A0 (outFilter0[320]), .A1 (nx8670), .B0 (
         outFilter1[320]), .B1 (nx8780)) ;
    ao22 ix887 (.Y (FilterToAlu_321), .A0 (outFilter0[321]), .A1 (nx8672), .B0 (
         outFilter1[321]), .B1 (nx8782)) ;
    ao22 ix893 (.Y (FilterToAlu_322), .A0 (outFilter0[322]), .A1 (nx8672), .B0 (
         outFilter1[322]), .B1 (nx8782)) ;
    ao22 ix899 (.Y (FilterToAlu_323), .A0 (outFilter0[323]), .A1 (nx8672), .B0 (
         outFilter1[323]), .B1 (nx8782)) ;
    ao22 ix905 (.Y (FilterToAlu_324), .A0 (outFilter0[324]), .A1 (nx8672), .B0 (
         outFilter1[324]), .B1 (nx8782)) ;
    ao22 ix911 (.Y (FilterToAlu_325), .A0 (outFilter0[325]), .A1 (nx8672), .B0 (
         outFilter1[325]), .B1 (nx8782)) ;
    ao22 ix917 (.Y (FilterToAlu_326), .A0 (outFilter0[326]), .A1 (nx8672), .B0 (
         outFilter1[326]), .B1 (nx8782)) ;
    ao22 ix923 (.Y (FilterToAlu_327), .A0 (outFilter0[327]), .A1 (nx8672), .B0 (
         outFilter1[327]), .B1 (nx8782)) ;
    ao22 ix929 (.Y (FilterToAlu_328), .A0 (outFilter0[328]), .A1 (nx8674), .B0 (
         outFilter1[328]), .B1 (nx8784)) ;
    nand02 ix305 (.Y (FilterToAlu_329), .A0 (nx8414), .A1 (nx8808)) ;
    mux21 ix8415 (.Y (nx8414), .A0 (outFilter0[329]), .A1 (outFilter1[329]), .S0 (
          nx8902)) ;
    ao22 ix935 (.Y (FilterToAlu_330), .A0 (outFilter0[330]), .A1 (nx8674), .B0 (
         outFilter1[330]), .B1 (nx8784)) ;
    ao22 ix941 (.Y (FilterToAlu_331), .A0 (outFilter0[331]), .A1 (nx8674), .B0 (
         outFilter1[331]), .B1 (nx8784)) ;
    ao22 ix947 (.Y (FilterToAlu_332), .A0 (outFilter0[332]), .A1 (nx8674), .B0 (
         outFilter1[332]), .B1 (nx8784)) ;
    ao22 ix953 (.Y (FilterToAlu_333), .A0 (outFilter0[333]), .A1 (nx8674), .B0 (
         outFilter1[333]), .B1 (nx8784)) ;
    ao22 ix959 (.Y (FilterToAlu_334), .A0 (outFilter0[334]), .A1 (nx8674), .B0 (
         outFilter1[334]), .B1 (nx8784)) ;
    ao22 ix965 (.Y (FilterToAlu_335), .A0 (outFilter0[335]), .A1 (nx8674), .B0 (
         outFilter1[335]), .B1 (nx8784)) ;
    ao22 ix791 (.Y (FilterToAlu_336), .A0 (outFilter0[336]), .A1 (nx8676), .B0 (
         outFilter1[336]), .B1 (nx8786)) ;
    ao22 ix797 (.Y (FilterToAlu_337), .A0 (outFilter0[337]), .A1 (nx8676), .B0 (
         outFilter1[337]), .B1 (nx8786)) ;
    ao22 ix803 (.Y (FilterToAlu_338), .A0 (outFilter0[338]), .A1 (nx8676), .B0 (
         outFilter1[338]), .B1 (nx8786)) ;
    ao22 ix809 (.Y (FilterToAlu_339), .A0 (outFilter0[339]), .A1 (nx8676), .B0 (
         outFilter1[339]), .B1 (nx8786)) ;
    ao22 ix815 (.Y (FilterToAlu_340), .A0 (outFilter0[340]), .A1 (nx8676), .B0 (
         outFilter1[340]), .B1 (nx8786)) ;
    ao22 ix821 (.Y (FilterToAlu_341), .A0 (outFilter0[341]), .A1 (nx8676), .B0 (
         outFilter1[341]), .B1 (nx8786)) ;
    ao22 ix827 (.Y (FilterToAlu_342), .A0 (outFilter0[342]), .A1 (nx8676), .B0 (
         outFilter1[342]), .B1 (nx8786)) ;
    ao22 ix833 (.Y (FilterToAlu_343), .A0 (outFilter0[343]), .A1 (nx8678), .B0 (
         outFilter1[343]), .B1 (nx8788)) ;
    ao22 ix839 (.Y (FilterToAlu_344), .A0 (outFilter0[344]), .A1 (nx8678), .B0 (
         outFilter1[344]), .B1 (nx8788)) ;
    nand02 ix295 (.Y (FilterToAlu_345), .A0 (nx8432), .A1 (nx8810)) ;
    mux21 ix8433 (.Y (nx8432), .A0 (outFilter0[345]), .A1 (outFilter1[345]), .S0 (
          nx8902)) ;
    ao22 ix845 (.Y (FilterToAlu_346), .A0 (outFilter0[346]), .A1 (nx8678), .B0 (
         outFilter1[346]), .B1 (nx8788)) ;
    ao22 ix851 (.Y (FilterToAlu_347), .A0 (outFilter0[347]), .A1 (nx8678), .B0 (
         outFilter1[347]), .B1 (nx8788)) ;
    ao22 ix857 (.Y (FilterToAlu_348), .A0 (outFilter0[348]), .A1 (nx8678), .B0 (
         outFilter1[348]), .B1 (nx8788)) ;
    ao22 ix863 (.Y (FilterToAlu_349), .A0 (outFilter0[349]), .A1 (nx8678), .B0 (
         outFilter1[349]), .B1 (nx8788)) ;
    ao22 ix869 (.Y (FilterToAlu_350), .A0 (outFilter0[350]), .A1 (nx8678), .B0 (
         outFilter1[350]), .B1 (nx8788)) ;
    ao22 ix875 (.Y (FilterToAlu_351), .A0 (outFilter0[351]), .A1 (nx8680), .B0 (
         outFilter1[351]), .B1 (nx8790)) ;
    ao22 ix701 (.Y (FilterToAlu_352), .A0 (outFilter0[352]), .A1 (nx8680), .B0 (
         outFilter1[352]), .B1 (nx8790)) ;
    ao22 ix707 (.Y (FilterToAlu_353), .A0 (outFilter0[353]), .A1 (nx8680), .B0 (
         outFilter1[353]), .B1 (nx8790)) ;
    ao22 ix713 (.Y (FilterToAlu_354), .A0 (outFilter0[354]), .A1 (nx8680), .B0 (
         outFilter1[354]), .B1 (nx8790)) ;
    ao22 ix719 (.Y (FilterToAlu_355), .A0 (outFilter0[355]), .A1 (nx8680), .B0 (
         outFilter1[355]), .B1 (nx8790)) ;
    ao22 ix725 (.Y (FilterToAlu_356), .A0 (outFilter0[356]), .A1 (nx8680), .B0 (
         outFilter1[356]), .B1 (nx8790)) ;
    ao22 ix731 (.Y (FilterToAlu_357), .A0 (outFilter0[357]), .A1 (nx8680), .B0 (
         outFilter1[357]), .B1 (nx8790)) ;
    ao22 ix737 (.Y (FilterToAlu_358), .A0 (outFilter0[358]), .A1 (nx8682), .B0 (
         outFilter1[358]), .B1 (nx8792)) ;
    ao22 ix743 (.Y (FilterToAlu_359), .A0 (outFilter0[359]), .A1 (nx8682), .B0 (
         outFilter1[359]), .B1 (nx8792)) ;
    ao22 ix749 (.Y (FilterToAlu_360), .A0 (outFilter0[360]), .A1 (nx8682), .B0 (
         outFilter1[360]), .B1 (nx8792)) ;
    nand02 ix285 (.Y (FilterToAlu_361), .A0 (nx8450), .A1 (nx8810)) ;
    mux21 ix8451 (.Y (nx8450), .A0 (outFilter0[361]), .A1 (outFilter1[361]), .S0 (
          nx8902)) ;
    ao22 ix755 (.Y (FilterToAlu_362), .A0 (outFilter0[362]), .A1 (nx8682), .B0 (
         outFilter1[362]), .B1 (nx8792)) ;
    ao22 ix761 (.Y (FilterToAlu_363), .A0 (outFilter0[363]), .A1 (nx8682), .B0 (
         outFilter1[363]), .B1 (nx8792)) ;
    ao22 ix767 (.Y (FilterToAlu_364), .A0 (outFilter0[364]), .A1 (nx8682), .B0 (
         outFilter1[364]), .B1 (nx8792)) ;
    ao22 ix773 (.Y (FilterToAlu_365), .A0 (outFilter0[365]), .A1 (nx8682), .B0 (
         outFilter1[365]), .B1 (nx8792)) ;
    ao22 ix779 (.Y (FilterToAlu_366), .A0 (outFilter0[366]), .A1 (nx8684), .B0 (
         outFilter1[366]), .B1 (nx8794)) ;
    ao22 ix785 (.Y (FilterToAlu_367), .A0 (outFilter0[367]), .A1 (nx8684), .B0 (
         outFilter1[367]), .B1 (nx8794)) ;
    ao22 ix611 (.Y (FilterToAlu_368), .A0 (outFilter0[368]), .A1 (nx8684), .B0 (
         outFilter1[368]), .B1 (nx8794)) ;
    ao22 ix617 (.Y (FilterToAlu_369), .A0 (outFilter0[369]), .A1 (nx8684), .B0 (
         outFilter1[369]), .B1 (nx8794)) ;
    ao22 ix623 (.Y (FilterToAlu_370), .A0 (outFilter0[370]), .A1 (nx8684), .B0 (
         outFilter1[370]), .B1 (nx8794)) ;
    ao22 ix629 (.Y (FilterToAlu_371), .A0 (outFilter0[371]), .A1 (nx8684), .B0 (
         outFilter1[371]), .B1 (nx8794)) ;
    ao22 ix635 (.Y (FilterToAlu_372), .A0 (outFilter0[372]), .A1 (nx8684), .B0 (
         outFilter1[372]), .B1 (nx8794)) ;
    ao22 ix641 (.Y (FilterToAlu_373), .A0 (outFilter0[373]), .A1 (nx8686), .B0 (
         outFilter1[373]), .B1 (nx8796)) ;
    ao22 ix647 (.Y (FilterToAlu_374), .A0 (outFilter0[374]), .A1 (nx8686), .B0 (
         outFilter1[374]), .B1 (nx8796)) ;
    ao22 ix653 (.Y (FilterToAlu_375), .A0 (outFilter0[375]), .A1 (nx8686), .B0 (
         outFilter1[375]), .B1 (nx8796)) ;
    ao22 ix659 (.Y (FilterToAlu_376), .A0 (outFilter0[376]), .A1 (nx8686), .B0 (
         outFilter1[376]), .B1 (nx8796)) ;
    nand02 ix275 (.Y (FilterToAlu_377), .A0 (nx8468), .A1 (nx8810)) ;
    mux21 ix8469 (.Y (nx8468), .A0 (outFilter0[377]), .A1 (outFilter1[377]), .S0 (
          nx8902)) ;
    ao22 ix665 (.Y (FilterToAlu_378), .A0 (outFilter0[378]), .A1 (nx8686), .B0 (
         outFilter1[378]), .B1 (nx8796)) ;
    ao22 ix671 (.Y (FilterToAlu_379), .A0 (outFilter0[379]), .A1 (nx8686), .B0 (
         outFilter1[379]), .B1 (nx8796)) ;
    ao22 ix677 (.Y (FilterToAlu_380), .A0 (outFilter0[380]), .A1 (nx8686), .B0 (
         outFilter1[380]), .B1 (nx8796)) ;
    ao22 ix683 (.Y (FilterToAlu_381), .A0 (outFilter0[381]), .A1 (nx8688), .B0 (
         outFilter1[381]), .B1 (nx8798)) ;
    ao22 ix689 (.Y (FilterToAlu_382), .A0 (outFilter0[382]), .A1 (nx8688), .B0 (
         outFilter1[382]), .B1 (nx8798)) ;
    ao22 ix695 (.Y (FilterToAlu_383), .A0 (outFilter0[383]), .A1 (nx8688), .B0 (
         outFilter1[383]), .B1 (nx8798)) ;
    ao22 ix521 (.Y (FilterToAlu_384), .A0 (outFilter0[384]), .A1 (nx8688), .B0 (
         outFilter1[384]), .B1 (nx8798)) ;
    ao22 ix527 (.Y (FilterToAlu_385), .A0 (outFilter0[385]), .A1 (nx8688), .B0 (
         outFilter1[385]), .B1 (nx8798)) ;
    ao22 ix533 (.Y (FilterToAlu_386), .A0 (outFilter0[386]), .A1 (nx8688), .B0 (
         outFilter1[386]), .B1 (nx8798)) ;
    ao22 ix539 (.Y (FilterToAlu_387), .A0 (outFilter0[387]), .A1 (nx8688), .B0 (
         outFilter1[387]), .B1 (nx8798)) ;
    ao22 ix545 (.Y (FilterToAlu_388), .A0 (outFilter0[388]), .A1 (nx8690), .B0 (
         outFilter1[388]), .B1 (nx8800)) ;
    ao22 ix551 (.Y (FilterToAlu_389), .A0 (outFilter0[389]), .A1 (nx8690), .B0 (
         outFilter1[389]), .B1 (nx8800)) ;
    ao22 ix557 (.Y (FilterToAlu_390), .A0 (outFilter0[390]), .A1 (nx8690), .B0 (
         outFilter1[390]), .B1 (nx8800)) ;
    ao22 ix563 (.Y (FilterToAlu_391), .A0 (outFilter0[391]), .A1 (nx8690), .B0 (
         outFilter1[391]), .B1 (nx8800)) ;
    ao22 ix569 (.Y (FilterToAlu_392), .A0 (outFilter0[392]), .A1 (nx8690), .B0 (
         outFilter1[392]), .B1 (nx8800)) ;
    nand02 ix265 (.Y (FilterToAlu_393), .A0 (nx8486), .A1 (nx8810)) ;
    mux21 ix8487 (.Y (nx8486), .A0 (outFilter0[393]), .A1 (outFilter1[393]), .S0 (
          nx8902)) ;
    ao22 ix575 (.Y (FilterToAlu_394), .A0 (outFilter0[394]), .A1 (nx8690), .B0 (
         outFilter1[394]), .B1 (nx8800)) ;
    ao22 ix581 (.Y (FilterToAlu_395), .A0 (outFilter0[395]), .A1 (nx8690), .B0 (
         outFilter1[395]), .B1 (nx8800)) ;
    ao22 ix587 (.Y (FilterToAlu_396), .A0 (outFilter0[396]), .A1 (nx8692), .B0 (
         outFilter1[396]), .B1 (nx8802)) ;
    ao22 ix593 (.Y (FilterToAlu_397), .A0 (outFilter0[397]), .A1 (nx8692), .B0 (
         outFilter1[397]), .B1 (nx8802)) ;
    ao22 ix599 (.Y (FilterToAlu_398), .A0 (outFilter0[398]), .A1 (nx8692), .B0 (
         outFilter1[398]), .B1 (nx8802)) ;
    ao22 ix605 (.Y (FilterToAlu_399), .A0 (outFilter0[399]), .A1 (nx8692), .B0 (
         outFilter1[399]), .B1 (nx8802)) ;
    nand02 ix55 (.Y (ConvOuput[0]), .A0 (nx8495), .A1 (nx8501)) ;
    aoi32 ix8496 (.Y (nx8495), .A0 (nx8916), .A1 (AddOut33_3), .A2 (nx8852), .B0 (
          nx32), .B1 (nx34)) ;
    mux21_ni ix33 (.Y (nx32), .A0 (AddOut33_5), .A1 (Final55_5), .S0 (nx8884)) ;
    aoi32 ix8502 (.Y (nx8501), .A0 (Final55_0), .A1 (nx8884), .A2 (nx8904), .B0 (
          AddOut33_0), .B1 (nx20)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (nx8852), .A1 (nx6)) ;
    mux21_ni ix7 (.Y (nx6), .A0 (AddOut33_15), .A1 (Final55_15), .S0 (nx8886)) ;
    nand02 ix85 (.Y (ConvOuput[1]), .A0 (nx8511), .A1 (nx8514)) ;
    aoi32 ix8512 (.Y (nx8511), .A0 (nx8916), .A1 (AddOut33_4), .A2 (nx8852), .B0 (
          nx68), .B1 (nx34)) ;
    mux21_ni ix69 (.Y (nx68), .A0 (AddOut33_6), .A1 (Final55_6), .S0 (nx8886)) ;
    aoi32 ix8515 (.Y (nx8514), .A0 (Final55_1), .A1 (nx8886), .A2 (nx8904), .B0 (
          AddOut33_1), .B1 (nx20)) ;
    nand02 ix107 (.Y (ConvOuput[2]), .A0 (nx8517), .A1 (nx8520)) ;
    aoi32 ix8518 (.Y (nx8517), .A0 (Final55_7), .A1 (nx8886), .A2 (nx8852), .B0 (
          nx32), .B1 (nx8908)) ;
    aoi32 ix8521 (.Y (nx8520), .A0 (Final55_2), .A1 (nx8886), .A2 (nx8904), .B0 (
          AddOut33_2), .B1 (nx20)) ;
    oai21 ix125 (.Y (ConvOuput[3]), .A0 (nx8523), .A1 (nx8812), .B0 (nx8525)) ;
    mux21 ix8524 (.Y (nx8523), .A0 (AddOut33_3), .A1 (Final55_3), .S0 (nx8886)
          ) ;
    aoi32 ix8526 (.Y (nx8525), .A0 (Final55_8), .A1 (nx8886), .A2 (nx8852), .B0 (
          nx68), .B1 (nx8908)) ;
    oai21 ix143 (.Y (ConvOuput[4]), .A0 (nx8528), .A1 (nx8812), .B0 (nx8530)) ;
    mux21 ix8529 (.Y (nx8528), .A0 (AddOut33_4), .A1 (Final55_4), .S0 (nx8888)
          ) ;
    aoi32 ix8531 (.Y (nx8530), .A0 (Final55_9), .A1 (nx8888), .A2 (nx8852), .B0 (
          nx98), .B1 (nx8908)) ;
    mux21_ni ix99 (.Y (nx98), .A0 (AddOut33_7), .A1 (Final55_7), .S0 (nx8888)) ;
    oai21 ix161 (.Y (ConvOuput[5]), .A0 (nx8534), .A1 (nx8812), .B0 (nx8536)) ;
    aoi32 ix8537 (.Y (nx8536), .A0 (Final55_10), .A1 (nx8888), .A2 (nx8854), .B0 (
          nx116), .B1 (nx8908)) ;
    mux21_ni ix117 (.Y (nx116), .A0 (AddOut33_8), .A1 (Final55_8), .S0 (nx8888)
             ) ;
    oai21 ix179 (.Y (ConvOuput[6]), .A0 (nx8540), .A1 (nx8812), .B0 (nx8542)) ;
    aoi32 ix8543 (.Y (nx8542), .A0 (Final55_11), .A1 (nx8888), .A2 (nx8854), .B0 (
          nx134), .B1 (nx8908)) ;
    mux21_ni ix135 (.Y (nx134), .A0 (AddOut33_9), .A1 (Final55_9), .S0 (nx8888)
             ) ;
    oai21 ix197 (.Y (ConvOuput[7]), .A0 (nx8546), .A1 (nx8812), .B0 (nx8548)) ;
    aoi32 ix8549 (.Y (nx8548), .A0 (Final55_12), .A1 (nx8890), .A2 (nx8854), .B0 (
          nx152), .B1 (nx8908)) ;
    mux21_ni ix153 (.Y (nx152), .A0 (AddOut33_10), .A1 (Final55_10), .S0 (nx8890
             )) ;
    oai21 ix215 (.Y (ConvOuput[8]), .A0 (nx8552), .A1 (nx8812), .B0 (nx8554)) ;
    aoi32 ix8555 (.Y (nx8554), .A0 (Final55_13), .A1 (nx8890), .A2 (nx8854), .B0 (
          nx170), .B1 (nx8908)) ;
    mux21_ni ix171 (.Y (nx170), .A0 (AddOut33_11), .A1 (Final55_11), .S0 (nx8890
             )) ;
    oai21 ix233 (.Y (ConvOuput[9]), .A0 (nx8558), .A1 (nx8814), .B0 (nx8560)) ;
    aoi32 ix8561 (.Y (nx8560), .A0 (Final55_14), .A1 (nx8890), .A2 (nx8854), .B0 (
          nx188), .B1 (nx8910)) ;
    mux21_ni ix189 (.Y (nx188), .A0 (AddOut33_12), .A1 (Final55_12), .S0 (nx8890
             )) ;
    oai21 ix243 (.Y (ConvOuput[10]), .A0 (nx8564), .A1 (nx8814), .B0 (nx8566)) ;
    aoi32 ix8567 (.Y (nx8566), .A0 (nx8916), .A1 (AddOut33_13), .A2 (nx8854), .B0 (
          nx6), .B1 (nx34)) ;
    oai21 ix253 (.Y (ConvOuput[11]), .A0 (nx8569), .A1 (nx8814), .B0 (nx8571)) ;
    aoi32 ix8572 (.Y (nx8571), .A0 (nx8916), .A1 (AddOut33_14), .A2 (nx8854), .B0 (
          nx6), .B1 (nx34)) ;
    ao21 ix2769 (.Y (ConvOuput[12]), .A0 (nx188), .A1 (nx8904), .B0 (
         ConvOuput[15])) ;
    ao21 ix2773 (.Y (ConvOuput[13]), .A0 (nx206), .A1 (nx8904), .B0 (
         ConvOuput[15])) ;
    mux21_ni ix207 (.Y (nx206), .A0 (AddOut33_13), .A1 (Final55_13), .S0 (nx8890
             )) ;
    ao21 ix2777 (.Y (ConvOuput[14]), .A0 (nx224), .A1 (nx8904), .B0 (
         ConvOuput[15])) ;
    mux21_ni ix225 (.Y (nx224), .A0 (AddOut33_14), .A1 (Final55_14), .S0 (nx8892
             )) ;
    inv01 ix8570 (.Y (nx8569), .A (nx170)) ;
    inv01 ix8565 (.Y (nx8564), .A (nx152)) ;
    inv01 ix8559 (.Y (nx8558), .A (nx134)) ;
    inv01 ix8553 (.Y (nx8552), .A (nx116)) ;
    inv01 ix8547 (.Y (nx8546), .A (nx98)) ;
    inv01 ix8541 (.Y (nx8540), .A (nx68)) ;
    inv01 ix8535 (.Y (nx8534), .A (nx32)) ;
    inv02 ix8585 (.Y (nx8586), .A (nx8816)) ;
    inv02 ix8587 (.Y (nx8588), .A (nx8816)) ;
    inv02 ix8589 (.Y (nx8590), .A (nx8816)) ;
    inv02 ix8591 (.Y (nx8592), .A (nx8816)) ;
    inv02 ix8593 (.Y (nx8594), .A (nx8816)) ;
    inv02 ix8595 (.Y (nx8596), .A (nx8816)) ;
    inv02 ix8597 (.Y (nx8598), .A (nx8816)) ;
    inv02 ix8599 (.Y (nx8600), .A (nx8818)) ;
    inv02 ix8601 (.Y (nx8602), .A (nx8818)) ;
    inv02 ix8603 (.Y (nx8604), .A (nx8818)) ;
    inv02 ix8605 (.Y (nx8606), .A (nx8818)) ;
    inv02 ix8607 (.Y (nx8608), .A (nx8818)) ;
    inv02 ix8609 (.Y (nx8610), .A (nx8818)) ;
    inv02 ix8611 (.Y (nx8612), .A (nx8818)) ;
    inv02 ix8613 (.Y (nx8614), .A (nx8820)) ;
    inv02 ix8615 (.Y (nx8616), .A (nx8820)) ;
    inv02 ix8617 (.Y (nx8618), .A (nx8820)) ;
    inv02 ix8619 (.Y (nx8620), .A (nx8820)) ;
    inv02 ix8621 (.Y (nx8622), .A (nx8820)) ;
    inv02 ix8623 (.Y (nx8624), .A (nx8820)) ;
    inv02 ix8625 (.Y (nx8626), .A (nx8820)) ;
    inv02 ix8627 (.Y (nx8628), .A (nx8822)) ;
    inv02 ix8629 (.Y (nx8630), .A (nx8822)) ;
    inv02 ix8631 (.Y (nx8632), .A (nx8822)) ;
    inv02 ix8633 (.Y (nx8634), .A (nx8822)) ;
    inv02 ix8635 (.Y (nx8636), .A (nx8822)) ;
    inv02 ix8637 (.Y (nx8638), .A (nx8822)) ;
    inv02 ix8639 (.Y (nx8640), .A (nx8822)) ;
    inv02 ix8641 (.Y (nx8642), .A (nx8824)) ;
    inv02 ix8643 (.Y (nx8644), .A (nx8824)) ;
    inv02 ix8645 (.Y (nx8646), .A (nx8824)) ;
    inv02 ix8647 (.Y (nx8648), .A (nx8824)) ;
    inv02 ix8649 (.Y (nx8650), .A (nx8824)) ;
    inv02 ix8651 (.Y (nx8652), .A (nx8824)) ;
    inv02 ix8653 (.Y (nx8654), .A (nx8824)) ;
    inv02 ix8655 (.Y (nx8656), .A (nx8826)) ;
    inv02 ix8657 (.Y (nx8658), .A (nx8826)) ;
    inv02 ix8659 (.Y (nx8660), .A (nx8826)) ;
    inv02 ix8661 (.Y (nx8662), .A (nx8826)) ;
    inv02 ix8663 (.Y (nx8664), .A (nx8826)) ;
    inv02 ix8665 (.Y (nx8666), .A (nx8826)) ;
    inv02 ix8667 (.Y (nx8668), .A (nx8826)) ;
    inv02 ix8669 (.Y (nx8670), .A (nx8828)) ;
    inv02 ix8671 (.Y (nx8672), .A (nx8828)) ;
    inv02 ix8673 (.Y (nx8674), .A (nx8828)) ;
    inv02 ix8675 (.Y (nx8676), .A (nx8828)) ;
    inv02 ix8677 (.Y (nx8678), .A (nx8828)) ;
    inv02 ix8679 (.Y (nx8680), .A (nx8828)) ;
    inv02 ix8681 (.Y (nx8682), .A (nx8828)) ;
    inv02 ix8683 (.Y (nx8684), .A (nx8830)) ;
    inv02 ix8685 (.Y (nx8686), .A (nx8830)) ;
    inv02 ix8687 (.Y (nx8688), .A (nx8830)) ;
    inv02 ix8689 (.Y (nx8690), .A (nx8830)) ;
    inv02 ix8691 (.Y (nx8692), .A (nx8830)) ;
    inv02 ix8695 (.Y (nx8696), .A (nx8926)) ;
    inv02 ix8697 (.Y (nx8698), .A (nx8926)) ;
    inv02 ix8699 (.Y (nx8700), .A (nx8926)) ;
    inv02 ix8701 (.Y (nx8702), .A (nx8926)) ;
    inv02 ix8703 (.Y (nx8704), .A (nx8926)) ;
    inv02 ix8705 (.Y (nx8706), .A (nx8926)) ;
    inv02 ix8707 (.Y (nx8708), .A (nx8832)) ;
    inv02 ix8709 (.Y (nx8710), .A (nx8834)) ;
    inv02 ix8711 (.Y (nx8712), .A (nx8834)) ;
    inv02 ix8713 (.Y (nx8714), .A (nx8834)) ;
    inv02 ix8715 (.Y (nx8716), .A (nx8834)) ;
    inv02 ix8717 (.Y (nx8718), .A (nx8834)) ;
    inv02 ix8719 (.Y (nx8720), .A (nx8834)) ;
    inv02 ix8721 (.Y (nx8722), .A (nx8834)) ;
    inv02 ix8723 (.Y (nx8724), .A (nx8836)) ;
    inv02 ix8725 (.Y (nx8726), .A (nx8836)) ;
    inv02 ix8727 (.Y (nx8728), .A (nx8836)) ;
    inv02 ix8729 (.Y (nx8730), .A (nx8836)) ;
    inv02 ix8731 (.Y (nx8732), .A (nx8836)) ;
    inv02 ix8733 (.Y (nx8734), .A (nx8836)) ;
    inv02 ix8735 (.Y (nx8736), .A (nx8836)) ;
    inv02 ix8737 (.Y (nx8738), .A (nx8838)) ;
    inv02 ix8739 (.Y (nx8740), .A (nx8838)) ;
    inv02 ix8741 (.Y (nx8742), .A (nx8838)) ;
    inv02 ix8743 (.Y (nx8744), .A (nx8838)) ;
    inv02 ix8745 (.Y (nx8746), .A (nx8838)) ;
    inv02 ix8747 (.Y (nx8748), .A (nx8838)) ;
    inv02 ix8749 (.Y (nx8750), .A (nx8838)) ;
    inv02 ix8751 (.Y (nx8752), .A (nx8840)) ;
    inv02 ix8753 (.Y (nx8754), .A (nx8840)) ;
    inv02 ix8755 (.Y (nx8756), .A (nx8840)) ;
    inv02 ix8757 (.Y (nx8758), .A (nx8840)) ;
    inv02 ix8759 (.Y (nx8760), .A (nx8840)) ;
    inv02 ix8761 (.Y (nx8762), .A (nx8840)) ;
    inv02 ix8763 (.Y (nx8764), .A (nx8840)) ;
    inv02 ix8765 (.Y (nx8766), .A (nx8842)) ;
    inv02 ix8767 (.Y (nx8768), .A (nx8842)) ;
    inv02 ix8769 (.Y (nx8770), .A (nx8842)) ;
    inv02 ix8771 (.Y (nx8772), .A (nx8842)) ;
    inv02 ix8773 (.Y (nx8774), .A (nx8842)) ;
    inv02 ix8775 (.Y (nx8776), .A (nx8842)) ;
    inv02 ix8777 (.Y (nx8778), .A (nx8842)) ;
    inv02 ix8779 (.Y (nx8780), .A (nx8844)) ;
    inv02 ix8781 (.Y (nx8782), .A (nx8844)) ;
    inv02 ix8783 (.Y (nx8784), .A (nx8844)) ;
    inv02 ix8785 (.Y (nx8786), .A (nx8844)) ;
    inv02 ix8787 (.Y (nx8788), .A (nx8844)) ;
    inv02 ix8789 (.Y (nx8790), .A (nx8844)) ;
    inv02 ix8791 (.Y (nx8792), .A (nx8844)) ;
    inv02 ix8793 (.Y (nx8794), .A (nx8846)) ;
    inv02 ix8795 (.Y (nx8796), .A (nx8846)) ;
    inv02 ix8797 (.Y (nx8798), .A (nx8846)) ;
    inv02 ix8799 (.Y (nx8800), .A (nx8846)) ;
    inv02 ix8801 (.Y (nx8802), .A (nx8846)) ;
    inv02 ix8803 (.Y (nx8804), .A (LayerInfo[15])) ;
    inv02 ix8805 (.Y (nx8806), .A (nx8856)) ;
    inv02 ix8807 (.Y (nx8808), .A (nx8856)) ;
    inv02 ix8809 (.Y (nx8810), .A (nx8856)) ;
    inv02 ix8811 (.Y (nx8812), .A (nx12)) ;
    inv02 ix8813 (.Y (nx8814), .A (nx8904)) ;
    inv02 ix8815 (.Y (nx8816), .A (nx510)) ;
    inv02 ix8817 (.Y (nx8818), .A (nx510)) ;
    inv02 ix8819 (.Y (nx8820), .A (nx510)) ;
    inv02 ix8821 (.Y (nx8822), .A (nx510)) ;
    inv02 ix8823 (.Y (nx8824), .A (nx510)) ;
    inv02 ix8825 (.Y (nx8826), .A (nx510)) ;
    inv02 ix8827 (.Y (nx8828), .A (nx510)) ;
    inv02 ix8829 (.Y (nx8830), .A (nx510)) ;
    inv02 ix8831 (.Y (nx8832), .A (nx516)) ;
    inv02 ix8833 (.Y (nx8834), .A (nx8912)) ;
    inv02 ix8835 (.Y (nx8836), .A (nx8912)) ;
    inv02 ix8837 (.Y (nx8838), .A (nx8912)) ;
    inv02 ix8839 (.Y (nx8840), .A (nx8912)) ;
    inv02 ix8841 (.Y (nx8842), .A (nx8912)) ;
    inv02 ix8843 (.Y (nx8844), .A (nx8914)) ;
    inv02 ix8845 (.Y (nx8846), .A (nx8914)) ;
    nor02ii ix517 (.Y (nx516), .A0 (nx8856), .A1 (nx8902)) ;
    and02 ix35 (.Y (nx34), .A0 (nx8892), .A1 (nx8856)) ;
    nor02ii ix21 (.Y (nx20), .A0 (nx8892), .A1 (nx8906)) ;
    nor02ii ix49 (.Y (nx48), .A0 (nx8892), .A1 (nx8856)) ;
    and02 ix255 (.Y (ConvOuput[15]), .A0 (nx8856), .A1 (nx6)) ;
    inv02 ix8851 (.Y (nx8852), .A (nx8804)) ;
    inv02 ix8853 (.Y (nx8854), .A (nx8804)) ;
    inv02 ix8855 (.Y (nx8856), .A (nx8804)) ;
    inv02 ix8857 (.Y (nx8858), .A (nx8916)) ;
    inv02 ix8859 (.Y (nx8860), .A (nx8916)) ;
    inv02 ix8861 (.Y (nx8862), .A (nx8916)) ;
    inv02 ix8863 (.Y (nx8864), .A (nx8918)) ;
    inv02 ix8865 (.Y (nx8866), .A (nx8918)) ;
    inv02 ix8867 (.Y (nx8868), .A (nx8918)) ;
    inv02 ix8869 (.Y (nx8870), .A (nx8918)) ;
    inv02 ix8871 (.Y (nx8872), .A (nx8918)) ;
    inv02 ix8873 (.Y (nx8874), .A (nx8918)) ;
    inv02 ix8875 (.Y (nx8876), .A (nx8918)) ;
    inv02 ix8877 (.Y (nx8878), .A (nx8920)) ;
    inv02 ix8879 (.Y (nx8880), .A (nx8920)) ;
    inv02 ix8881 (.Y (nx8882), .A (nx8920)) ;
    inv02 ix8883 (.Y (nx8884), .A (nx8920)) ;
    inv02 ix8885 (.Y (nx8886), .A (nx8920)) ;
    inv02 ix8887 (.Y (nx8888), .A (nx8920)) ;
    inv02 ix8889 (.Y (nx8890), .A (nx8920)) ;
    inv02 ix8891 (.Y (nx8892), .A (nx8922)) ;
    inv01 ix8893 (.Y (nx8894), .A (QImgStat)) ;
    inv02 ix8895 (.Y (nx8896), .A (nx8894)) ;
    inv02 ix8897 (.Y (nx8898), .A (nx8894)) ;
    inv02 ix8899 (.Y (nx8900), .A (nx8894)) ;
    inv02 ix8901 (.Y (nx8902), .A (nx8894)) ;
    inv02 ix8903 (.Y (nx8904), .A (nx8812)) ;
    inv02 ix8905 (.Y (nx8906), .A (nx8812)) ;
    buf02 ix8907 (.Y (nx8908), .A (nx48)) ;
    buf02 ix8909 (.Y (nx8910), .A (nx48)) ;
    inv01 ix8911 (.Y (nx8912), .A (nx8926)) ;
    inv01 ix8913 (.Y (nx8914), .A (nx8832)) ;
    inv02 ix8915 (.Y (nx8916), .A (LayerInfo[14])) ;
    inv02 ix8917 (.Y (nx8918), .A (LayerInfo[14])) ;
    inv02 ix8919 (.Y (nx8920), .A (LayerInfo[14])) ;
    inv02 ix8921 (.Y (nx8922), .A (LayerInfo[14])) ;
    inv02 ix8923 (.Y (nx8924), .A (LayerInfo[15])) ;
    inv02 ix8925 (.Y (nx8926), .A (nx516)) ;
endmodule


module Multiplier_16 ( A, B, F ) ;

    input [15:0]A ;
    input [15:0]B ;
    output [31:0]F ;

    wire addout_0__31, addout_0__30, addout_0__29, addout_0__28, addout_0__27, 
         addout_0__26, addout_0__25, addout_0__24, addout_0__23, addout_0__22, 
         addout_0__21, addout_0__20, addout_0__19, addout_0__18, addout_0__17, 
         addout_0__16, addout_0__15, addout_0__14, addout_0__13, addout_0__12, 
         addout_0__11, addout_0__10, addout_0__9, addout_0__8, addout_0__7, 
         addout_0__6, addout_0__5, addout_0__4, addout_0__3, addout_0__2, 
         addout_0__1, addout_0__0, addout_1__31, addout_1__30, addout_1__29, 
         addout_1__28, addout_1__27, addout_1__26, addout_1__25, addout_1__24, 
         addout_1__23, addout_1__22, addout_1__21, addout_1__20, addout_1__19, 
         addout_1__18, addout_1__17, addout_1__16, addout_1__15, addout_1__14, 
         addout_1__13, addout_1__12, addout_1__11, addout_1__10, addout_1__9, 
         addout_1__8, addout_1__7, addout_1__6, addout_1__5, addout_1__4, 
         addout_1__3, addout_1__2, addout_1__1, addout_1__0, addout_2__31, 
         addout_2__30, addout_2__29, addout_2__28, addout_2__27, addout_2__26, 
         addout_2__25, addout_2__24, addout_2__23, addout_2__22, addout_2__21, 
         addout_2__20, addout_2__19, addout_2__18, addout_2__17, addout_2__16, 
         addout_2__15, addout_2__14, addout_2__13, addout_2__12, addout_2__11, 
         addout_2__10, addout_2__9, addout_2__8, addout_2__7, addout_2__6, 
         addout_2__5, addout_2__4, addout_2__3, addout_2__2, addout_2__1, 
         addout_2__0, addout_3__31, addout_3__30, addout_3__29, addout_3__28, 
         addout_3__27, addout_3__26, addout_3__25, addout_3__24, addout_3__23, 
         addout_3__22, addout_3__21, addout_3__20, addout_3__19, addout_3__18, 
         addout_3__17, addout_3__16, addout_3__15, addout_3__14, addout_3__13, 
         addout_3__12, addout_3__11, addout_3__10, addout_3__9, addout_3__8, 
         addout_3__7, addout_3__6, addout_3__5, addout_3__4, addout_3__3, 
         addout_3__2, addout_3__1, addout_3__0, addout_4__31, addout_4__30, 
         addout_4__29, addout_4__28, addout_4__27, addout_4__26, addout_4__25, 
         addout_4__24, addout_4__23, addout_4__22, addout_4__21, addout_4__20, 
         addout_4__19, addout_4__18, addout_4__17, addout_4__16, addout_4__15, 
         addout_4__14, addout_4__13, addout_4__12, addout_4__11, addout_4__10, 
         addout_4__9, addout_4__8, addout_4__7, addout_4__6, addout_4__5, 
         addout_4__4, addout_4__3, addout_4__2, addout_4__1, addout_4__0, 
         addout_5__31, addout_5__30, addout_5__29, addout_5__28, addout_5__27, 
         addout_5__26, addout_5__25, addout_5__24, addout_5__23, addout_5__22, 
         addout_5__21, addout_5__20, addout_5__19, addout_5__18, addout_5__17, 
         addout_5__16, addout_5__15, addout_5__14, addout_5__13, addout_5__12, 
         addout_5__11, addout_5__10, addout_5__9, addout_5__8, addout_5__7, 
         addout_5__6, addout_5__5, addout_5__4, addout_5__3, addout_5__2, 
         addout_5__1, addout_5__0, addout_6__31, addout_6__30, addout_6__29, 
         addout_6__28, addout_6__27, addout_6__26, addout_6__25, addout_6__24, 
         addout_6__23, addout_6__22, addout_6__21, addout_6__20, addout_6__19, 
         addout_6__18, addout_6__17, addout_6__16, addout_6__15, addout_6__14, 
         addout_6__13, addout_6__12, addout_6__11, addout_6__10, addout_6__9, 
         addout_6__8, addout_6__7, addout_6__6, addout_6__5, addout_6__4, 
         addout_6__3, addout_6__2, addout_6__1, addout_6__0, addout_7__31, 
         addout_7__30, addout_7__29, addout_7__28, addout_7__27, addout_7__26, 
         addout_7__25, addout_7__24, addout_7__23, addout_7__22, addout_7__21, 
         addout_7__20, addout_7__19, addout_7__18, addout_7__17, addout_7__16, 
         addout_7__15, addout_7__14, addout_7__13, addout_7__12, addout_7__11, 
         addout_7__10, addout_7__9, addout_7__8, addout_7__7, addout_7__6, 
         addout_7__5, addout_7__4, addout_7__3, addout_7__2, addout_7__1, 
         addout_7__0, addout_8__31, addout_8__30, addout_8__29, addout_8__28, 
         addout_8__27, addout_8__26, addout_8__25, addout_8__24, addout_8__23, 
         addout_8__22, addout_8__21, addout_8__20, addout_8__19, addout_8__18, 
         addout_8__17, addout_8__16, addout_8__15, addout_8__14, addout_8__13, 
         addout_8__12, addout_8__11, addout_8__10, addout_8__9, addout_8__8, 
         addout_8__7, addout_8__6, addout_8__5, addout_8__4, addout_8__3, 
         addout_8__2, addout_8__1, addout_8__0, addout_9__31, addout_9__30, 
         addout_9__29, addout_9__28, addout_9__27, addout_9__26, addout_9__25, 
         addout_9__24, addout_9__23, addout_9__22, addout_9__21, addout_9__20, 
         addout_9__19, addout_9__18, addout_9__17, addout_9__16, addout_9__15, 
         addout_9__14, addout_9__13, addout_9__12, addout_9__11, addout_9__10, 
         addout_9__9, addout_9__8, addout_9__7, addout_9__6, addout_9__5, 
         addout_9__4, addout_9__3, addout_9__2, addout_9__1, addout_9__0, 
         addout_10__31, addout_10__30, addout_10__29, addout_10__28, 
         addout_10__27, addout_10__26, addout_10__25, addout_10__24, 
         addout_10__23, addout_10__22, addout_10__21, addout_10__20, 
         addout_10__19, addout_10__18, addout_10__17, addout_10__16, 
         addout_10__15, addout_10__14, addout_10__13, addout_10__12, 
         addout_10__11, addout_10__10, addout_10__9, addout_10__8, addout_10__7, 
         addout_10__6, addout_10__5, addout_10__4, addout_10__3, addout_10__2, 
         addout_10__1, addout_10__0, addout_11__31, addout_11__30, addout_11__29, 
         addout_11__28, addout_11__27, addout_11__26, addout_11__25, 
         addout_11__24, addout_11__23, addout_11__22, addout_11__21, 
         addout_11__20, addout_11__19, addout_11__18, addout_11__17, 
         addout_11__16, addout_11__15, addout_11__14, addout_11__13, 
         addout_11__12, addout_11__11, addout_11__10, addout_11__9, addout_11__8, 
         addout_11__7, addout_11__6, addout_11__5, addout_11__4, addout_11__3, 
         addout_11__2, addout_11__1, addout_11__0, addout_12__31, addout_12__30, 
         addout_12__29, addout_12__28, addout_12__27, addout_12__26, 
         addout_12__25, addout_12__24, addout_12__23, addout_12__22, 
         addout_12__21, addout_12__20, addout_12__19, addout_12__18, 
         addout_12__17, addout_12__16, addout_12__15, addout_12__14, 
         addout_12__13, addout_12__12, addout_12__11, addout_12__10, 
         addout_12__9, addout_12__8, addout_12__7, addout_12__6, addout_12__5, 
         addout_12__4, addout_12__3, addout_12__2, addout_12__1, addout_12__0, 
         addout_13__31, addout_13__30, addout_13__29, addout_13__28, 
         addout_13__27, addout_13__26, addout_13__25, addout_13__24, 
         addout_13__23, addout_13__22, addout_13__21, addout_13__20, 
         addout_13__19, addout_13__18, addout_13__17, addout_13__16, 
         addout_13__15, addout_13__14, addout_13__13, addout_13__12, 
         addout_13__11, addout_13__10, addout_13__9, addout_13__8, addout_13__7, 
         addout_13__6, addout_13__5, addout_13__4, addout_13__3, addout_13__2, 
         addout_13__1, addout_13__0, addout_14__31, addout_14__30, addout_14__29, 
         addout_14__28, addout_14__27, addout_14__26, addout_14__25, 
         addout_14__24, addout_14__23, addout_14__22, addout_14__21, 
         addout_14__20, addout_14__19, addout_14__18, addout_14__17, 
         addout_14__16, addout_14__15, addout_14__14, addout_14__13, 
         addout_14__12, addout_14__11, addout_14__10, addout_14__9, addout_14__8, 
         addout_14__7, addout_14__6, addout_14__5, addout_14__4, addout_14__3, 
         addout_14__2, addout_14__1, addout_14__0, addout_15__31, addout_15__30, 
         addout_15__29, addout_15__28, addout_15__27, addout_15__26, 
         addout_15__25, addout_15__24, addout_15__23, addout_15__22, 
         addout_15__21, addout_15__20, addout_15__19, addout_15__18, 
         addout_15__17, addout_15__16, addout_15__15, addout_15__14, 
         addout_15__13, addout_15__12, addout_15__11, addout_15__10, 
         addout_15__9, addout_15__8, addout_15__7, addout_15__6, addout_15__5, 
         addout_15__4, addout_15__3, addout_15__2, addout_15__1, addout_15__0, 
         addout_16__31, addout_16__30, addout_16__29, addout_16__28, 
         addout_16__27, addout_16__26, addout_16__25, addout_16__24, 
         addout_16__23, addout_16__22, addout_16__21, addout_16__20, 
         addout_16__19, addout_16__18, addout_16__17, addout_16__16, 
         addout_16__15, addout_16__14, addout_16__13, addout_16__12, 
         addout_16__11, addout_16__10, addout_16__9, addout_16__8, addout_16__7, 
         addout_16__6, addout_16__5, addout_16__4, addout_16__3, addout_16__2, 
         addout_16__1, addout_16__0, addout_17__31, addout_17__30, addout_17__29, 
         addout_17__28, addout_17__27, addout_17__26, addout_17__25, 
         addout_17__24, addout_17__23, addout_17__22, addout_17__21, 
         addout_17__20, addout_17__19, addout_17__18, addout_17__17, 
         addout_17__16, addout_17__15, addout_17__14, addout_17__13, 
         addout_17__12, addout_17__11, addout_17__10, addout_17__9, addout_17__8, 
         addout_17__7, addout_17__6, addout_17__5, addout_17__4, addout_17__3, 
         addout_17__2, addout_17__1, addout_17__0, addout_18__31, addout_18__30, 
         addout_18__29, addout_18__28, addout_18__27, addout_18__26, 
         addout_18__25, addout_18__24, addout_18__23, addout_18__22, 
         addout_18__21, addout_18__20, addout_18__19, addout_18__18, 
         addout_18__17, addout_18__16, addout_18__15, addout_18__14, 
         addout_18__13, addout_18__12, addout_18__11, addout_18__10, 
         addout_18__9, addout_18__8, addout_18__7, addout_18__6, addout_18__5, 
         addout_18__4, addout_18__3, addout_18__2, addout_18__1, addout_18__0, 
         addout_19__31, addout_19__30, addout_19__29, addout_19__28, 
         addout_19__27, addout_19__26, addout_19__25, addout_19__24, 
         addout_19__23, addout_19__22, addout_19__21, addout_19__20, 
         addout_19__19, addout_19__18, addout_19__17, addout_19__16, 
         addout_19__15, addout_19__14, addout_19__13, addout_19__12, 
         addout_19__11, addout_19__10, addout_19__9, addout_19__8, addout_19__7, 
         addout_19__6, addout_19__5, addout_19__4, addout_19__3, addout_19__2, 
         addout_19__1, addout_19__0, addout_20__31, addout_20__30, addout_20__29, 
         addout_20__28, addout_20__27, addout_20__26, addout_20__25, 
         addout_20__24, addout_20__23, addout_20__22, addout_20__21, 
         addout_20__20, addout_20__19, addout_20__18, addout_20__17, 
         addout_20__16, addout_20__15, addout_20__14, addout_20__13, 
         addout_20__12, addout_20__11, addout_20__10, addout_20__9, addout_20__8, 
         addout_20__7, addout_20__6, addout_20__5, addout_20__4, addout_20__3, 
         addout_20__2, addout_20__1, addout_20__0, addout_21__31, addout_21__30, 
         addout_21__29, addout_21__28, addout_21__27, addout_21__26, 
         addout_21__25, addout_21__24, addout_21__23, addout_21__22, 
         addout_21__21, addout_21__20, addout_21__19, addout_21__18, 
         addout_21__17, addout_21__16, addout_21__15, addout_21__14, 
         addout_21__13, addout_21__12, addout_21__11, addout_21__10, 
         addout_21__9, addout_21__8, addout_21__7, addout_21__6, addout_21__5, 
         addout_21__4, addout_21__3, addout_21__2, addout_21__1, addout_21__0, 
         addout_22__31, addout_22__30, addout_22__29, addout_22__28, 
         addout_22__27, addout_22__26, addout_22__25, addout_22__24, 
         addout_22__23, addout_22__22, addout_22__21, addout_22__20, 
         addout_22__19, addout_22__18, addout_22__17, addout_22__16, 
         addout_22__15, addout_22__14, addout_22__13, addout_22__12, 
         addout_22__11, addout_22__10, addout_22__9, addout_22__8, addout_22__7, 
         addout_22__6, addout_22__5, addout_22__4, addout_22__3, addout_22__2, 
         addout_22__1, addout_22__0, addout_23__31, addout_23__30, addout_23__29, 
         addout_23__28, addout_23__27, addout_23__26, addout_23__25, 
         addout_23__24, addout_23__23, addout_23__22, addout_23__21, 
         addout_23__20, addout_23__19, addout_23__18, addout_23__17, 
         addout_23__16, addout_23__15, addout_23__14, addout_23__13, 
         addout_23__12, addout_23__11, addout_23__10, addout_23__9, addout_23__8, 
         addout_23__7, addout_23__6, addout_23__5, addout_23__4, addout_23__3, 
         addout_23__2, addout_23__1, addout_23__0, addout_24__31, addout_24__30, 
         addout_24__29, addout_24__28, addout_24__27, addout_24__26, 
         addout_24__25, addout_24__24, addout_24__23, addout_24__22, 
         addout_24__21, addout_24__20, addout_24__19, addout_24__18, 
         addout_24__17, addout_24__16, addout_24__15, addout_24__14, 
         addout_24__13, addout_24__12, addout_24__11, addout_24__10, 
         addout_24__9, addout_24__8, addout_24__7, addout_24__6, addout_24__5, 
         addout_24__4, addout_24__3, addout_24__2, addout_24__1, addout_24__0, 
         addout_25__31, addout_25__30, addout_25__29, addout_25__28, 
         addout_25__27, addout_25__26, addout_25__25, addout_25__24, 
         addout_25__23, addout_25__22, addout_25__21, addout_25__20, 
         addout_25__19, addout_25__18, addout_25__17, addout_25__16, 
         addout_25__15, addout_25__14, addout_25__13, addout_25__12, 
         addout_25__11, addout_25__10, addout_25__9, addout_25__8, addout_25__7, 
         addout_25__6, addout_25__5, addout_25__4, addout_25__3, addout_25__2, 
         addout_25__1, addout_25__0, addout_26__31, addout_26__30, addout_26__29, 
         addout_26__28, addout_26__27, addout_26__26, addout_26__25, 
         addout_26__24, addout_26__23, addout_26__22, addout_26__21, 
         addout_26__20, addout_26__19, addout_26__18, addout_26__17, 
         addout_26__16, addout_26__15, addout_26__14, addout_26__13, 
         addout_26__12, addout_26__11, addout_26__10, addout_26__9, addout_26__8, 
         addout_26__7, addout_26__6, addout_26__5, addout_26__4, addout_26__3, 
         addout_26__2, addout_26__1, addout_26__0, addout_27__31, addout_27__30, 
         addout_27__29, addout_27__28, addout_27__27, addout_27__26, 
         addout_27__25, addout_27__24, addout_27__23, addout_27__22, 
         addout_27__21, addout_27__20, addout_27__19, addout_27__18, 
         addout_27__17, addout_27__16, addout_27__15, addout_27__14, 
         addout_27__13, addout_27__12, addout_27__11, addout_27__10, 
         addout_27__9, addout_27__8, addout_27__7, addout_27__6, addout_27__5, 
         addout_27__4, addout_27__3, addout_27__2, addout_27__1, addout_27__0, 
         addout_28__31, addout_28__30, addout_28__29, addout_28__28, 
         addout_28__27, addout_28__26, addout_28__25, addout_28__24, 
         addout_28__23, addout_28__22, addout_28__21, addout_28__20, 
         addout_28__19, addout_28__18, addout_28__17, addout_28__16, 
         addout_28__15, addout_28__14, addout_28__13, addout_28__12, 
         addout_28__11, addout_28__10, addout_28__9, addout_28__8, addout_28__7, 
         addout_28__6, addout_28__5, addout_28__4, addout_28__3, addout_28__2, 
         addout_28__1, addout_28__0, addout_29__31, addout_29__30, addout_29__29, 
         addout_29__28, addout_29__27, addout_29__26, addout_29__25, 
         addout_29__24, addout_29__23, addout_29__22, addout_29__21, 
         addout_29__20, addout_29__19, addout_29__18, addout_29__17, 
         addout_29__16, addout_29__15, addout_29__14, addout_29__13, 
         addout_29__12, addout_29__11, addout_29__10, addout_29__9, addout_29__8, 
         addout_29__7, addout_29__6, addout_29__5, addout_29__4, addout_29__3, 
         addout_29__2, addout_29__1, addout_29__0, op2_0__15, op2_0__14, 
         op2_0__13, op2_0__12, op2_0__11, op2_0__10, op2_0__9, op2_0__8, 
         op2_0__7, op2_0__6, op2_0__5, op2_0__4, op2_0__3, op2_0__2, op2_0__1, 
         op2_1__16, op2_1__15, op2_1__14, op2_1__13, op2_1__12, op2_1__11, 
         op2_1__10, op2_1__9, op2_1__8, op2_1__7, op2_1__6, op2_1__5, op2_1__4, 
         op2_1__3, op2_1__2, op2_2__17, op2_2__16, op2_2__15, op2_2__14, 
         op2_2__13, op2_2__12, op2_2__11, op2_2__10, op2_2__9, op2_2__8, 
         op2_2__7, op2_2__6, op2_2__5, op2_2__4, op2_2__3, op2_3__18, op2_3__17, 
         op2_3__16, op2_3__15, op2_3__14, op2_3__13, op2_3__12, op2_3__11, 
         op2_3__10, op2_3__9, op2_3__8, op2_3__7, op2_3__6, op2_3__5, op2_3__4, 
         op2_4__19, op2_4__18, op2_4__17, op2_4__16, op2_4__15, op2_4__14, 
         op2_4__13, op2_4__12, op2_4__11, op2_4__10, op2_4__9, op2_4__8, 
         op2_4__7, op2_4__6, op2_4__5, op2_5__20, op2_5__19, op2_5__18, 
         op2_5__17, op2_5__16, op2_5__15, op2_5__14, op2_5__13, op2_5__12, 
         op2_5__11, op2_5__10, op2_5__9, op2_5__8, op2_5__7, op2_5__6, op2_6__21, 
         op2_6__20, op2_6__19, op2_6__18, op2_6__17, op2_6__16, op2_6__15, 
         op2_6__14, op2_6__13, op2_6__12, op2_6__11, op2_6__10, op2_6__9, 
         op2_6__8, op2_6__7, op2_7__22, op2_7__21, op2_7__20, op2_7__19, 
         op2_7__18, op2_7__17, op2_7__16, op2_7__15, op2_7__14, op2_7__13, 
         op2_7__12, op2_7__11, op2_7__10, op2_7__9, op2_7__8, op2_8__23, 
         op2_8__22, op2_8__21, op2_8__20, op2_8__19, op2_8__18, op2_8__17, 
         op2_8__16, op2_8__15, op2_8__14, op2_8__13, op2_8__12, op2_8__11, 
         op2_8__10, op2_8__9, op2_9__24, op2_9__23, op2_9__22, op2_9__21, 
         op2_9__20, op2_9__19, op2_9__18, op2_9__17, op2_9__16, op2_9__15, 
         op2_9__14, op2_9__13, op2_9__12, op2_9__11, op2_9__10, op2_10__26, 
         op2_10__25, op2_10__24, op2_10__23, op2_10__22, op2_10__21, op2_10__20, 
         op2_10__19, op2_10__18, op2_10__17, op2_10__16, op2_10__15, op2_10__14, 
         op2_10__13, op2_10__12, op2_10__11, op2_11__27, op2_11__26, op2_11__25, 
         op2_11__24, op2_11__23, op2_11__22, op2_11__21, op2_11__20, op2_11__19, 
         op2_11__18, op2_11__17, op2_11__16, op2_11__15, op2_11__14, op2_11__13, 
         op2_11__12, op2_12__28, op2_12__27, op2_12__26, op2_12__25, op2_12__24, 
         op2_12__23, op2_12__22, op2_12__21, op2_12__20, op2_12__19, op2_12__18, 
         op2_12__17, op2_12__16, op2_12__15, op2_12__14, op2_12__13, op2_13__29, 
         op2_13__28, op2_13__27, op2_13__26, op2_13__25, op2_13__24, op2_13__23, 
         op2_13__22, op2_13__21, op2_13__20, op2_13__19, op2_13__18, op2_13__17, 
         op2_13__16, op2_13__15, op2_13__14, op2_14__30, op2_14__29, op2_14__28, 
         op2_14__27, op2_14__26, op1_14, op1_13, op1_12, op1_11, op1_10, op1_9, 
         op1_8, op1_7, op1_6, op1_5, op1_4, op1_3, op1_2, op1_1, op1_0, 
         addout_31__31, nx5768, nx5770, nx5772, nx5774, nx5776, nx5778, nx5780, 
         nx5782, nx5784, nx5786, nx5788, nx5790, nx5792, nx5794, nx5796, nx5798, 
         nx5800, nx5802, nx5804, nx5806, nx5808, nx5810, nx5812, nx5814, nx5816, 
         nx5818, nx5820, nx5822, nx5824, nx5826, nx5828, nx5830, nx5832, nx5834, 
         nx5836, nx5838, nx5840, nx5842, nx5844, nx5846, nx5848, nx5850, nx5852, 
         nx5854, nx5856, nx5858, nx5860, nx5862, nx5864, nx5866, nx5868, nx5870, 
         nx5872, nx5874, nx5876, nx5878, nx5880, nx5882, nx5884, nx5886, nx5888, 
         nx5890, nx5892, nx5894, nx5896, nx5898, nx5900, nx5902, nx5904, nx5906, 
         nx5908, nx5910, nx5912, nx5914, nx5916, nx5918, nx5920, nx5922, nx5924, 
         nx5926, nx5928, nx5930, nx5932, nx5934, nx5936, nx5938, nx5940, nx5942, 
         nx5944, nx5946, nx5948, nx5950, nx5952, nx5954, nx5956, nx5958, nx5960, 
         nx5962, nx5964, nx5966, nx5968, nx5970, nx5972, nx5974, nx5976, nx5978, 
         nx5980, nx5982, nx5984, nx5986, nx5988, nx5990, nx5992, nx5994, nx5996, 
         nx5998, nx6000, nx6002, nx6004, nx6006, nx6008, nx6010, nx6012, nx6014, 
         nx6016, nx6018, nx6020, nx6022, nx6024, nx6026, nx6224, nx6226, nx6228, 
         nx6230, nx6232, nx6234, nx6236, nx6238, nx6240, nx6242, nx6244, nx6246, 
         nx6248, nx6250, nx6252, nx6254, nx6256, nx6258, nx6260, nx6262, nx6264, 
         nx6266, nx6268, nx6270, nx6272, nx6274, nx6276, nx6278, nx6280, nx6282, 
         nx6284, nx6286, nx6288, nx6290, nx6292, nx6294, nx6296, nx6298, nx6300, 
         nx6302, nx6304, nx6306, nx6308, nx6310, nx6312, nx6314, nx6316, nx6318, 
         nx6320, nx6322, nx6324, nx6326, nx6328, nx6330, nx6332, nx6334, nx6336, 
         nx6338, nx6340, nx6342, nx6344, nx6346, nx6348, nx6350, nx6352, nx6354, 
         nx6356, nx6358, nx6360, nx6362, nx6364, nx6366, nx6368, nx6370, nx6372, 
         nx6374, nx6376, nx6378, nx6380, nx6382, nx6384, nx6386, nx6388, nx6390, 
         nx6392, nx6394, nx6396, nx6398, nx6400, nx6402, nx6404, nx6406, nx6408, 
         nx6410, nx6412, nx6414, nx6416, nx6418, nx6420, nx6422, nx6424, nx6426, 
         nx6428, nx6430, nx6432, nx6434, nx6436, nx6438, nx6440, nx6442, nx6444, 
         nx6446, nx6448, nx6450, nx6452, nx6454, nx6456, nx6458, nx6460, nx6462, 
         nx6464, nx6466, nx6468, nx6470, nx6472, nx6474, nx6476, nx6478, nx6480, 
         nx6482, nx6484;



    FC_nadder_32 f0 (.aa ({nx6026,nx6026,nx6024,nx6024,nx6024,nx6022,nx6022,
                 nx6022,nx6020,nx6020,nx6020,nx6018,nx6018,nx6018,nx6016,nx6016,
                 nx6016,op1_14,op1_13,op1_12,op1_11,op1_10,op1_9,op1_8,op1_7,
                 op1_6,op1_5,op1_4,op1_3,op1_2,op1_1,op1_0}), .bb ({nx5780,
                 nx5778,nx5778,nx5778,nx5776,nx5776,nx5776,nx5774,nx5774,nx5774,
                 nx5772,nx5772,nx5772,nx5770,nx5770,nx5770,op2_0__15,op2_0__14,
                 op2_0__13,op2_0__12,op2_0__11,op2_0__10,op2_0__9,op2_0__8,
                 op2_0__7,op2_0__6,op2_0__5,op2_0__4,op2_0__3,op2_0__2,op2_0__1,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({addout_0__31,
                 addout_0__30,addout_0__29,addout_0__28,addout_0__27,
                 addout_0__26,addout_0__25,addout_0__24,addout_0__23,
                 addout_0__22,addout_0__21,addout_0__20,addout_0__19,
                 addout_0__18,addout_0__17,addout_0__16,addout_0__15,
                 addout_0__14,addout_0__13,addout_0__12,addout_0__11,
                 addout_0__10,addout_0__9,addout_0__8,addout_0__7,addout_0__6,
                 addout_0__5,addout_0__4,addout_0__3,addout_0__2,addout_0__1,
                 addout_0__0})) ;
    FC_nadder_32 loop3_1_fx (.aa ({addout_0__31,addout_0__30,addout_0__29,
                 addout_0__28,addout_0__27,addout_0__26,addout_0__25,
                 addout_0__24,addout_0__23,addout_0__22,addout_0__21,
                 addout_0__20,addout_0__19,addout_0__18,addout_0__17,
                 addout_0__16,addout_0__15,addout_0__14,addout_0__13,
                 addout_0__12,addout_0__11,addout_0__10,addout_0__9,addout_0__8,
                 addout_0__7,addout_0__6,addout_0__5,addout_0__4,addout_0__3,
                 addout_0__2,addout_0__1,addout_0__0}), .bb ({nx5792,nx5792,
                 nx5792,nx5790,nx5790,nx5790,nx5788,nx5788,nx5788,nx5786,nx5786,
                 nx5786,nx5784,nx5784,nx5784,op2_1__16,op2_1__15,op2_1__14,
                 op2_1__13,op2_1__12,op2_1__11,op2_1__10,op2_1__9,op2_1__8,
                 op2_1__7,op2_1__6,op2_1__5,op2_1__4,op2_1__3,op2_1__2,
                 addout_31__31,addout_31__31}), .c_cin (addout_31__31), .ff ({
                 addout_1__31,addout_1__30,addout_1__29,addout_1__28,
                 addout_1__27,addout_1__26,addout_1__25,addout_1__24,
                 addout_1__23,addout_1__22,addout_1__21,addout_1__20,
                 addout_1__19,addout_1__18,addout_1__17,addout_1__16,
                 addout_1__15,addout_1__14,addout_1__13,addout_1__12,
                 addout_1__11,addout_1__10,addout_1__9,addout_1__8,addout_1__7,
                 addout_1__6,addout_1__5,addout_1__4,addout_1__3,addout_1__2,
                 addout_1__1,addout_1__0})) ;
    FC_nadder_32 loop3_2_fx (.aa ({addout_1__31,addout_1__30,addout_1__29,
                 addout_1__28,addout_1__27,addout_1__26,addout_1__25,
                 addout_1__24,addout_1__23,addout_1__22,addout_1__21,
                 addout_1__20,addout_1__19,addout_1__18,addout_1__17,
                 addout_1__16,addout_1__15,addout_1__14,addout_1__13,
                 addout_1__12,addout_1__11,addout_1__10,addout_1__9,addout_1__8,
                 addout_1__7,addout_1__6,addout_1__5,addout_1__4,addout_1__3,
                 addout_1__2,addout_1__1,addout_1__0}), .bb ({nx5804,nx5804,
                 nx5802,nx5802,nx5802,nx5800,nx5800,nx5800,nx5798,nx5798,nx5798,
                 nx5796,nx5796,nx5796,op2_2__17,op2_2__16,op2_2__15,op2_2__14,
                 op2_2__13,op2_2__12,op2_2__11,op2_2__10,op2_2__9,op2_2__8,
                 op2_2__7,op2_2__6,op2_2__5,op2_2__4,op2_2__3,addout_31__31,
                 addout_31__31,addout_31__31}), .c_cin (addout_31__31), .ff ({
                 addout_2__31,addout_2__30,addout_2__29,addout_2__28,
                 addout_2__27,addout_2__26,addout_2__25,addout_2__24,
                 addout_2__23,addout_2__22,addout_2__21,addout_2__20,
                 addout_2__19,addout_2__18,addout_2__17,addout_2__16,
                 addout_2__15,addout_2__14,addout_2__13,addout_2__12,
                 addout_2__11,addout_2__10,addout_2__9,addout_2__8,addout_2__7,
                 addout_2__6,addout_2__5,addout_2__4,addout_2__3,addout_2__2,
                 addout_2__1,addout_2__0})) ;
    FC_nadder_32 loop3_3_fx (.aa ({addout_2__31,addout_2__30,addout_2__29,
                 addout_2__28,addout_2__27,addout_2__26,addout_2__25,
                 addout_2__24,addout_2__23,addout_2__22,addout_2__21,
                 addout_2__20,addout_2__19,addout_2__18,addout_2__17,
                 addout_2__16,addout_2__15,addout_2__14,addout_2__13,
                 addout_2__12,addout_2__11,addout_2__10,addout_2__9,addout_2__8,
                 addout_2__7,addout_2__6,addout_2__5,addout_2__4,addout_2__3,
                 addout_2__2,addout_2__1,addout_2__0}), .bb ({nx5816,nx5814,
                 nx5814,nx5814,nx5812,nx5812,nx5812,nx5810,nx5810,nx5810,nx5808,
                 nx5808,nx5808,op2_3__18,op2_3__17,op2_3__16,op2_3__15,op2_3__14
                 ,op2_3__13,op2_3__12,op2_3__11,op2_3__10,op2_3__9,op2_3__8,
                 op2_3__7,op2_3__6,op2_3__5,op2_3__4,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31}), .c_cin (addout_31__31), .ff ({
                 addout_3__31,addout_3__30,addout_3__29,addout_3__28,
                 addout_3__27,addout_3__26,addout_3__25,addout_3__24,
                 addout_3__23,addout_3__22,addout_3__21,addout_3__20,
                 addout_3__19,addout_3__18,addout_3__17,addout_3__16,
                 addout_3__15,addout_3__14,addout_3__13,addout_3__12,
                 addout_3__11,addout_3__10,addout_3__9,addout_3__8,addout_3__7,
                 addout_3__6,addout_3__5,addout_3__4,addout_3__3,addout_3__2,
                 addout_3__1,addout_3__0})) ;
    FC_nadder_32 loop3_4_fx (.aa ({addout_3__31,addout_3__30,addout_3__29,
                 addout_3__28,addout_3__27,addout_3__26,addout_3__25,
                 addout_3__24,addout_3__23,addout_3__22,addout_3__21,
                 addout_3__20,addout_3__19,addout_3__18,addout_3__17,
                 addout_3__16,addout_3__15,addout_3__14,addout_3__13,
                 addout_3__12,addout_3__11,addout_3__10,addout_3__9,addout_3__8,
                 addout_3__7,addout_3__6,addout_3__5,addout_3__4,addout_3__3,
                 addout_3__2,addout_3__1,addout_3__0}), .bb ({nx5826,nx5826,
                 nx5826,nx5824,nx5824,nx5824,nx5822,nx5822,nx5822,nx5820,nx5820,
                 nx5820,op2_4__19,op2_4__18,op2_4__17,op2_4__16,op2_4__15,
                 op2_4__14,op2_4__13,op2_4__12,op2_4__11,op2_4__10,op2_4__9,
                 op2_4__8,op2_4__7,op2_4__6,op2_4__5,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_4__31,addout_4__30,addout_4__29,
                 addout_4__28,addout_4__27,addout_4__26,addout_4__25,
                 addout_4__24,addout_4__23,addout_4__22,addout_4__21,
                 addout_4__20,addout_4__19,addout_4__18,addout_4__17,
                 addout_4__16,addout_4__15,addout_4__14,addout_4__13,
                 addout_4__12,addout_4__11,addout_4__10,addout_4__9,addout_4__8,
                 addout_4__7,addout_4__6,addout_4__5,addout_4__4,addout_4__3,
                 addout_4__2,addout_4__1,addout_4__0})) ;
    FC_nadder_32 loop3_5_fx (.aa ({addout_4__31,addout_4__30,addout_4__29,
                 addout_4__28,addout_4__27,addout_4__26,addout_4__25,
                 addout_4__24,addout_4__23,addout_4__22,addout_4__21,
                 addout_4__20,addout_4__19,addout_4__18,addout_4__17,
                 addout_4__16,addout_4__15,addout_4__14,addout_4__13,
                 addout_4__12,addout_4__11,addout_4__10,addout_4__9,addout_4__8,
                 addout_4__7,addout_4__6,addout_4__5,addout_4__4,addout_4__3,
                 addout_4__2,addout_4__1,addout_4__0}), .bb ({nx5836,nx5836,
                 nx5834,nx5834,nx5834,nx5832,nx5832,nx5832,nx5830,nx5830,nx5830,
                 op2_5__20,op2_5__19,op2_5__18,op2_5__17,op2_5__16,op2_5__15,
                 op2_5__14,op2_5__13,op2_5__12,op2_5__11,op2_5__10,op2_5__9,
                 op2_5__8,op2_5__7,op2_5__6,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_5__31,addout_5__30,addout_5__29,
                 addout_5__28,addout_5__27,addout_5__26,addout_5__25,
                 addout_5__24,addout_5__23,addout_5__22,addout_5__21,
                 addout_5__20,addout_5__19,addout_5__18,addout_5__17,
                 addout_5__16,addout_5__15,addout_5__14,addout_5__13,
                 addout_5__12,addout_5__11,addout_5__10,addout_5__9,addout_5__8,
                 addout_5__7,addout_5__6,addout_5__5,addout_5__4,addout_5__3,
                 addout_5__2,addout_5__1,addout_5__0})) ;
    FC_nadder_32 loop3_6_fx (.aa ({addout_5__31,addout_5__30,addout_5__29,
                 addout_5__28,addout_5__27,addout_5__26,addout_5__25,
                 addout_5__24,addout_5__23,addout_5__22,addout_5__21,
                 addout_5__20,addout_5__19,addout_5__18,addout_5__17,
                 addout_5__16,addout_5__15,addout_5__14,addout_5__13,
                 addout_5__12,addout_5__11,addout_5__10,addout_5__9,addout_5__8,
                 addout_5__7,addout_5__6,addout_5__5,addout_5__4,addout_5__3,
                 addout_5__2,addout_5__1,addout_5__0}), .bb ({nx5846,nx5844,
                 nx5844,nx5844,nx5842,nx5842,nx5842,nx5840,nx5840,nx5840,
                 op2_6__21,op2_6__20,op2_6__19,op2_6__18,op2_6__17,op2_6__16,
                 op2_6__15,op2_6__14,op2_6__13,op2_6__12,op2_6__11,op2_6__10,
                 op2_6__9,op2_6__8,op2_6__7,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({addout_6__31,
                 addout_6__30,addout_6__29,addout_6__28,addout_6__27,
                 addout_6__26,addout_6__25,addout_6__24,addout_6__23,
                 addout_6__22,addout_6__21,addout_6__20,addout_6__19,
                 addout_6__18,addout_6__17,addout_6__16,addout_6__15,
                 addout_6__14,addout_6__13,addout_6__12,addout_6__11,
                 addout_6__10,addout_6__9,addout_6__8,addout_6__7,addout_6__6,
                 addout_6__5,addout_6__4,addout_6__3,addout_6__2,addout_6__1,
                 addout_6__0})) ;
    FC_nadder_32 loop3_7_fx (.aa ({addout_6__31,addout_6__30,addout_6__29,
                 addout_6__28,addout_6__27,addout_6__26,addout_6__25,
                 addout_6__24,addout_6__23,addout_6__22,addout_6__21,
                 addout_6__20,addout_6__19,addout_6__18,addout_6__17,
                 addout_6__16,addout_6__15,addout_6__14,addout_6__13,
                 addout_6__12,addout_6__11,addout_6__10,addout_6__9,addout_6__8,
                 addout_6__7,addout_6__6,addout_6__5,addout_6__4,addout_6__3,
                 addout_6__2,addout_6__1,addout_6__0}), .bb ({nx5854,nx5854,
                 nx5854,nx5852,nx5852,nx5852,nx5850,nx5850,nx5850,op2_7__22,
                 op2_7__21,op2_7__20,op2_7__19,op2_7__18,op2_7__17,op2_7__16,
                 op2_7__15,op2_7__14,op2_7__13,op2_7__12,op2_7__11,op2_7__10,
                 op2_7__9,op2_7__8,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({addout_7__31,
                 addout_7__30,addout_7__29,addout_7__28,addout_7__27,
                 addout_7__26,addout_7__25,addout_7__24,addout_7__23,
                 addout_7__22,addout_7__21,addout_7__20,addout_7__19,
                 addout_7__18,addout_7__17,addout_7__16,addout_7__15,
                 addout_7__14,addout_7__13,addout_7__12,addout_7__11,
                 addout_7__10,addout_7__9,addout_7__8,addout_7__7,addout_7__6,
                 addout_7__5,addout_7__4,addout_7__3,addout_7__2,addout_7__1,
                 addout_7__0})) ;
    FC_nadder_32 loop3_8_fx (.aa ({addout_7__31,addout_7__30,addout_7__29,
                 addout_7__28,addout_7__27,addout_7__26,addout_7__25,
                 addout_7__24,addout_7__23,addout_7__22,addout_7__21,
                 addout_7__20,addout_7__19,addout_7__18,addout_7__17,
                 addout_7__16,addout_7__15,addout_7__14,addout_7__13,
                 addout_7__12,addout_7__11,addout_7__10,addout_7__9,addout_7__8,
                 addout_7__7,addout_7__6,addout_7__5,addout_7__4,addout_7__3,
                 addout_7__2,addout_7__1,addout_7__0}), .bb ({nx5862,nx5862,
                 nx5860,nx5860,nx5860,nx5858,nx5858,nx5858,op2_8__23,op2_8__22,
                 op2_8__21,op2_8__20,op2_8__19,op2_8__18,op2_8__17,op2_8__16,
                 op2_8__15,op2_8__14,op2_8__13,op2_8__12,op2_8__11,op2_8__10,
                 op2_8__9,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31}), .c_cin (addout_31__31), .ff ({
                 addout_8__31,addout_8__30,addout_8__29,addout_8__28,
                 addout_8__27,addout_8__26,addout_8__25,addout_8__24,
                 addout_8__23,addout_8__22,addout_8__21,addout_8__20,
                 addout_8__19,addout_8__18,addout_8__17,addout_8__16,
                 addout_8__15,addout_8__14,addout_8__13,addout_8__12,
                 addout_8__11,addout_8__10,addout_8__9,addout_8__8,addout_8__7,
                 addout_8__6,addout_8__5,addout_8__4,addout_8__3,addout_8__2,
                 addout_8__1,addout_8__0})) ;
    FC_nadder_32 loop3_9_fx (.aa ({addout_8__31,addout_8__30,addout_8__29,
                 addout_8__28,addout_8__27,addout_8__26,addout_8__25,
                 addout_8__24,addout_8__23,addout_8__22,addout_8__21,
                 addout_8__20,addout_8__19,addout_8__18,addout_8__17,
                 addout_8__16,addout_8__15,addout_8__14,addout_8__13,
                 addout_8__12,addout_8__11,addout_8__10,addout_8__9,addout_8__8,
                 addout_8__7,addout_8__6,addout_8__5,addout_8__4,addout_8__3,
                 addout_8__2,addout_8__1,addout_8__0}), .bb ({nx5870,nx5868,
                 nx5868,nx5868,nx5866,nx5866,nx5866,op2_9__24,op2_9__23,
                 op2_9__22,op2_9__21,op2_9__20,op2_9__19,op2_9__18,op2_9__17,
                 op2_9__16,op2_9__15,op2_9__14,op2_9__13,op2_9__12,op2_9__11,
                 op2_9__10,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_9__31,addout_9__30,addout_9__29,
                 addout_9__28,addout_9__27,addout_9__26,addout_9__25,
                 addout_9__24,addout_9__23,addout_9__22,addout_9__21,
                 addout_9__20,addout_9__19,addout_9__18,addout_9__17,
                 addout_9__16,addout_9__15,addout_9__14,addout_9__13,
                 addout_9__12,addout_9__11,addout_9__10,addout_9__9,addout_9__8,
                 addout_9__7,addout_9__6,addout_9__5,addout_9__4,addout_9__3,
                 addout_9__2,addout_9__1,addout_9__0})) ;
    FC_nadder_32 loop3_10_fx (.aa ({addout_9__31,addout_9__30,addout_9__29,
                 addout_9__28,addout_9__27,addout_9__26,addout_9__25,
                 addout_9__24,addout_9__23,addout_9__22,addout_9__21,
                 addout_9__20,addout_9__19,addout_9__18,addout_9__17,
                 addout_9__16,addout_9__15,addout_9__14,addout_9__13,
                 addout_9__12,addout_9__11,addout_9__10,addout_9__9,addout_9__8,
                 addout_9__7,addout_9__6,addout_9__5,addout_9__4,addout_9__3,
                 addout_9__2,addout_9__1,addout_9__0}), .bb ({nx5874,nx5874,
                 nx5874,nx5872,nx5872,nx5872,op2_10__25,op2_10__24,op2_10__23,
                 op2_10__22,op2_10__21,op2_10__20,op2_10__19,op2_10__18,
                 op2_10__17,op2_10__16,op2_10__15,op2_10__14,op2_10__13,
                 op2_10__12,op2_10__11,addout_31__31,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_10__31,addout_10__30,addout_10__29
                 ,addout_10__28,addout_10__27,addout_10__26,addout_10__25,
                 addout_10__24,addout_10__23,addout_10__22,addout_10__21,
                 addout_10__20,addout_10__19,addout_10__18,addout_10__17,
                 addout_10__16,addout_10__15,addout_10__14,addout_10__13,
                 addout_10__12,addout_10__11,addout_10__10,addout_10__9,
                 addout_10__8,addout_10__7,addout_10__6,addout_10__5,
                 addout_10__4,addout_10__3,addout_10__2,addout_10__1,
                 addout_10__0})) ;
    FC_nadder_32 loop3_11_fx (.aa ({addout_10__31,addout_10__30,addout_10__29,
                 addout_10__28,addout_10__27,addout_10__26,addout_10__25,
                 addout_10__24,addout_10__23,addout_10__22,addout_10__21,
                 addout_10__20,addout_10__19,addout_10__18,addout_10__17,
                 addout_10__16,addout_10__15,addout_10__14,addout_10__13,
                 addout_10__12,addout_10__11,addout_10__10,addout_10__9,
                 addout_10__8,addout_10__7,addout_10__6,addout_10__5,
                 addout_10__4,addout_10__3,addout_10__2,addout_10__1,
                 addout_10__0}), .bb ({nx5878,nx5878,nx5876,nx5876,nx5876,
                 op2_11__26,op2_11__25,op2_11__24,op2_11__23,op2_11__22,
                 op2_11__21,op2_11__20,op2_11__19,op2_11__18,op2_11__17,
                 op2_11__16,op2_11__15,op2_11__14,op2_11__13,op2_11__12,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_11__31,addout_11__30,addout_11__29
                 ,addout_11__28,addout_11__27,addout_11__26,addout_11__25,
                 addout_11__24,addout_11__23,addout_11__22,addout_11__21,
                 addout_11__20,addout_11__19,addout_11__18,addout_11__17,
                 addout_11__16,addout_11__15,addout_11__14,addout_11__13,
                 addout_11__12,addout_11__11,addout_11__10,addout_11__9,
                 addout_11__8,addout_11__7,addout_11__6,addout_11__5,
                 addout_11__4,addout_11__3,addout_11__2,addout_11__1,
                 addout_11__0})) ;
    FC_nadder_32 loop3_12_fx (.aa ({addout_11__31,addout_11__30,addout_11__29,
                 addout_11__28,addout_11__27,addout_11__26,addout_11__25,
                 addout_11__24,addout_11__23,addout_11__22,addout_11__21,
                 addout_11__20,addout_11__19,addout_11__18,addout_11__17,
                 addout_11__16,addout_11__15,addout_11__14,addout_11__13,
                 addout_11__12,addout_11__11,addout_11__10,addout_11__9,
                 addout_11__8,addout_11__7,addout_11__6,addout_11__5,
                 addout_11__4,addout_11__3,addout_11__2,addout_11__1,
                 addout_11__0}), .bb ({nx5882,nx5880,nx5880,nx5880,op2_12__27,
                 op2_12__26,op2_12__25,op2_12__24,op2_12__23,op2_12__22,
                 op2_12__21,op2_12__20,op2_12__19,op2_12__18,op2_12__17,
                 op2_12__16,op2_12__15,op2_12__14,op2_12__13,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_12__31,addout_12__30,addout_12__29
                 ,addout_12__28,addout_12__27,addout_12__26,addout_12__25,
                 addout_12__24,addout_12__23,addout_12__22,addout_12__21,
                 addout_12__20,addout_12__19,addout_12__18,addout_12__17,
                 addout_12__16,addout_12__15,addout_12__14,addout_12__13,
                 addout_12__12,addout_12__11,addout_12__10,addout_12__9,
                 addout_12__8,addout_12__7,addout_12__6,addout_12__5,
                 addout_12__4,addout_12__3,addout_12__2,addout_12__1,
                 addout_12__0})) ;
    FC_nadder_32 loop3_13_fx (.aa ({addout_12__31,addout_12__30,addout_12__29,
                 addout_12__28,addout_12__27,addout_12__26,addout_12__25,
                 addout_12__24,addout_12__23,addout_12__22,addout_12__21,
                 addout_12__20,addout_12__19,addout_12__18,addout_12__17,
                 addout_12__16,addout_12__15,addout_12__14,addout_12__13,
                 addout_12__12,addout_12__11,addout_12__10,addout_12__9,
                 addout_12__8,addout_12__7,addout_12__6,addout_12__5,
                 addout_12__4,addout_12__3,addout_12__2,addout_12__1,
                 addout_12__0}), .bb ({nx6480,nx6480,nx6480,op2_13__28,
                 op2_13__27,op2_13__26,op2_13__25,op2_13__24,op2_13__23,
                 op2_13__22,op2_13__21,op2_13__20,op2_13__19,op2_13__18,
                 op2_13__17,op2_13__16,op2_13__15,op2_13__14,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({addout_13__31,
                 addout_13__30,addout_13__29,addout_13__28,addout_13__27,
                 addout_13__26,addout_13__25,addout_13__24,addout_13__23,
                 addout_13__22,addout_13__21,addout_13__20,addout_13__19,
                 addout_13__18,addout_13__17,addout_13__16,addout_13__15,
                 addout_13__14,addout_13__13,addout_13__12,addout_13__11,
                 addout_13__10,addout_13__9,addout_13__8,addout_13__7,
                 addout_13__6,addout_13__5,addout_13__4,addout_13__3,
                 addout_13__2,addout_13__1,addout_13__0})) ;
    FC_nadder_32 loop3_14_fx (.aa ({addout_13__31,addout_13__30,addout_13__29,
                 addout_13__28,addout_13__27,addout_13__26,addout_13__25,
                 addout_13__24,addout_13__23,addout_13__22,addout_13__21,
                 addout_13__20,addout_13__19,addout_13__18,addout_13__17,
                 addout_13__16,addout_13__15,addout_13__14,addout_13__13,
                 addout_13__12,addout_13__11,addout_13__10,addout_13__9,
                 addout_13__8,addout_13__7,addout_13__6,addout_13__5,
                 addout_13__4,addout_13__3,addout_13__2,addout_13__1,
                 addout_13__0}), .bb ({nx6482,nx6482,nx6484,nx5884,nx5888,nx5892
                 ,nx5898,nx5906,nx5914,nx5922,nx5932,nx5942,nx5952,nx5964,nx5976
                 ,nx5988,nx6002,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_14__31,addout_14__30,addout_14__29
                 ,addout_14__28,addout_14__27,addout_14__26,addout_14__25,
                 addout_14__24,addout_14__23,addout_14__22,addout_14__21,
                 addout_14__20,addout_14__19,addout_14__18,addout_14__17,
                 addout_14__16,addout_14__15,addout_14__14,addout_14__13,
                 addout_14__12,addout_14__11,addout_14__10,addout_14__9,
                 addout_14__8,addout_14__7,addout_14__6,addout_14__5,
                 addout_14__4,addout_14__3,addout_14__2,addout_14__1,
                 addout_14__0})) ;
    FC_nadder_32 loop3_15_fx (.aa ({addout_14__31,addout_14__30,addout_14__29,
                 addout_14__28,addout_14__27,addout_14__26,addout_14__25,
                 addout_14__24,addout_14__23,addout_14__22,addout_14__21,
                 addout_14__20,addout_14__19,addout_14__18,addout_14__17,
                 addout_14__16,addout_14__15,addout_14__14,addout_14__13,
                 addout_14__12,addout_14__11,addout_14__10,addout_14__9,
                 addout_14__8,addout_14__7,addout_14__6,addout_14__5,
                 addout_14__4,addout_14__3,addout_14__2,addout_14__1,
                 addout_14__0}), .bb ({nx6482,nx6484,nx5884,nx5888,nx5892,nx5898
                 ,nx5906,nx5914,nx5922,nx5932,nx5942,nx5952,nx5964,nx5976,nx5988
                 ,nx6002,addout_31__31,addout_31__31,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_15__31,addout_15__30,addout_15__29
                 ,addout_15__28,addout_15__27,addout_15__26,addout_15__25,
                 addout_15__24,addout_15__23,addout_15__22,addout_15__21,
                 addout_15__20,addout_15__19,addout_15__18,addout_15__17,
                 addout_15__16,addout_15__15,addout_15__14,addout_15__13,
                 addout_15__12,addout_15__11,addout_15__10,addout_15__9,
                 addout_15__8,addout_15__7,addout_15__6,addout_15__5,
                 addout_15__4,addout_15__3,addout_15__2,addout_15__1,
                 addout_15__0})) ;
    FC_nadder_32 loop3_16_fx (.aa ({addout_15__31,addout_15__30,addout_15__29,
                 addout_15__28,addout_15__27,addout_15__26,addout_15__25,
                 addout_15__24,addout_15__23,addout_15__22,addout_15__21,
                 addout_15__20,addout_15__19,addout_15__18,addout_15__17,
                 addout_15__16,addout_15__15,addout_15__14,addout_15__13,
                 addout_15__12,addout_15__11,addout_15__10,addout_15__9,
                 addout_15__8,addout_15__7,addout_15__6,addout_15__5,
                 addout_15__4,addout_15__3,addout_15__2,addout_15__1,
                 addout_15__0}), .bb ({nx6484,nx5884,nx5888,nx5892,nx5898,nx5906
                 ,nx5914,nx5922,nx5932,nx5942,nx5952,nx5964,nx5976,nx5988,nx6002
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({addout_16__31,
                 addout_16__30,addout_16__29,addout_16__28,addout_16__27,
                 addout_16__26,addout_16__25,addout_16__24,addout_16__23,
                 addout_16__22,addout_16__21,addout_16__20,addout_16__19,
                 addout_16__18,addout_16__17,addout_16__16,addout_16__15,
                 addout_16__14,addout_16__13,addout_16__12,addout_16__11,
                 addout_16__10,addout_16__9,addout_16__8,addout_16__7,
                 addout_16__6,addout_16__5,addout_16__4,addout_16__3,
                 addout_16__2,addout_16__1,addout_16__0})) ;
    FC_nadder_32 loop3_17_fx (.aa ({addout_16__31,addout_16__30,addout_16__29,
                 addout_16__28,addout_16__27,addout_16__26,addout_16__25,
                 addout_16__24,addout_16__23,addout_16__22,addout_16__21,
                 addout_16__20,addout_16__19,addout_16__18,addout_16__17,
                 addout_16__16,addout_16__15,addout_16__14,addout_16__13,
                 addout_16__12,addout_16__11,addout_16__10,addout_16__9,
                 addout_16__8,addout_16__7,addout_16__6,addout_16__5,
                 addout_16__4,addout_16__3,addout_16__2,addout_16__1,
                 addout_16__0}), .bb ({nx5886,nx5890,nx5894,nx5900,nx5908,nx5916
                 ,nx5924,nx5934,nx5944,nx5954,nx5966,nx5978,nx5990,nx6004,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31}), .c_cin (addout_31__31), .ff ({
                 addout_17__31,addout_17__30,addout_17__29,addout_17__28,
                 addout_17__27,addout_17__26,addout_17__25,addout_17__24,
                 addout_17__23,addout_17__22,addout_17__21,addout_17__20,
                 addout_17__19,addout_17__18,addout_17__17,addout_17__16,
                 addout_17__15,addout_17__14,addout_17__13,addout_17__12,
                 addout_17__11,addout_17__10,addout_17__9,addout_17__8,
                 addout_17__7,addout_17__6,addout_17__5,addout_17__4,
                 addout_17__3,addout_17__2,addout_17__1,addout_17__0})) ;
    FC_nadder_32 loop3_18_fx (.aa ({addout_17__31,addout_17__30,addout_17__29,
                 addout_17__28,addout_17__27,addout_17__26,addout_17__25,
                 addout_17__24,addout_17__23,addout_17__22,addout_17__21,
                 addout_17__20,addout_17__19,addout_17__18,addout_17__17,
                 addout_17__16,addout_17__15,addout_17__14,addout_17__13,
                 addout_17__12,addout_17__11,addout_17__10,addout_17__9,
                 addout_17__8,addout_17__7,addout_17__6,addout_17__5,
                 addout_17__4,addout_17__3,addout_17__2,addout_17__1,
                 addout_17__0}), .bb ({nx5890,nx5894,nx5900,nx5908,nx5916,nx5924
                 ,nx5934,nx5944,nx5954,nx5966,nx5978,nx5990,nx6004,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31}), .c_cin (addout_31__31), .ff ({
                 addout_18__31,addout_18__30,addout_18__29,addout_18__28,
                 addout_18__27,addout_18__26,addout_18__25,addout_18__24,
                 addout_18__23,addout_18__22,addout_18__21,addout_18__20,
                 addout_18__19,addout_18__18,addout_18__17,addout_18__16,
                 addout_18__15,addout_18__14,addout_18__13,addout_18__12,
                 addout_18__11,addout_18__10,addout_18__9,addout_18__8,
                 addout_18__7,addout_18__6,addout_18__5,addout_18__4,
                 addout_18__3,addout_18__2,addout_18__1,addout_18__0})) ;
    FC_nadder_32 loop3_19_fx (.aa ({addout_18__31,addout_18__30,addout_18__29,
                 addout_18__28,addout_18__27,addout_18__26,addout_18__25,
                 addout_18__24,addout_18__23,addout_18__22,addout_18__21,
                 addout_18__20,addout_18__19,addout_18__18,addout_18__17,
                 addout_18__16,addout_18__15,addout_18__14,addout_18__13,
                 addout_18__12,addout_18__11,addout_18__10,addout_18__9,
                 addout_18__8,addout_18__7,addout_18__6,addout_18__5,
                 addout_18__4,addout_18__3,addout_18__2,addout_18__1,
                 addout_18__0}), .bb ({nx5894,nx5900,nx5908,nx5916,nx5924,nx5934
                 ,nx5944,nx5954,nx5966,nx5978,nx5990,nx6004,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_19__31,addout_19__30,addout_19__29
                 ,addout_19__28,addout_19__27,addout_19__26,addout_19__25,
                 addout_19__24,addout_19__23,addout_19__22,addout_19__21,
                 addout_19__20,addout_19__19,addout_19__18,addout_19__17,
                 addout_19__16,addout_19__15,addout_19__14,addout_19__13,
                 addout_19__12,addout_19__11,addout_19__10,addout_19__9,
                 addout_19__8,addout_19__7,addout_19__6,addout_19__5,
                 addout_19__4,addout_19__3,addout_19__2,addout_19__1,
                 addout_19__0})) ;
    FC_nadder_32 loop3_20_fx (.aa ({addout_19__31,addout_19__30,addout_19__29,
                 addout_19__28,addout_19__27,addout_19__26,addout_19__25,
                 addout_19__24,addout_19__23,addout_19__22,addout_19__21,
                 addout_19__20,addout_19__19,addout_19__18,addout_19__17,
                 addout_19__16,addout_19__15,addout_19__14,addout_19__13,
                 addout_19__12,addout_19__11,addout_19__10,addout_19__9,
                 addout_19__8,addout_19__7,addout_19__6,addout_19__5,
                 addout_19__4,addout_19__3,addout_19__2,addout_19__1,
                 addout_19__0}), .bb ({nx5902,nx5910,nx5918,nx5926,nx5936,nx5946
                 ,nx5956,nx5968,nx5980,nx5992,nx6006,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_20__31,addout_20__30,addout_20__29
                 ,addout_20__28,addout_20__27,addout_20__26,addout_20__25,
                 addout_20__24,addout_20__23,addout_20__22,addout_20__21,
                 addout_20__20,addout_20__19,addout_20__18,addout_20__17,
                 addout_20__16,addout_20__15,addout_20__14,addout_20__13,
                 addout_20__12,addout_20__11,addout_20__10,addout_20__9,
                 addout_20__8,addout_20__7,addout_20__6,addout_20__5,
                 addout_20__4,addout_20__3,addout_20__2,addout_20__1,
                 addout_20__0})) ;
    FC_nadder_32 loop3_21_fx (.aa ({addout_20__31,addout_20__30,addout_20__29,
                 addout_20__28,addout_20__27,addout_20__26,addout_20__25,
                 addout_20__24,addout_20__23,addout_20__22,addout_20__21,
                 addout_20__20,addout_20__19,addout_20__18,addout_20__17,
                 addout_20__16,addout_20__15,addout_20__14,addout_20__13,
                 addout_20__12,addout_20__11,addout_20__10,addout_20__9,
                 addout_20__8,addout_20__7,addout_20__6,addout_20__5,
                 addout_20__4,addout_20__3,addout_20__2,addout_20__1,
                 addout_20__0}), .bb ({nx5910,nx5918,nx5926,nx5936,nx5946,nx5956
                 ,nx5968,nx5980,nx5992,nx6006,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_21__31,addout_21__30,addout_21__29
                 ,addout_21__28,addout_21__27,addout_21__26,addout_21__25,
                 addout_21__24,addout_21__23,addout_21__22,addout_21__21,
                 addout_21__20,addout_21__19,addout_21__18,addout_21__17,
                 addout_21__16,addout_21__15,addout_21__14,addout_21__13,
                 addout_21__12,addout_21__11,addout_21__10,addout_21__9,
                 addout_21__8,addout_21__7,addout_21__6,addout_21__5,
                 addout_21__4,addout_21__3,addout_21__2,addout_21__1,
                 addout_21__0})) ;
    FC_nadder_32 loop3_22_fx (.aa ({addout_21__31,addout_21__30,addout_21__29,
                 addout_21__28,addout_21__27,addout_21__26,addout_21__25,
                 addout_21__24,addout_21__23,addout_21__22,addout_21__21,
                 addout_21__20,addout_21__19,addout_21__18,addout_21__17,
                 addout_21__16,addout_21__15,addout_21__14,addout_21__13,
                 addout_21__12,addout_21__11,addout_21__10,addout_21__9,
                 addout_21__8,addout_21__7,addout_21__6,addout_21__5,
                 addout_21__4,addout_21__3,addout_21__2,addout_21__1,
                 addout_21__0}), .bb ({nx5918,nx5926,nx5936,nx5946,nx5956,nx5968
                 ,nx5980,nx5992,nx6006,addout_31__31,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_22__31,addout_22__30,addout_22__29
                 ,addout_22__28,addout_22__27,addout_22__26,addout_22__25,
                 addout_22__24,addout_22__23,addout_22__22,addout_22__21,
                 addout_22__20,addout_22__19,addout_22__18,addout_22__17,
                 addout_22__16,addout_22__15,addout_22__14,addout_22__13,
                 addout_22__12,addout_22__11,addout_22__10,addout_22__9,
                 addout_22__8,addout_22__7,addout_22__6,addout_22__5,
                 addout_22__4,addout_22__3,addout_22__2,addout_22__1,
                 addout_22__0})) ;
    FC_nadder_32 loop3_23_fx (.aa ({addout_22__31,addout_22__30,addout_22__29,
                 addout_22__28,addout_22__27,addout_22__26,addout_22__25,
                 addout_22__24,addout_22__23,addout_22__22,addout_22__21,
                 addout_22__20,addout_22__19,addout_22__18,addout_22__17,
                 addout_22__16,addout_22__15,addout_22__14,addout_22__13,
                 addout_22__12,addout_22__11,addout_22__10,addout_22__9,
                 addout_22__8,addout_22__7,addout_22__6,addout_22__5,
                 addout_22__4,addout_22__3,addout_22__2,addout_22__1,
                 addout_22__0}), .bb ({nx5928,nx5938,nx5948,nx5958,nx5970,nx5982
                 ,nx5994,nx6008,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({addout_23__31,
                 addout_23__30,addout_23__29,addout_23__28,addout_23__27,
                 addout_23__26,addout_23__25,addout_23__24,addout_23__23,
                 addout_23__22,addout_23__21,addout_23__20,addout_23__19,
                 addout_23__18,addout_23__17,addout_23__16,addout_23__15,
                 addout_23__14,addout_23__13,addout_23__12,addout_23__11,
                 addout_23__10,addout_23__9,addout_23__8,addout_23__7,
                 addout_23__6,addout_23__5,addout_23__4,addout_23__3,
                 addout_23__2,addout_23__1,addout_23__0})) ;
    FC_nadder_32 loop3_24_fx (.aa ({addout_23__31,addout_23__30,addout_23__29,
                 addout_23__28,addout_23__27,addout_23__26,addout_23__25,
                 addout_23__24,addout_23__23,addout_23__22,addout_23__21,
                 addout_23__20,addout_23__19,addout_23__18,addout_23__17,
                 addout_23__16,addout_23__15,addout_23__14,addout_23__13,
                 addout_23__12,addout_23__11,addout_23__10,addout_23__9,
                 addout_23__8,addout_23__7,addout_23__6,addout_23__5,
                 addout_23__4,addout_23__3,addout_23__2,addout_23__1,
                 addout_23__0}), .bb ({nx5938,nx5948,nx5958,nx5970,nx5982,nx5994
                 ,nx6008,addout_31__31,addout_31__31,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({addout_24__31,
                 addout_24__30,addout_24__29,addout_24__28,addout_24__27,
                 addout_24__26,addout_24__25,addout_24__24,addout_24__23,
                 addout_24__22,addout_24__21,addout_24__20,addout_24__19,
                 addout_24__18,addout_24__17,addout_24__16,addout_24__15,
                 addout_24__14,addout_24__13,addout_24__12,addout_24__11,
                 addout_24__10,addout_24__9,addout_24__8,addout_24__7,
                 addout_24__6,addout_24__5,addout_24__4,addout_24__3,
                 addout_24__2,addout_24__1,addout_24__0})) ;
    FC_nadder_32 loop3_25_fx (.aa ({addout_24__31,addout_24__30,addout_24__29,
                 addout_24__28,addout_24__27,addout_24__26,addout_24__25,
                 addout_24__24,addout_24__23,addout_24__22,addout_24__21,
                 addout_24__20,addout_24__19,addout_24__18,addout_24__17,
                 addout_24__16,addout_24__15,addout_24__14,addout_24__13,
                 addout_24__12,addout_24__11,addout_24__10,addout_24__9,
                 addout_24__8,addout_24__7,addout_24__6,addout_24__5,
                 addout_24__4,addout_24__3,addout_24__2,addout_24__1,
                 addout_24__0}), .bb ({nx5948,nx5958,nx5970,nx5982,nx5994,nx6008
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31}), .c_cin (addout_31__31), .ff ({
                 addout_25__31,addout_25__30,addout_25__29,addout_25__28,
                 addout_25__27,addout_25__26,addout_25__25,addout_25__24,
                 addout_25__23,addout_25__22,addout_25__21,addout_25__20,
                 addout_25__19,addout_25__18,addout_25__17,addout_25__16,
                 addout_25__15,addout_25__14,addout_25__13,addout_25__12,
                 addout_25__11,addout_25__10,addout_25__9,addout_25__8,
                 addout_25__7,addout_25__6,addout_25__5,addout_25__4,
                 addout_25__3,addout_25__2,addout_25__1,addout_25__0})) ;
    FC_nadder_32 loop3_26_fx (.aa ({addout_25__31,addout_25__30,addout_25__29,
                 addout_25__28,addout_25__27,addout_25__26,addout_25__25,
                 addout_25__24,addout_25__23,addout_25__22,addout_25__21,
                 addout_25__20,addout_25__19,addout_25__18,addout_25__17,
                 addout_25__16,addout_25__15,addout_25__14,addout_25__13,
                 addout_25__12,addout_25__11,addout_25__10,addout_25__9,
                 addout_25__8,addout_25__7,addout_25__6,addout_25__5,
                 addout_25__4,addout_25__3,addout_25__2,addout_25__1,
                 addout_25__0}), .bb ({nx5960,nx5972,nx5984,nx5996,nx6010,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_26__31,addout_26__30,addout_26__29
                 ,addout_26__28,addout_26__27,addout_26__26,addout_26__25,
                 addout_26__24,addout_26__23,addout_26__22,addout_26__21,
                 addout_26__20,addout_26__19,addout_26__18,addout_26__17,
                 addout_26__16,addout_26__15,addout_26__14,addout_26__13,
                 addout_26__12,addout_26__11,addout_26__10,addout_26__9,
                 addout_26__8,addout_26__7,addout_26__6,addout_26__5,
                 addout_26__4,addout_26__3,addout_26__2,addout_26__1,
                 addout_26__0})) ;
    FC_nadder_32 loop3_27_fx (.aa ({addout_26__31,addout_26__30,addout_26__29,
                 addout_26__28,addout_26__27,addout_26__26,addout_26__25,
                 addout_26__24,addout_26__23,addout_26__22,addout_26__21,
                 addout_26__20,addout_26__19,addout_26__18,addout_26__17,
                 addout_26__16,addout_26__15,addout_26__14,addout_26__13,
                 addout_26__12,addout_26__11,addout_26__10,addout_26__9,
                 addout_26__8,addout_26__7,addout_26__6,addout_26__5,
                 addout_26__4,addout_26__3,addout_26__2,addout_26__1,
                 addout_26__0}), .bb ({nx5972,nx5984,nx5996,nx6010,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_27__31,addout_27__30,addout_27__29
                 ,addout_27__28,addout_27__27,addout_27__26,addout_27__25,
                 addout_27__24,addout_27__23,addout_27__22,addout_27__21,
                 addout_27__20,addout_27__19,addout_27__18,addout_27__17,
                 addout_27__16,addout_27__15,addout_27__14,addout_27__13,
                 addout_27__12,addout_27__11,addout_27__10,addout_27__9,
                 addout_27__8,addout_27__7,addout_27__6,addout_27__5,
                 addout_27__4,addout_27__3,addout_27__2,addout_27__1,
                 addout_27__0})) ;
    FC_nadder_32 loop3_28_fx (.aa ({addout_27__31,addout_27__30,addout_27__29,
                 addout_27__28,addout_27__27,addout_27__26,addout_27__25,
                 addout_27__24,addout_27__23,addout_27__22,addout_27__21,
                 addout_27__20,addout_27__19,addout_27__18,addout_27__17,
                 addout_27__16,addout_27__15,addout_27__14,addout_27__13,
                 addout_27__12,addout_27__11,addout_27__10,addout_27__9,
                 addout_27__8,addout_27__7,addout_27__6,addout_27__5,
                 addout_27__4,addout_27__3,addout_27__2,addout_27__1,
                 addout_27__0}), .bb ({nx5984,nx5996,nx6010,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_28__31,addout_28__30,addout_28__29
                 ,addout_28__28,addout_28__27,addout_28__26,addout_28__25,
                 addout_28__24,addout_28__23,addout_28__22,addout_28__21,
                 addout_28__20,addout_28__19,addout_28__18,addout_28__17,
                 addout_28__16,addout_28__15,addout_28__14,addout_28__13,
                 addout_28__12,addout_28__11,addout_28__10,addout_28__9,
                 addout_28__8,addout_28__7,addout_28__6,addout_28__5,
                 addout_28__4,addout_28__3,addout_28__2,addout_28__1,
                 addout_28__0})) ;
    FC_nadder_32 loop3_29_fx (.aa ({addout_28__31,addout_28__30,addout_28__29,
                 addout_28__28,addout_28__27,addout_28__26,addout_28__25,
                 addout_28__24,addout_28__23,addout_28__22,addout_28__21,
                 addout_28__20,addout_28__19,addout_28__18,addout_28__17,
                 addout_28__16,addout_28__15,addout_28__14,addout_28__13,
                 addout_28__12,addout_28__11,addout_28__10,addout_28__9,
                 addout_28__8,addout_28__7,addout_28__6,addout_28__5,
                 addout_28__4,addout_28__3,addout_28__2,addout_28__1,
                 addout_28__0}), .bb ({nx5998,nx6012,addout_31__31,addout_31__31
                 ,addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31}), .c_cin (
                 addout_31__31), .ff ({addout_29__31,addout_29__30,addout_29__29
                 ,addout_29__28,addout_29__27,addout_29__26,addout_29__25,
                 addout_29__24,addout_29__23,addout_29__22,addout_29__21,
                 addout_29__20,addout_29__19,addout_29__18,addout_29__17,
                 addout_29__16,addout_29__15,addout_29__14,addout_29__13,
                 addout_29__12,addout_29__11,addout_29__10,addout_29__9,
                 addout_29__8,addout_29__7,addout_29__6,addout_29__5,
                 addout_29__4,addout_29__3,addout_29__2,addout_29__1,
                 addout_29__0})) ;
    FC_nadder_32 loop3_30_fx (.aa ({addout_29__31,addout_29__30,addout_29__29,
                 addout_29__28,addout_29__27,addout_29__26,addout_29__25,
                 addout_29__24,addout_29__23,addout_29__22,addout_29__21,
                 addout_29__20,addout_29__19,addout_29__18,addout_29__17,
                 addout_29__16,addout_29__15,addout_29__14,addout_29__13,
                 addout_29__12,addout_29__11,addout_29__10,addout_29__9,
                 addout_29__8,addout_29__7,addout_29__6,addout_29__5,
                 addout_29__4,addout_29__3,addout_29__2,addout_29__1,
                 addout_29__0}), .bb ({nx6012,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31,addout_31__31,addout_31__31,addout_31__31,
                 addout_31__31}), .c_cin (addout_31__31), .ff ({F[31],F[30],
                 F[29],F[28],F[27],F[26],F[25],F[24],F[23],F[22],F[21],F[20],
                 F[19],F[18],F[17],F[16],F[15],F[14],F[13],F[12],F[11],F[10],
                 F[9],F[8],F[7],F[6],F[5],F[4],F[3],F[2],F[1],F[0]})) ;
    fake_gnd ix5404 (.Y (addout_31__31)) ;
    inv02 ix5769 (.Y (nx5770), .A (nx5768)) ;
    inv02 ix5771 (.Y (nx5772), .A (nx5768)) ;
    inv02 ix5773 (.Y (nx5774), .A (nx5768)) ;
    inv02 ix5775 (.Y (nx5776), .A (nx5768)) ;
    inv02 ix5777 (.Y (nx5778), .A (nx5768)) ;
    inv02 ix5779 (.Y (nx5780), .A (nx5768)) ;
    inv02 ix5783 (.Y (nx5784), .A (nx5782)) ;
    inv02 ix5785 (.Y (nx5786), .A (nx5782)) ;
    inv02 ix5787 (.Y (nx5788), .A (nx5782)) ;
    inv02 ix5789 (.Y (nx5790), .A (nx5782)) ;
    inv02 ix5791 (.Y (nx5792), .A (nx5782)) ;
    inv02 ix5795 (.Y (nx5796), .A (nx5794)) ;
    inv02 ix5797 (.Y (nx5798), .A (nx5794)) ;
    inv02 ix5799 (.Y (nx5800), .A (nx5794)) ;
    inv02 ix5801 (.Y (nx5802), .A (nx5794)) ;
    inv02 ix5803 (.Y (nx5804), .A (nx5794)) ;
    inv02 ix5807 (.Y (nx5808), .A (nx5806)) ;
    inv02 ix5809 (.Y (nx5810), .A (nx5806)) ;
    inv02 ix5811 (.Y (nx5812), .A (nx5806)) ;
    inv02 ix5813 (.Y (nx5814), .A (nx5806)) ;
    inv02 ix5815 (.Y (nx5816), .A (nx5806)) ;
    inv02 ix5819 (.Y (nx5820), .A (nx5818)) ;
    inv02 ix5821 (.Y (nx5822), .A (nx5818)) ;
    inv02 ix5823 (.Y (nx5824), .A (nx5818)) ;
    inv02 ix5825 (.Y (nx5826), .A (nx5818)) ;
    inv02 ix5829 (.Y (nx5830), .A (nx5828)) ;
    inv02 ix5831 (.Y (nx5832), .A (nx5828)) ;
    inv02 ix5833 (.Y (nx5834), .A (nx5828)) ;
    inv02 ix5835 (.Y (nx5836), .A (nx5828)) ;
    inv02 ix5839 (.Y (nx5840), .A (nx5838)) ;
    inv02 ix5841 (.Y (nx5842), .A (nx5838)) ;
    inv02 ix5843 (.Y (nx5844), .A (nx5838)) ;
    inv02 ix5845 (.Y (nx5846), .A (nx5838)) ;
    inv02 ix5849 (.Y (nx5850), .A (nx5848)) ;
    inv02 ix5851 (.Y (nx5852), .A (nx5848)) ;
    inv02 ix5853 (.Y (nx5854), .A (nx5848)) ;
    inv02 ix5857 (.Y (nx5858), .A (nx5856)) ;
    inv02 ix5859 (.Y (nx5860), .A (nx5856)) ;
    inv02 ix5861 (.Y (nx5862), .A (nx5856)) ;
    inv02 ix5865 (.Y (nx5866), .A (nx5864)) ;
    inv02 ix5867 (.Y (nx5868), .A (nx5864)) ;
    inv02 ix5869 (.Y (nx5870), .A (nx5864)) ;
    buf02 ix5871 (.Y (nx5872), .A (op2_10__26)) ;
    buf02 ix5873 (.Y (nx5874), .A (op2_10__26)) ;
    buf02 ix5875 (.Y (nx5876), .A (op2_11__27)) ;
    buf02 ix5877 (.Y (nx5878), .A (op2_11__27)) ;
    buf02 ix5879 (.Y (nx5880), .A (op2_12__28)) ;
    buf02 ix5881 (.Y (nx5882), .A (op2_12__28)) ;
    buf02 ix5883 (.Y (nx5884), .A (op2_14__28)) ;
    buf02 ix5885 (.Y (nx5886), .A (op2_14__28)) ;
    buf02 ix5887 (.Y (nx5888), .A (op2_14__27)) ;
    buf02 ix5889 (.Y (nx5890), .A (op2_14__27)) ;
    buf02 ix5891 (.Y (nx5892), .A (op2_14__26)) ;
    buf02 ix5893 (.Y (nx5894), .A (op2_14__26)) ;
    inv02 ix5897 (.Y (nx5898), .A (nx5896)) ;
    inv02 ix5899 (.Y (nx5900), .A (nx5896)) ;
    inv02 ix5901 (.Y (nx5902), .A (nx5896)) ;
    inv02 ix5905 (.Y (nx5906), .A (nx5904)) ;
    inv02 ix5907 (.Y (nx5908), .A (nx5904)) ;
    inv02 ix5909 (.Y (nx5910), .A (nx5904)) ;
    inv02 ix5913 (.Y (nx5914), .A (nx5912)) ;
    inv02 ix5915 (.Y (nx5916), .A (nx5912)) ;
    inv02 ix5917 (.Y (nx5918), .A (nx5912)) ;
    inv02 ix5921 (.Y (nx5922), .A (nx5920)) ;
    inv02 ix5923 (.Y (nx5924), .A (nx5920)) ;
    inv02 ix5925 (.Y (nx5926), .A (nx5920)) ;
    inv02 ix5927 (.Y (nx5928), .A (nx5920)) ;
    inv02 ix5931 (.Y (nx5932), .A (nx5930)) ;
    inv02 ix5933 (.Y (nx5934), .A (nx5930)) ;
    inv02 ix5935 (.Y (nx5936), .A (nx5930)) ;
    inv02 ix5937 (.Y (nx5938), .A (nx5930)) ;
    inv02 ix5941 (.Y (nx5942), .A (nx5940)) ;
    inv02 ix5943 (.Y (nx5944), .A (nx5940)) ;
    inv02 ix5945 (.Y (nx5946), .A (nx5940)) ;
    inv02 ix5947 (.Y (nx5948), .A (nx5940)) ;
    inv02 ix5951 (.Y (nx5952), .A (nx5950)) ;
    inv02 ix5953 (.Y (nx5954), .A (nx5950)) ;
    inv02 ix5955 (.Y (nx5956), .A (nx5950)) ;
    inv02 ix5957 (.Y (nx5958), .A (nx5950)) ;
    inv02 ix5959 (.Y (nx5960), .A (nx5950)) ;
    inv02 ix5963 (.Y (nx5964), .A (nx5962)) ;
    inv02 ix5965 (.Y (nx5966), .A (nx5962)) ;
    inv02 ix5967 (.Y (nx5968), .A (nx5962)) ;
    inv02 ix5969 (.Y (nx5970), .A (nx5962)) ;
    inv02 ix5971 (.Y (nx5972), .A (nx5962)) ;
    inv02 ix5975 (.Y (nx5976), .A (nx5974)) ;
    inv02 ix5977 (.Y (nx5978), .A (nx5974)) ;
    inv02 ix5979 (.Y (nx5980), .A (nx5974)) ;
    inv02 ix5981 (.Y (nx5982), .A (nx5974)) ;
    inv02 ix5983 (.Y (nx5984), .A (nx5974)) ;
    inv02 ix5987 (.Y (nx5988), .A (nx5986)) ;
    inv02 ix5989 (.Y (nx5990), .A (nx5986)) ;
    inv02 ix5991 (.Y (nx5992), .A (nx5986)) ;
    inv02 ix5993 (.Y (nx5994), .A (nx5986)) ;
    inv02 ix5995 (.Y (nx5996), .A (nx5986)) ;
    inv02 ix5997 (.Y (nx5998), .A (nx5986)) ;
    inv02 ix6001 (.Y (nx6002), .A (nx6000)) ;
    inv02 ix6003 (.Y (nx6004), .A (nx6000)) ;
    inv02 ix6005 (.Y (nx6006), .A (nx6000)) ;
    inv02 ix6007 (.Y (nx6008), .A (nx6000)) ;
    inv02 ix6009 (.Y (nx6010), .A (nx6000)) ;
    inv02 ix6011 (.Y (nx6012), .A (nx6000)) ;
    inv02 ix6015 (.Y (nx6016), .A (nx6014)) ;
    inv02 ix6017 (.Y (nx6018), .A (nx6014)) ;
    inv02 ix6019 (.Y (nx6020), .A (nx6014)) ;
    inv02 ix6021 (.Y (nx6022), .A (nx6014)) ;
    inv02 ix6023 (.Y (nx6024), .A (nx6014)) ;
    inv02 ix6025 (.Y (nx6026), .A (nx6014)) ;
    and02 ix481 (.Y (op1_0), .A0 (nx6346), .A1 (nx6474)) ;
    and02 ix483 (.Y (op1_1), .A0 (nx6338), .A1 (nx6474)) ;
    and02 ix485 (.Y (op1_2), .A0 (nx6330), .A1 (nx6474)) ;
    and02 ix487 (.Y (op1_3), .A0 (nx6322), .A1 (nx6474)) ;
    and02 ix489 (.Y (op1_4), .A0 (nx6314), .A1 (nx6474)) ;
    and02 ix491 (.Y (op1_5), .A0 (nx6306), .A1 (nx6474)) ;
    and02 ix493 (.Y (op1_6), .A0 (nx6298), .A1 (nx6474)) ;
    and02 ix495 (.Y (op1_7), .A0 (nx6290), .A1 (nx6476)) ;
    and02 ix497 (.Y (op1_8), .A0 (nx6282), .A1 (nx6476)) ;
    and02 ix499 (.Y (op1_9), .A0 (nx6274), .A1 (nx6476)) ;
    and02 ix501 (.Y (op1_10), .A0 (nx6266), .A1 (nx6476)) ;
    and02 ix503 (.Y (op1_11), .A0 (nx6258), .A1 (nx6476)) ;
    and02 ix505 (.Y (op1_12), .A0 (nx6250), .A1 (nx6476)) ;
    and02 ix507 (.Y (op1_13), .A0 (nx6242), .A1 (nx6476)) ;
    and02 ix509 (.Y (op1_14), .A0 (nx6234), .A1 (nx6478)) ;
    nand02 ix511 (.Y (nx6014), .A0 (nx6478), .A1 (nx6226)) ;
    nand02 ix1 (.Y (nx6000), .A0 (nx6354), .A1 (nx6346)) ;
    nand02 ix3 (.Y (nx5986), .A0 (nx6354), .A1 (nx6338)) ;
    nand02 ix5 (.Y (nx5974), .A0 (nx6354), .A1 (nx6330)) ;
    nand02 ix7 (.Y (nx5962), .A0 (nx6354), .A1 (nx6322)) ;
    nand02 ix9 (.Y (nx5950), .A0 (nx6354), .A1 (nx6314)) ;
    nand02 ix11 (.Y (nx5940), .A0 (nx6354), .A1 (nx6306)) ;
    nand02 ix13 (.Y (nx5930), .A0 (nx6354), .A1 (nx6298)) ;
    nand02 ix15 (.Y (nx5920), .A0 (nx6356), .A1 (nx6290)) ;
    nand02 ix17 (.Y (nx5912), .A0 (nx6356), .A1 (nx6282)) ;
    nand02 ix19 (.Y (nx5904), .A0 (nx6356), .A1 (nx6274)) ;
    nand02 ix21 (.Y (nx5896), .A0 (nx6356), .A1 (nx6266)) ;
    and02 ix23 (.Y (op2_14__26), .A0 (nx6356), .A1 (nx6258)) ;
    and02 ix25 (.Y (op2_14__27), .A0 (nx6356), .A1 (nx6250)) ;
    and02 ix27 (.Y (op2_14__28), .A0 (nx6356), .A1 (nx6242)) ;
    and02 ix29 (.Y (op2_14__29), .A0 (nx6358), .A1 (nx6234)) ;
    and02 ix31 (.Y (op2_14__30), .A0 (nx6358), .A1 (nx6226)) ;
    and02 ix33 (.Y (op2_13__14), .A0 (nx6362), .A1 (nx6346)) ;
    and02 ix35 (.Y (op2_13__15), .A0 (nx6362), .A1 (nx6338)) ;
    and02 ix37 (.Y (op2_13__16), .A0 (nx6362), .A1 (nx6330)) ;
    and02 ix39 (.Y (op2_13__17), .A0 (nx6362), .A1 (nx6322)) ;
    and02 ix41 (.Y (op2_13__18), .A0 (nx6362), .A1 (nx6314)) ;
    and02 ix43 (.Y (op2_13__19), .A0 (nx6362), .A1 (nx6306)) ;
    and02 ix45 (.Y (op2_13__20), .A0 (nx6362), .A1 (nx6298)) ;
    and02 ix47 (.Y (op2_13__21), .A0 (nx6364), .A1 (nx6290)) ;
    and02 ix49 (.Y (op2_13__22), .A0 (nx6364), .A1 (nx6282)) ;
    and02 ix51 (.Y (op2_13__23), .A0 (nx6364), .A1 (nx6274)) ;
    and02 ix53 (.Y (op2_13__24), .A0 (nx6364), .A1 (nx6266)) ;
    and02 ix55 (.Y (op2_13__25), .A0 (nx6364), .A1 (nx6258)) ;
    and02 ix57 (.Y (op2_13__26), .A0 (nx6364), .A1 (nx6250)) ;
    and02 ix59 (.Y (op2_13__27), .A0 (nx6364), .A1 (nx6242)) ;
    and02 ix61 (.Y (op2_13__28), .A0 (nx6366), .A1 (nx6234)) ;
    and02 ix63 (.Y (op2_13__29), .A0 (nx6366), .A1 (nx6226)) ;
    and02 ix65 (.Y (op2_12__13), .A0 (nx6370), .A1 (nx6346)) ;
    and02 ix67 (.Y (op2_12__14), .A0 (nx6370), .A1 (nx6338)) ;
    and02 ix69 (.Y (op2_12__15), .A0 (nx6370), .A1 (nx6330)) ;
    and02 ix71 (.Y (op2_12__16), .A0 (nx6370), .A1 (nx6322)) ;
    and02 ix73 (.Y (op2_12__17), .A0 (nx6370), .A1 (nx6314)) ;
    and02 ix75 (.Y (op2_12__18), .A0 (nx6370), .A1 (nx6306)) ;
    and02 ix77 (.Y (op2_12__19), .A0 (nx6370), .A1 (nx6298)) ;
    and02 ix79 (.Y (op2_12__20), .A0 (nx6372), .A1 (nx6290)) ;
    and02 ix81 (.Y (op2_12__21), .A0 (nx6372), .A1 (nx6282)) ;
    and02 ix83 (.Y (op2_12__22), .A0 (nx6372), .A1 (nx6274)) ;
    and02 ix85 (.Y (op2_12__23), .A0 (nx6372), .A1 (nx6266)) ;
    and02 ix87 (.Y (op2_12__24), .A0 (nx6372), .A1 (nx6258)) ;
    and02 ix89 (.Y (op2_12__25), .A0 (nx6372), .A1 (nx6250)) ;
    and02 ix91 (.Y (op2_12__26), .A0 (nx6372), .A1 (nx6242)) ;
    and02 ix93 (.Y (op2_12__27), .A0 (nx6374), .A1 (nx6234)) ;
    and02 ix95 (.Y (op2_12__28), .A0 (nx6374), .A1 (nx6226)) ;
    and02 ix97 (.Y (op2_11__12), .A0 (nx6378), .A1 (nx6346)) ;
    and02 ix99 (.Y (op2_11__13), .A0 (nx6378), .A1 (nx6338)) ;
    and02 ix101 (.Y (op2_11__14), .A0 (nx6378), .A1 (nx6330)) ;
    and02 ix103 (.Y (op2_11__15), .A0 (nx6378), .A1 (nx6322)) ;
    and02 ix105 (.Y (op2_11__16), .A0 (nx6378), .A1 (nx6314)) ;
    and02 ix107 (.Y (op2_11__17), .A0 (nx6378), .A1 (nx6306)) ;
    and02 ix109 (.Y (op2_11__18), .A0 (nx6378), .A1 (nx6298)) ;
    and02 ix111 (.Y (op2_11__19), .A0 (nx6380), .A1 (nx6290)) ;
    and02 ix113 (.Y (op2_11__20), .A0 (nx6380), .A1 (nx6282)) ;
    and02 ix115 (.Y (op2_11__21), .A0 (nx6380), .A1 (nx6274)) ;
    and02 ix117 (.Y (op2_11__22), .A0 (nx6380), .A1 (nx6266)) ;
    and02 ix119 (.Y (op2_11__23), .A0 (nx6380), .A1 (nx6258)) ;
    and02 ix121 (.Y (op2_11__24), .A0 (nx6380), .A1 (nx6250)) ;
    and02 ix123 (.Y (op2_11__25), .A0 (nx6380), .A1 (nx6242)) ;
    and02 ix125 (.Y (op2_11__26), .A0 (nx6382), .A1 (nx6234)) ;
    and02 ix127 (.Y (op2_11__27), .A0 (nx6382), .A1 (nx6226)) ;
    and02 ix129 (.Y (op2_10__11), .A0 (nx6386), .A1 (nx6346)) ;
    and02 ix131 (.Y (op2_10__12), .A0 (nx6386), .A1 (nx6338)) ;
    and02 ix133 (.Y (op2_10__13), .A0 (nx6386), .A1 (nx6330)) ;
    and02 ix135 (.Y (op2_10__14), .A0 (nx6386), .A1 (nx6322)) ;
    and02 ix137 (.Y (op2_10__15), .A0 (nx6386), .A1 (nx6314)) ;
    and02 ix139 (.Y (op2_10__16), .A0 (nx6386), .A1 (nx6306)) ;
    and02 ix141 (.Y (op2_10__17), .A0 (nx6386), .A1 (nx6298)) ;
    and02 ix143 (.Y (op2_10__18), .A0 (nx6388), .A1 (nx6290)) ;
    and02 ix145 (.Y (op2_10__19), .A0 (nx6388), .A1 (nx6282)) ;
    and02 ix147 (.Y (op2_10__20), .A0 (nx6388), .A1 (nx6274)) ;
    and02 ix149 (.Y (op2_10__21), .A0 (nx6388), .A1 (nx6266)) ;
    and02 ix151 (.Y (op2_10__22), .A0 (nx6388), .A1 (nx6258)) ;
    and02 ix153 (.Y (op2_10__23), .A0 (nx6388), .A1 (nx6250)) ;
    and02 ix155 (.Y (op2_10__24), .A0 (nx6388), .A1 (nx6242)) ;
    and02 ix157 (.Y (op2_10__25), .A0 (nx6390), .A1 (nx6234)) ;
    and02 ix159 (.Y (op2_10__26), .A0 (nx6390), .A1 (nx6226)) ;
    and02 ix161 (.Y (op2_9__10), .A0 (nx6394), .A1 (nx6346)) ;
    and02 ix163 (.Y (op2_9__11), .A0 (nx6394), .A1 (nx6338)) ;
    and02 ix165 (.Y (op2_9__12), .A0 (nx6394), .A1 (nx6330)) ;
    and02 ix167 (.Y (op2_9__13), .A0 (nx6394), .A1 (nx6322)) ;
    and02 ix169 (.Y (op2_9__14), .A0 (nx6394), .A1 (nx6314)) ;
    and02 ix171 (.Y (op2_9__15), .A0 (nx6394), .A1 (nx6306)) ;
    and02 ix173 (.Y (op2_9__16), .A0 (nx6394), .A1 (nx6298)) ;
    and02 ix175 (.Y (op2_9__17), .A0 (nx6396), .A1 (nx6290)) ;
    and02 ix177 (.Y (op2_9__18), .A0 (nx6396), .A1 (nx6282)) ;
    and02 ix179 (.Y (op2_9__19), .A0 (nx6396), .A1 (nx6274)) ;
    and02 ix181 (.Y (op2_9__20), .A0 (nx6396), .A1 (nx6266)) ;
    and02 ix183 (.Y (op2_9__21), .A0 (nx6396), .A1 (nx6258)) ;
    and02 ix185 (.Y (op2_9__22), .A0 (nx6396), .A1 (nx6250)) ;
    and02 ix187 (.Y (op2_9__23), .A0 (nx6396), .A1 (nx6242)) ;
    and02 ix189 (.Y (op2_9__24), .A0 (nx6398), .A1 (nx6234)) ;
    nand02 ix191 (.Y (nx5864), .A0 (nx6398), .A1 (nx6226)) ;
    and02 ix193 (.Y (op2_8__9), .A0 (nx6402), .A1 (nx6348)) ;
    and02 ix195 (.Y (op2_8__10), .A0 (nx6402), .A1 (nx6340)) ;
    and02 ix197 (.Y (op2_8__11), .A0 (nx6402), .A1 (nx6332)) ;
    and02 ix199 (.Y (op2_8__12), .A0 (nx6402), .A1 (nx6324)) ;
    and02 ix201 (.Y (op2_8__13), .A0 (nx6402), .A1 (nx6316)) ;
    and02 ix203 (.Y (op2_8__14), .A0 (nx6402), .A1 (nx6308)) ;
    and02 ix205 (.Y (op2_8__15), .A0 (nx6402), .A1 (nx6300)) ;
    and02 ix207 (.Y (op2_8__16), .A0 (nx6404), .A1 (nx6292)) ;
    and02 ix209 (.Y (op2_8__17), .A0 (nx6404), .A1 (nx6284)) ;
    and02 ix211 (.Y (op2_8__18), .A0 (nx6404), .A1 (nx6276)) ;
    and02 ix213 (.Y (op2_8__19), .A0 (nx6404), .A1 (nx6268)) ;
    and02 ix215 (.Y (op2_8__20), .A0 (nx6404), .A1 (nx6260)) ;
    and02 ix217 (.Y (op2_8__21), .A0 (nx6404), .A1 (nx6252)) ;
    and02 ix219 (.Y (op2_8__22), .A0 (nx6404), .A1 (nx6244)) ;
    and02 ix221 (.Y (op2_8__23), .A0 (nx6406), .A1 (nx6236)) ;
    nand02 ix223 (.Y (nx5856), .A0 (nx6406), .A1 (nx6228)) ;
    and02 ix225 (.Y (op2_7__8), .A0 (nx6410), .A1 (nx6348)) ;
    and02 ix227 (.Y (op2_7__9), .A0 (nx6410), .A1 (nx6340)) ;
    and02 ix229 (.Y (op2_7__10), .A0 (nx6410), .A1 (nx6332)) ;
    and02 ix231 (.Y (op2_7__11), .A0 (nx6410), .A1 (nx6324)) ;
    and02 ix233 (.Y (op2_7__12), .A0 (nx6410), .A1 (nx6316)) ;
    and02 ix235 (.Y (op2_7__13), .A0 (nx6410), .A1 (nx6308)) ;
    and02 ix237 (.Y (op2_7__14), .A0 (nx6410), .A1 (nx6300)) ;
    and02 ix239 (.Y (op2_7__15), .A0 (nx6412), .A1 (nx6292)) ;
    and02 ix241 (.Y (op2_7__16), .A0 (nx6412), .A1 (nx6284)) ;
    and02 ix243 (.Y (op2_7__17), .A0 (nx6412), .A1 (nx6276)) ;
    and02 ix245 (.Y (op2_7__18), .A0 (nx6412), .A1 (nx6268)) ;
    and02 ix247 (.Y (op2_7__19), .A0 (nx6412), .A1 (nx6260)) ;
    and02 ix249 (.Y (op2_7__20), .A0 (nx6412), .A1 (nx6252)) ;
    and02 ix251 (.Y (op2_7__21), .A0 (nx6412), .A1 (nx6244)) ;
    and02 ix253 (.Y (op2_7__22), .A0 (nx6414), .A1 (nx6236)) ;
    nand02 ix255 (.Y (nx5848), .A0 (nx6414), .A1 (nx6228)) ;
    and02 ix257 (.Y (op2_6__7), .A0 (nx6418), .A1 (nx6348)) ;
    and02 ix259 (.Y (op2_6__8), .A0 (nx6418), .A1 (nx6340)) ;
    and02 ix261 (.Y (op2_6__9), .A0 (nx6418), .A1 (nx6332)) ;
    and02 ix263 (.Y (op2_6__10), .A0 (nx6418), .A1 (nx6324)) ;
    and02 ix265 (.Y (op2_6__11), .A0 (nx6418), .A1 (nx6316)) ;
    and02 ix267 (.Y (op2_6__12), .A0 (nx6418), .A1 (nx6308)) ;
    and02 ix269 (.Y (op2_6__13), .A0 (nx6418), .A1 (nx6300)) ;
    and02 ix271 (.Y (op2_6__14), .A0 (nx6420), .A1 (nx6292)) ;
    and02 ix273 (.Y (op2_6__15), .A0 (nx6420), .A1 (nx6284)) ;
    and02 ix275 (.Y (op2_6__16), .A0 (nx6420), .A1 (nx6276)) ;
    and02 ix277 (.Y (op2_6__17), .A0 (nx6420), .A1 (nx6268)) ;
    and02 ix279 (.Y (op2_6__18), .A0 (nx6420), .A1 (nx6260)) ;
    and02 ix281 (.Y (op2_6__19), .A0 (nx6420), .A1 (nx6252)) ;
    and02 ix283 (.Y (op2_6__20), .A0 (nx6420), .A1 (nx6244)) ;
    and02 ix285 (.Y (op2_6__21), .A0 (nx6422), .A1 (nx6236)) ;
    nand02 ix287 (.Y (nx5838), .A0 (nx6422), .A1 (nx6228)) ;
    and02 ix289 (.Y (op2_5__6), .A0 (nx6426), .A1 (nx6348)) ;
    and02 ix291 (.Y (op2_5__7), .A0 (nx6426), .A1 (nx6340)) ;
    and02 ix293 (.Y (op2_5__8), .A0 (nx6426), .A1 (nx6332)) ;
    and02 ix295 (.Y (op2_5__9), .A0 (nx6426), .A1 (nx6324)) ;
    and02 ix297 (.Y (op2_5__10), .A0 (nx6426), .A1 (nx6316)) ;
    and02 ix299 (.Y (op2_5__11), .A0 (nx6426), .A1 (nx6308)) ;
    and02 ix301 (.Y (op2_5__12), .A0 (nx6426), .A1 (nx6300)) ;
    and02 ix303 (.Y (op2_5__13), .A0 (nx6428), .A1 (nx6292)) ;
    and02 ix305 (.Y (op2_5__14), .A0 (nx6428), .A1 (nx6284)) ;
    and02 ix307 (.Y (op2_5__15), .A0 (nx6428), .A1 (nx6276)) ;
    and02 ix309 (.Y (op2_5__16), .A0 (nx6428), .A1 (nx6268)) ;
    and02 ix311 (.Y (op2_5__17), .A0 (nx6428), .A1 (nx6260)) ;
    and02 ix313 (.Y (op2_5__18), .A0 (nx6428), .A1 (nx6252)) ;
    and02 ix315 (.Y (op2_5__19), .A0 (nx6428), .A1 (nx6244)) ;
    and02 ix317 (.Y (op2_5__20), .A0 (nx6430), .A1 (nx6236)) ;
    nand02 ix319 (.Y (nx5828), .A0 (nx6430), .A1 (nx6228)) ;
    and02 ix321 (.Y (op2_4__5), .A0 (nx6434), .A1 (nx6348)) ;
    and02 ix323 (.Y (op2_4__6), .A0 (nx6434), .A1 (nx6340)) ;
    and02 ix325 (.Y (op2_4__7), .A0 (nx6434), .A1 (nx6332)) ;
    and02 ix327 (.Y (op2_4__8), .A0 (nx6434), .A1 (nx6324)) ;
    and02 ix329 (.Y (op2_4__9), .A0 (nx6434), .A1 (nx6316)) ;
    and02 ix331 (.Y (op2_4__10), .A0 (nx6434), .A1 (nx6308)) ;
    and02 ix333 (.Y (op2_4__11), .A0 (nx6434), .A1 (nx6300)) ;
    and02 ix335 (.Y (op2_4__12), .A0 (nx6436), .A1 (nx6292)) ;
    and02 ix337 (.Y (op2_4__13), .A0 (nx6436), .A1 (nx6284)) ;
    and02 ix339 (.Y (op2_4__14), .A0 (nx6436), .A1 (nx6276)) ;
    and02 ix341 (.Y (op2_4__15), .A0 (nx6436), .A1 (nx6268)) ;
    and02 ix343 (.Y (op2_4__16), .A0 (nx6436), .A1 (nx6260)) ;
    and02 ix345 (.Y (op2_4__17), .A0 (nx6436), .A1 (nx6252)) ;
    and02 ix347 (.Y (op2_4__18), .A0 (nx6436), .A1 (nx6244)) ;
    and02 ix349 (.Y (op2_4__19), .A0 (nx6438), .A1 (nx6236)) ;
    nand02 ix351 (.Y (nx5818), .A0 (nx6438), .A1 (nx6228)) ;
    and02 ix353 (.Y (op2_3__4), .A0 (nx6442), .A1 (nx6348)) ;
    and02 ix355 (.Y (op2_3__5), .A0 (nx6442), .A1 (nx6340)) ;
    and02 ix357 (.Y (op2_3__6), .A0 (nx6442), .A1 (nx6332)) ;
    and02 ix359 (.Y (op2_3__7), .A0 (nx6442), .A1 (nx6324)) ;
    and02 ix361 (.Y (op2_3__8), .A0 (nx6442), .A1 (nx6316)) ;
    and02 ix363 (.Y (op2_3__9), .A0 (nx6442), .A1 (nx6308)) ;
    and02 ix365 (.Y (op2_3__10), .A0 (nx6442), .A1 (nx6300)) ;
    and02 ix367 (.Y (op2_3__11), .A0 (nx6444), .A1 (nx6292)) ;
    and02 ix369 (.Y (op2_3__12), .A0 (nx6444), .A1 (nx6284)) ;
    and02 ix371 (.Y (op2_3__13), .A0 (nx6444), .A1 (nx6276)) ;
    and02 ix373 (.Y (op2_3__14), .A0 (nx6444), .A1 (nx6268)) ;
    and02 ix375 (.Y (op2_3__15), .A0 (nx6444), .A1 (nx6260)) ;
    and02 ix377 (.Y (op2_3__16), .A0 (nx6444), .A1 (nx6252)) ;
    and02 ix379 (.Y (op2_3__17), .A0 (nx6444), .A1 (nx6244)) ;
    and02 ix381 (.Y (op2_3__18), .A0 (nx6446), .A1 (nx6236)) ;
    nand02 ix383 (.Y (nx5806), .A0 (nx6446), .A1 (nx6228)) ;
    and02 ix385 (.Y (op2_2__3), .A0 (nx6450), .A1 (nx6348)) ;
    and02 ix387 (.Y (op2_2__4), .A0 (nx6450), .A1 (nx6340)) ;
    and02 ix389 (.Y (op2_2__5), .A0 (nx6450), .A1 (nx6332)) ;
    and02 ix391 (.Y (op2_2__6), .A0 (nx6450), .A1 (nx6324)) ;
    and02 ix393 (.Y (op2_2__7), .A0 (nx6450), .A1 (nx6316)) ;
    and02 ix395 (.Y (op2_2__8), .A0 (nx6450), .A1 (nx6308)) ;
    and02 ix397 (.Y (op2_2__9), .A0 (nx6450), .A1 (nx6300)) ;
    and02 ix399 (.Y (op2_2__10), .A0 (nx6452), .A1 (nx6292)) ;
    and02 ix401 (.Y (op2_2__11), .A0 (nx6452), .A1 (nx6284)) ;
    and02 ix403 (.Y (op2_2__12), .A0 (nx6452), .A1 (nx6276)) ;
    and02 ix405 (.Y (op2_2__13), .A0 (nx6452), .A1 (nx6268)) ;
    and02 ix407 (.Y (op2_2__14), .A0 (nx6452), .A1 (nx6260)) ;
    and02 ix409 (.Y (op2_2__15), .A0 (nx6452), .A1 (nx6252)) ;
    and02 ix411 (.Y (op2_2__16), .A0 (nx6452), .A1 (nx6244)) ;
    and02 ix413 (.Y (op2_2__17), .A0 (nx6454), .A1 (nx6236)) ;
    nand02 ix415 (.Y (nx5794), .A0 (nx6454), .A1 (nx6228)) ;
    and02 ix417 (.Y (op2_1__2), .A0 (nx6458), .A1 (nx6350)) ;
    and02 ix419 (.Y (op2_1__3), .A0 (nx6458), .A1 (nx6342)) ;
    and02 ix421 (.Y (op2_1__4), .A0 (nx6458), .A1 (nx6334)) ;
    and02 ix423 (.Y (op2_1__5), .A0 (nx6458), .A1 (nx6326)) ;
    and02 ix425 (.Y (op2_1__6), .A0 (nx6458), .A1 (nx6318)) ;
    and02 ix427 (.Y (op2_1__7), .A0 (nx6458), .A1 (nx6310)) ;
    and02 ix429 (.Y (op2_1__8), .A0 (nx6458), .A1 (nx6302)) ;
    and02 ix431 (.Y (op2_1__9), .A0 (nx6460), .A1 (nx6294)) ;
    and02 ix433 (.Y (op2_1__10), .A0 (nx6460), .A1 (nx6286)) ;
    and02 ix435 (.Y (op2_1__11), .A0 (nx6460), .A1 (nx6278)) ;
    and02 ix437 (.Y (op2_1__12), .A0 (nx6460), .A1 (nx6270)) ;
    and02 ix439 (.Y (op2_1__13), .A0 (nx6460), .A1 (nx6262)) ;
    and02 ix441 (.Y (op2_1__14), .A0 (nx6460), .A1 (nx6254)) ;
    and02 ix443 (.Y (op2_1__15), .A0 (nx6460), .A1 (nx6246)) ;
    and02 ix445 (.Y (op2_1__16), .A0 (nx6462), .A1 (nx6238)) ;
    nand02 ix447 (.Y (nx5782), .A0 (nx6462), .A1 (nx6230)) ;
    and02 ix449 (.Y (op2_0__1), .A0 (nx6466), .A1 (nx6350)) ;
    and02 ix451 (.Y (op2_0__2), .A0 (nx6466), .A1 (nx6342)) ;
    and02 ix453 (.Y (op2_0__3), .A0 (nx6466), .A1 (nx6334)) ;
    and02 ix455 (.Y (op2_0__4), .A0 (nx6466), .A1 (nx6326)) ;
    and02 ix457 (.Y (op2_0__5), .A0 (nx6466), .A1 (nx6318)) ;
    and02 ix459 (.Y (op2_0__6), .A0 (nx6466), .A1 (nx6310)) ;
    and02 ix461 (.Y (op2_0__7), .A0 (nx6466), .A1 (nx6302)) ;
    and02 ix463 (.Y (op2_0__8), .A0 (nx6468), .A1 (nx6294)) ;
    and02 ix465 (.Y (op2_0__9), .A0 (nx6468), .A1 (nx6286)) ;
    and02 ix467 (.Y (op2_0__10), .A0 (nx6468), .A1 (nx6278)) ;
    and02 ix469 (.Y (op2_0__11), .A0 (nx6468), .A1 (nx6270)) ;
    and02 ix471 (.Y (op2_0__12), .A0 (nx6468), .A1 (nx6262)) ;
    and02 ix473 (.Y (op2_0__13), .A0 (nx6468), .A1 (nx6254)) ;
    and02 ix475 (.Y (op2_0__14), .A0 (nx6468), .A1 (nx6246)) ;
    and02 ix477 (.Y (op2_0__15), .A0 (nx6470), .A1 (nx6238)) ;
    nand02 ix479 (.Y (nx5768), .A0 (nx6470), .A1 (nx6230)) ;
    inv01 ix6223 (.Y (nx6224), .A (A[15])) ;
    inv02 ix6225 (.Y (nx6226), .A (nx6224)) ;
    inv02 ix6227 (.Y (nx6228), .A (nx6224)) ;
    inv02 ix6229 (.Y (nx6230), .A (nx6224)) ;
    inv01 ix6231 (.Y (nx6232), .A (A[14])) ;
    inv02 ix6233 (.Y (nx6234), .A (nx6232)) ;
    inv02 ix6235 (.Y (nx6236), .A (nx6232)) ;
    inv02 ix6237 (.Y (nx6238), .A (nx6232)) ;
    inv01 ix6239 (.Y (nx6240), .A (A[13])) ;
    inv02 ix6241 (.Y (nx6242), .A (nx6240)) ;
    inv02 ix6243 (.Y (nx6244), .A (nx6240)) ;
    inv02 ix6245 (.Y (nx6246), .A (nx6240)) ;
    inv01 ix6247 (.Y (nx6248), .A (A[12])) ;
    inv02 ix6249 (.Y (nx6250), .A (nx6248)) ;
    inv02 ix6251 (.Y (nx6252), .A (nx6248)) ;
    inv02 ix6253 (.Y (nx6254), .A (nx6248)) ;
    inv01 ix6255 (.Y (nx6256), .A (A[11])) ;
    inv02 ix6257 (.Y (nx6258), .A (nx6256)) ;
    inv02 ix6259 (.Y (nx6260), .A (nx6256)) ;
    inv02 ix6261 (.Y (nx6262), .A (nx6256)) ;
    inv01 ix6263 (.Y (nx6264), .A (A[10])) ;
    inv02 ix6265 (.Y (nx6266), .A (nx6264)) ;
    inv02 ix6267 (.Y (nx6268), .A (nx6264)) ;
    inv02 ix6269 (.Y (nx6270), .A (nx6264)) ;
    inv01 ix6271 (.Y (nx6272), .A (A[9])) ;
    inv02 ix6273 (.Y (nx6274), .A (nx6272)) ;
    inv02 ix6275 (.Y (nx6276), .A (nx6272)) ;
    inv02 ix6277 (.Y (nx6278), .A (nx6272)) ;
    inv01 ix6279 (.Y (nx6280), .A (A[8])) ;
    inv02 ix6281 (.Y (nx6282), .A (nx6280)) ;
    inv02 ix6283 (.Y (nx6284), .A (nx6280)) ;
    inv02 ix6285 (.Y (nx6286), .A (nx6280)) ;
    inv01 ix6287 (.Y (nx6288), .A (A[7])) ;
    inv02 ix6289 (.Y (nx6290), .A (nx6288)) ;
    inv02 ix6291 (.Y (nx6292), .A (nx6288)) ;
    inv02 ix6293 (.Y (nx6294), .A (nx6288)) ;
    inv01 ix6295 (.Y (nx6296), .A (A[6])) ;
    inv02 ix6297 (.Y (nx6298), .A (nx6296)) ;
    inv02 ix6299 (.Y (nx6300), .A (nx6296)) ;
    inv02 ix6301 (.Y (nx6302), .A (nx6296)) ;
    inv01 ix6303 (.Y (nx6304), .A (A[5])) ;
    inv02 ix6305 (.Y (nx6306), .A (nx6304)) ;
    inv02 ix6307 (.Y (nx6308), .A (nx6304)) ;
    inv02 ix6309 (.Y (nx6310), .A (nx6304)) ;
    inv01 ix6311 (.Y (nx6312), .A (A[4])) ;
    inv02 ix6313 (.Y (nx6314), .A (nx6312)) ;
    inv02 ix6315 (.Y (nx6316), .A (nx6312)) ;
    inv02 ix6317 (.Y (nx6318), .A (nx6312)) ;
    inv01 ix6319 (.Y (nx6320), .A (A[3])) ;
    inv02 ix6321 (.Y (nx6322), .A (nx6320)) ;
    inv02 ix6323 (.Y (nx6324), .A (nx6320)) ;
    inv02 ix6325 (.Y (nx6326), .A (nx6320)) ;
    inv01 ix6327 (.Y (nx6328), .A (A[2])) ;
    inv02 ix6329 (.Y (nx6330), .A (nx6328)) ;
    inv02 ix6331 (.Y (nx6332), .A (nx6328)) ;
    inv02 ix6333 (.Y (nx6334), .A (nx6328)) ;
    inv01 ix6335 (.Y (nx6336), .A (A[1])) ;
    inv02 ix6337 (.Y (nx6338), .A (nx6336)) ;
    inv02 ix6339 (.Y (nx6340), .A (nx6336)) ;
    inv02 ix6341 (.Y (nx6342), .A (nx6336)) ;
    inv01 ix6343 (.Y (nx6344), .A (A[0])) ;
    inv02 ix6345 (.Y (nx6346), .A (nx6344)) ;
    inv02 ix6347 (.Y (nx6348), .A (nx6344)) ;
    inv02 ix6349 (.Y (nx6350), .A (nx6344)) ;
    inv01 ix6351 (.Y (nx6352), .A (B[15])) ;
    inv01 ix6353 (.Y (nx6354), .A (nx6352)) ;
    inv01 ix6355 (.Y (nx6356), .A (nx6352)) ;
    inv01 ix6357 (.Y (nx6358), .A (nx6352)) ;
    inv01 ix6359 (.Y (nx6360), .A (B[14])) ;
    inv01 ix6361 (.Y (nx6362), .A (nx6360)) ;
    inv01 ix6363 (.Y (nx6364), .A (nx6360)) ;
    inv01 ix6365 (.Y (nx6366), .A (nx6360)) ;
    inv01 ix6367 (.Y (nx6368), .A (B[13])) ;
    inv01 ix6369 (.Y (nx6370), .A (nx6368)) ;
    inv01 ix6371 (.Y (nx6372), .A (nx6368)) ;
    inv01 ix6373 (.Y (nx6374), .A (nx6368)) ;
    inv01 ix6375 (.Y (nx6376), .A (B[12])) ;
    inv01 ix6377 (.Y (nx6378), .A (nx6376)) ;
    inv01 ix6379 (.Y (nx6380), .A (nx6376)) ;
    inv01 ix6381 (.Y (nx6382), .A (nx6376)) ;
    inv01 ix6383 (.Y (nx6384), .A (B[11])) ;
    inv01 ix6385 (.Y (nx6386), .A (nx6384)) ;
    inv01 ix6387 (.Y (nx6388), .A (nx6384)) ;
    inv01 ix6389 (.Y (nx6390), .A (nx6384)) ;
    inv01 ix6391 (.Y (nx6392), .A (B[10])) ;
    inv01 ix6393 (.Y (nx6394), .A (nx6392)) ;
    inv01 ix6395 (.Y (nx6396), .A (nx6392)) ;
    inv01 ix6397 (.Y (nx6398), .A (nx6392)) ;
    inv01 ix6399 (.Y (nx6400), .A (B[9])) ;
    inv01 ix6401 (.Y (nx6402), .A (nx6400)) ;
    inv01 ix6403 (.Y (nx6404), .A (nx6400)) ;
    inv01 ix6405 (.Y (nx6406), .A (nx6400)) ;
    inv01 ix6407 (.Y (nx6408), .A (B[8])) ;
    inv01 ix6409 (.Y (nx6410), .A (nx6408)) ;
    inv01 ix6411 (.Y (nx6412), .A (nx6408)) ;
    inv01 ix6413 (.Y (nx6414), .A (nx6408)) ;
    inv01 ix6415 (.Y (nx6416), .A (B[7])) ;
    inv01 ix6417 (.Y (nx6418), .A (nx6416)) ;
    inv01 ix6419 (.Y (nx6420), .A (nx6416)) ;
    inv01 ix6421 (.Y (nx6422), .A (nx6416)) ;
    inv01 ix6423 (.Y (nx6424), .A (B[6])) ;
    inv01 ix6425 (.Y (nx6426), .A (nx6424)) ;
    inv01 ix6427 (.Y (nx6428), .A (nx6424)) ;
    inv01 ix6429 (.Y (nx6430), .A (nx6424)) ;
    inv01 ix6431 (.Y (nx6432), .A (B[5])) ;
    inv01 ix6433 (.Y (nx6434), .A (nx6432)) ;
    inv01 ix6435 (.Y (nx6436), .A (nx6432)) ;
    inv01 ix6437 (.Y (nx6438), .A (nx6432)) ;
    inv01 ix6439 (.Y (nx6440), .A (B[4])) ;
    inv01 ix6441 (.Y (nx6442), .A (nx6440)) ;
    inv01 ix6443 (.Y (nx6444), .A (nx6440)) ;
    inv01 ix6445 (.Y (nx6446), .A (nx6440)) ;
    inv01 ix6447 (.Y (nx6448), .A (B[3])) ;
    inv01 ix6449 (.Y (nx6450), .A (nx6448)) ;
    inv01 ix6451 (.Y (nx6452), .A (nx6448)) ;
    inv01 ix6453 (.Y (nx6454), .A (nx6448)) ;
    inv01 ix6455 (.Y (nx6456), .A (B[2])) ;
    inv01 ix6457 (.Y (nx6458), .A (nx6456)) ;
    inv01 ix6459 (.Y (nx6460), .A (nx6456)) ;
    inv01 ix6461 (.Y (nx6462), .A (nx6456)) ;
    inv01 ix6463 (.Y (nx6464), .A (B[1])) ;
    inv01 ix6465 (.Y (nx6466), .A (nx6464)) ;
    inv01 ix6467 (.Y (nx6468), .A (nx6464)) ;
    inv01 ix6469 (.Y (nx6470), .A (nx6464)) ;
    inv01 ix6471 (.Y (nx6472), .A (B[0])) ;
    inv02 ix6473 (.Y (nx6474), .A (nx6472)) ;
    inv02 ix6475 (.Y (nx6476), .A (nx6472)) ;
    inv02 ix6477 (.Y (nx6478), .A (nx6472)) ;
    buf02 ix6479 (.Y (nx6480), .A (op2_13__29)) ;
    buf02 ix6481 (.Y (nx6482), .A (op2_14__30)) ;
    buf02 ix6483 (.Y (nx6484), .A (op2_14__29)) ;
endmodule


module FC_nadder_32 ( aa, bb, c_cin, ff ) ;

    input [31:0]aa ;
    input [31:0]bb ;
    input c_cin ;
    output [31:0]ff ;

    wire temp_30, temp_29, temp_28, temp_27, temp_26, temp_25, temp_24, temp_23, 
         temp_22, temp_21, temp_20, temp_19, temp_18, temp_17, temp_16, temp_15, 
         temp_14, temp_13, temp_12, temp_11, temp_10, temp_9, temp_8, temp_7, 
         temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0;
    wire [0:0] \$dummy ;




    FC_adder f0 (.a (aa[0]), .b (bb[0]), .cin (c_cin), .f (ff[0]), .cout (temp_0
             )) ;
    FC_adder loop1_1_fx (.a (aa[1]), .b (bb[1]), .cin (temp_0), .f (ff[1]), .cout (
             temp_1)) ;
    FC_adder loop1_2_fx (.a (aa[2]), .b (bb[2]), .cin (temp_1), .f (ff[2]), .cout (
             temp_2)) ;
    FC_adder loop1_3_fx (.a (aa[3]), .b (bb[3]), .cin (temp_2), .f (ff[3]), .cout (
             temp_3)) ;
    FC_adder loop1_4_fx (.a (aa[4]), .b (bb[4]), .cin (temp_3), .f (ff[4]), .cout (
             temp_4)) ;
    FC_adder loop1_5_fx (.a (aa[5]), .b (bb[5]), .cin (temp_4), .f (ff[5]), .cout (
             temp_5)) ;
    FC_adder loop1_6_fx (.a (aa[6]), .b (bb[6]), .cin (temp_5), .f (ff[6]), .cout (
             temp_6)) ;
    FC_adder loop1_7_fx (.a (aa[7]), .b (bb[7]), .cin (temp_6), .f (ff[7]), .cout (
             temp_7)) ;
    FC_adder loop1_8_fx (.a (aa[8]), .b (bb[8]), .cin (temp_7), .f (ff[8]), .cout (
             temp_8)) ;
    FC_adder loop1_9_fx (.a (aa[9]), .b (bb[9]), .cin (temp_8), .f (ff[9]), .cout (
             temp_9)) ;
    FC_adder loop1_10_fx (.a (aa[10]), .b (bb[10]), .cin (temp_9), .f (ff[10]), 
             .cout (temp_10)) ;
    FC_adder loop1_11_fx (.a (aa[11]), .b (bb[11]), .cin (temp_10), .f (ff[11])
             , .cout (temp_11)) ;
    FC_adder loop1_12_fx (.a (aa[12]), .b (bb[12]), .cin (temp_11), .f (ff[12])
             , .cout (temp_12)) ;
    FC_adder loop1_13_fx (.a (aa[13]), .b (bb[13]), .cin (temp_12), .f (ff[13])
             , .cout (temp_13)) ;
    FC_adder loop1_14_fx (.a (aa[14]), .b (bb[14]), .cin (temp_13), .f (ff[14])
             , .cout (temp_14)) ;
    FC_adder loop1_15_fx (.a (aa[15]), .b (bb[15]), .cin (temp_14), .f (ff[15])
             , .cout (temp_15)) ;
    FC_adder loop1_16_fx (.a (aa[16]), .b (bb[16]), .cin (temp_15), .f (ff[16])
             , .cout (temp_16)) ;
    FC_adder loop1_17_fx (.a (aa[17]), .b (bb[17]), .cin (temp_16), .f (ff[17])
             , .cout (temp_17)) ;
    FC_adder loop1_18_fx (.a (aa[18]), .b (bb[18]), .cin (temp_17), .f (ff[18])
             , .cout (temp_18)) ;
    FC_adder loop1_19_fx (.a (aa[19]), .b (bb[19]), .cin (temp_18), .f (ff[19])
             , .cout (temp_19)) ;
    FC_adder loop1_20_fx (.a (aa[20]), .b (bb[20]), .cin (temp_19), .f (ff[20])
             , .cout (temp_20)) ;
    FC_adder loop1_21_fx (.a (aa[21]), .b (bb[21]), .cin (temp_20), .f (ff[21])
             , .cout (temp_21)) ;
    FC_adder loop1_22_fx (.a (aa[22]), .b (bb[22]), .cin (temp_21), .f (ff[22])
             , .cout (temp_22)) ;
    FC_adder loop1_23_fx (.a (aa[23]), .b (bb[23]), .cin (temp_22), .f (ff[23])
             , .cout (temp_23)) ;
    FC_adder loop1_24_fx (.a (aa[24]), .b (bb[24]), .cin (temp_23), .f (ff[24])
             , .cout (temp_24)) ;
    FC_adder loop1_25_fx (.a (aa[25]), .b (bb[25]), .cin (temp_24), .f (ff[25])
             , .cout (temp_25)) ;
    FC_adder loop1_26_fx (.a (aa[26]), .b (bb[26]), .cin (temp_25), .f (ff[26])
             , .cout (temp_26)) ;
    FC_adder loop1_27_fx (.a (aa[27]), .b (bb[27]), .cin (temp_26), .f (ff[27])
             , .cout (temp_27)) ;
    FC_adder loop1_28_fx (.a (aa[28]), .b (bb[28]), .cin (temp_27), .f (ff[28])
             , .cout (temp_28)) ;
    FC_adder loop1_29_fx (.a (aa[29]), .b (bb[29]), .cin (temp_28), .f (ff[29])
             , .cout (temp_29)) ;
    FC_adder loop1_30_fx (.a (aa[30]), .b (bb[30]), .cin (temp_29), .f (ff[30])
             , .cout (temp_30)) ;
    FC_adder loop1_31_fx (.a (aa[31]), .b (bb[31]), .cin (temp_30), .f (ff[31])
             , .cout (\$dummy [0])) ;
endmodule


module FC_adder ( a, b, cin, f, cout ) ;

    input a ;
    input b ;
    input cin ;
    output f ;
    output cout ;

    wire nx0, nx69;



    ao22 ix7 (.Y (cout), .A0 (b), .A1 (a), .B0 (cin), .B1 (nx0)) ;
    xnor2 ix9 (.Y (f), .A0 (nx69), .A1 (cin)) ;
    xnor2 ix70 (.Y (nx69), .A0 (a), .A1 (b)) ;
    inv01 ix1 (.Y (nx0), .A (nx69)) ;
endmodule


module ReadImage ( WI, current_state, CLK, RST, ACK, ImgAddress, ImgWidth, DATA, 
                   OutputImg0, OutputImg1, OutputImg2, OutputImg3, OutputImg4, 
                   OutputImg5, ImgCounterOuput, ImgAddToDma, UpdatedAddress, 
                   ImgIndic, ImgEn, dontTrust ) ;

    input WI ;
    input [14:0]current_state ;
    input CLK ;
    input RST ;
    input ACK ;
    input [12:0]ImgAddress ;
    input [15:0]ImgWidth ;
    input [447:0]DATA ;
    output [447:0]OutputImg0 ;
    output [447:0]OutputImg1 ;
    output [447:0]OutputImg2 ;
    output [447:0]OutputImg3 ;
    output [447:0]OutputImg4 ;
    output [447:0]OutputImg5 ;
    output [2:0]ImgCounterOuput ;
    output [12:0]ImgAddToDma ;
    output [12:0]UpdatedAddress ;
    output [0:0]ImgIndic ;
    output [5:0]ImgEn ;
    input dontTrust ;

    wire newAdd16_12, newAdd16_11, newAdd16_10, newAdd16_9, newAdd16_8, 
         newAdd16_7, newAdd16_6, newAdd16_5, newAdd16_4, newAdd16_3, newAdd16_2, 
         newAdd16_1, newAdd16_0, DFFCLK, DecOutput_5, DecOutput_4, DecOutput_3, 
         DecOutput_2, DecOutput_1, DecOutput_0, ImgReg0IN_447, ImgReg0IN_446, 
         ImgReg0IN_445, ImgReg0IN_444, ImgReg0IN_443, ImgReg0IN_442, 
         ImgReg0IN_441, ImgReg0IN_440, ImgReg0IN_439, ImgReg0IN_438, 
         ImgReg0IN_437, ImgReg0IN_436, ImgReg0IN_435, ImgReg0IN_434, 
         ImgReg0IN_433, ImgReg0IN_432, ImgReg0IN_431, ImgReg0IN_430, 
         ImgReg0IN_429, ImgReg0IN_428, ImgReg0IN_427, ImgReg0IN_426, 
         ImgReg0IN_425, ImgReg0IN_424, ImgReg0IN_423, ImgReg0IN_422, 
         ImgReg0IN_421, ImgReg0IN_420, ImgReg0IN_419, ImgReg0IN_418, 
         ImgReg0IN_417, ImgReg0IN_416, ImgReg0IN_415, ImgReg0IN_414, 
         ImgReg0IN_413, ImgReg0IN_412, ImgReg0IN_411, ImgReg0IN_410, 
         ImgReg0IN_409, ImgReg0IN_408, ImgReg0IN_407, ImgReg0IN_406, 
         ImgReg0IN_405, ImgReg0IN_404, ImgReg0IN_403, ImgReg0IN_402, 
         ImgReg0IN_401, ImgReg0IN_400, ImgReg0IN_399, ImgReg0IN_398, 
         ImgReg0IN_397, ImgReg0IN_396, ImgReg0IN_395, ImgReg0IN_394, 
         ImgReg0IN_393, ImgReg0IN_392, ImgReg0IN_391, ImgReg0IN_390, 
         ImgReg0IN_389, ImgReg0IN_388, ImgReg0IN_387, ImgReg0IN_386, 
         ImgReg0IN_385, ImgReg0IN_384, ImgReg0IN_383, ImgReg0IN_382, 
         ImgReg0IN_381, ImgReg0IN_380, ImgReg0IN_379, ImgReg0IN_378, 
         ImgReg0IN_377, ImgReg0IN_376, ImgReg0IN_375, ImgReg0IN_374, 
         ImgReg0IN_373, ImgReg0IN_372, ImgReg0IN_371, ImgReg0IN_370, 
         ImgReg0IN_369, ImgReg0IN_368, ImgReg0IN_367, ImgReg0IN_366, 
         ImgReg0IN_365, ImgReg0IN_364, ImgReg0IN_363, ImgReg0IN_362, 
         ImgReg0IN_361, ImgReg0IN_360, ImgReg0IN_359, ImgReg0IN_358, 
         ImgReg0IN_357, ImgReg0IN_356, ImgReg0IN_355, ImgReg0IN_354, 
         ImgReg0IN_353, ImgReg0IN_352, ImgReg0IN_351, ImgReg0IN_350, 
         ImgReg0IN_349, ImgReg0IN_348, ImgReg0IN_347, ImgReg0IN_346, 
         ImgReg0IN_345, ImgReg0IN_344, ImgReg0IN_343, ImgReg0IN_342, 
         ImgReg0IN_341, ImgReg0IN_340, ImgReg0IN_339, ImgReg0IN_338, 
         ImgReg0IN_337, ImgReg0IN_336, ImgReg0IN_335, ImgReg0IN_334, 
         ImgReg0IN_333, ImgReg0IN_332, ImgReg0IN_331, ImgReg0IN_330, 
         ImgReg0IN_329, ImgReg0IN_328, ImgReg0IN_327, ImgReg0IN_326, 
         ImgReg0IN_325, ImgReg0IN_324, ImgReg0IN_323, ImgReg0IN_322, 
         ImgReg0IN_321, ImgReg0IN_320, ImgReg0IN_319, ImgReg0IN_318, 
         ImgReg0IN_317, ImgReg0IN_316, ImgReg0IN_315, ImgReg0IN_314, 
         ImgReg0IN_313, ImgReg0IN_312, ImgReg0IN_311, ImgReg0IN_310, 
         ImgReg0IN_309, ImgReg0IN_308, ImgReg0IN_307, ImgReg0IN_306, 
         ImgReg0IN_305, ImgReg0IN_304, ImgReg0IN_303, ImgReg0IN_302, 
         ImgReg0IN_301, ImgReg0IN_300, ImgReg0IN_299, ImgReg0IN_298, 
         ImgReg0IN_297, ImgReg0IN_296, ImgReg0IN_295, ImgReg0IN_294, 
         ImgReg0IN_293, ImgReg0IN_292, ImgReg0IN_291, ImgReg0IN_290, 
         ImgReg0IN_289, ImgReg0IN_288, ImgReg0IN_287, ImgReg0IN_286, 
         ImgReg0IN_285, ImgReg0IN_284, ImgReg0IN_283, ImgReg0IN_282, 
         ImgReg0IN_281, ImgReg0IN_280, ImgReg0IN_279, ImgReg0IN_278, 
         ImgReg0IN_277, ImgReg0IN_276, ImgReg0IN_275, ImgReg0IN_274, 
         ImgReg0IN_273, ImgReg0IN_272, ImgReg0IN_271, ImgReg0IN_270, 
         ImgReg0IN_269, ImgReg0IN_268, ImgReg0IN_267, ImgReg0IN_266, 
         ImgReg0IN_265, ImgReg0IN_264, ImgReg0IN_263, ImgReg0IN_262, 
         ImgReg0IN_261, ImgReg0IN_260, ImgReg0IN_259, ImgReg0IN_258, 
         ImgReg0IN_257, ImgReg0IN_256, ImgReg0IN_255, ImgReg0IN_254, 
         ImgReg0IN_253, ImgReg0IN_252, ImgReg0IN_251, ImgReg0IN_250, 
         ImgReg0IN_249, ImgReg0IN_248, ImgReg0IN_247, ImgReg0IN_246, 
         ImgReg0IN_245, ImgReg0IN_244, ImgReg0IN_243, ImgReg0IN_242, 
         ImgReg0IN_241, ImgReg0IN_240, ImgReg0IN_239, ImgReg0IN_238, 
         ImgReg0IN_237, ImgReg0IN_236, ImgReg0IN_235, ImgReg0IN_234, 
         ImgReg0IN_233, ImgReg0IN_232, ImgReg0IN_231, ImgReg0IN_230, 
         ImgReg0IN_229, ImgReg0IN_228, ImgReg0IN_227, ImgReg0IN_226, 
         ImgReg0IN_225, ImgReg0IN_224, ImgReg0IN_223, ImgReg0IN_222, 
         ImgReg0IN_221, ImgReg0IN_220, ImgReg0IN_219, ImgReg0IN_218, 
         ImgReg0IN_217, ImgReg0IN_216, ImgReg0IN_215, ImgReg0IN_214, 
         ImgReg0IN_213, ImgReg0IN_212, ImgReg0IN_211, ImgReg0IN_210, 
         ImgReg0IN_209, ImgReg0IN_208, ImgReg0IN_207, ImgReg0IN_206, 
         ImgReg0IN_205, ImgReg0IN_204, ImgReg0IN_203, ImgReg0IN_202, 
         ImgReg0IN_201, ImgReg0IN_200, ImgReg0IN_199, ImgReg0IN_198, 
         ImgReg0IN_197, ImgReg0IN_196, ImgReg0IN_195, ImgReg0IN_194, 
         ImgReg0IN_193, ImgReg0IN_192, ImgReg0IN_191, ImgReg0IN_190, 
         ImgReg0IN_189, ImgReg0IN_188, ImgReg0IN_187, ImgReg0IN_186, 
         ImgReg0IN_185, ImgReg0IN_184, ImgReg0IN_183, ImgReg0IN_182, 
         ImgReg0IN_181, ImgReg0IN_180, ImgReg0IN_179, ImgReg0IN_178, 
         ImgReg0IN_177, ImgReg0IN_176, ImgReg0IN_175, ImgReg0IN_174, 
         ImgReg0IN_173, ImgReg0IN_172, ImgReg0IN_171, ImgReg0IN_170, 
         ImgReg0IN_169, ImgReg0IN_168, ImgReg0IN_167, ImgReg0IN_166, 
         ImgReg0IN_165, ImgReg0IN_164, ImgReg0IN_163, ImgReg0IN_162, 
         ImgReg0IN_161, ImgReg0IN_160, ImgReg0IN_159, ImgReg0IN_158, 
         ImgReg0IN_157, ImgReg0IN_156, ImgReg0IN_155, ImgReg0IN_154, 
         ImgReg0IN_153, ImgReg0IN_152, ImgReg0IN_151, ImgReg0IN_150, 
         ImgReg0IN_149, ImgReg0IN_148, ImgReg0IN_147, ImgReg0IN_146, 
         ImgReg0IN_145, ImgReg0IN_144, ImgReg0IN_143, ImgReg0IN_142, 
         ImgReg0IN_141, ImgReg0IN_140, ImgReg0IN_139, ImgReg0IN_138, 
         ImgReg0IN_137, ImgReg0IN_136, ImgReg0IN_135, ImgReg0IN_134, 
         ImgReg0IN_133, ImgReg0IN_132, ImgReg0IN_131, ImgReg0IN_130, 
         ImgReg0IN_129, ImgReg0IN_128, ImgReg0IN_127, ImgReg0IN_126, 
         ImgReg0IN_125, ImgReg0IN_124, ImgReg0IN_123, ImgReg0IN_122, 
         ImgReg0IN_121, ImgReg0IN_120, ImgReg0IN_119, ImgReg0IN_118, 
         ImgReg0IN_117, ImgReg0IN_116, ImgReg0IN_115, ImgReg0IN_114, 
         ImgReg0IN_113, ImgReg0IN_112, ImgReg0IN_111, ImgReg0IN_110, 
         ImgReg0IN_109, ImgReg0IN_108, ImgReg0IN_107, ImgReg0IN_106, 
         ImgReg0IN_105, ImgReg0IN_104, ImgReg0IN_103, ImgReg0IN_102, 
         ImgReg0IN_101, ImgReg0IN_100, ImgReg0IN_99, ImgReg0IN_98, ImgReg0IN_97, 
         ImgReg0IN_96, ImgReg0IN_95, ImgReg0IN_94, ImgReg0IN_93, ImgReg0IN_92, 
         ImgReg0IN_91, ImgReg0IN_90, ImgReg0IN_89, ImgReg0IN_88, ImgReg0IN_87, 
         ImgReg0IN_86, ImgReg0IN_85, ImgReg0IN_84, ImgReg0IN_83, ImgReg0IN_82, 
         ImgReg0IN_81, ImgReg0IN_80, ImgReg0IN_79, ImgReg0IN_78, ImgReg0IN_77, 
         ImgReg0IN_76, ImgReg0IN_75, ImgReg0IN_74, ImgReg0IN_73, ImgReg0IN_72, 
         ImgReg0IN_71, ImgReg0IN_70, ImgReg0IN_69, ImgReg0IN_68, ImgReg0IN_67, 
         ImgReg0IN_66, ImgReg0IN_65, ImgReg0IN_64, ImgReg0IN_63, ImgReg0IN_62, 
         ImgReg0IN_61, ImgReg0IN_60, ImgReg0IN_59, ImgReg0IN_58, ImgReg0IN_57, 
         ImgReg0IN_56, ImgReg0IN_55, ImgReg0IN_54, ImgReg0IN_53, ImgReg0IN_52, 
         ImgReg0IN_51, ImgReg0IN_50, ImgReg0IN_49, ImgReg0IN_48, ImgReg0IN_47, 
         ImgReg0IN_46, ImgReg0IN_45, ImgReg0IN_44, ImgReg0IN_43, ImgReg0IN_42, 
         ImgReg0IN_41, ImgReg0IN_40, ImgReg0IN_39, ImgReg0IN_38, ImgReg0IN_37, 
         ImgReg0IN_36, ImgReg0IN_35, ImgReg0IN_34, ImgReg0IN_33, ImgReg0IN_32, 
         ImgReg0IN_31, ImgReg0IN_30, ImgReg0IN_29, ImgReg0IN_28, ImgReg0IN_27, 
         ImgReg0IN_26, ImgReg0IN_25, ImgReg0IN_24, ImgReg0IN_23, ImgReg0IN_22, 
         ImgReg0IN_21, ImgReg0IN_20, ImgReg0IN_19, ImgReg0IN_18, ImgReg0IN_17, 
         ImgReg0IN_16, ImgReg0IN_15, ImgReg0IN_14, ImgReg0IN_13, ImgReg0IN_12, 
         ImgReg0IN_11, ImgReg0IN_10, ImgReg0IN_9, ImgReg0IN_8, ImgReg0IN_7, 
         ImgReg0IN_6, ImgReg0IN_5, ImgReg0IN_4, ImgReg0IN_3, ImgReg0IN_2, 
         ImgReg0IN_1, ImgReg0IN_0, ImgReg1IN_447, ImgReg1IN_446, ImgReg1IN_445, 
         ImgReg1IN_444, ImgReg1IN_443, ImgReg1IN_442, ImgReg1IN_441, 
         ImgReg1IN_440, ImgReg1IN_439, ImgReg1IN_438, ImgReg1IN_437, 
         ImgReg1IN_436, ImgReg1IN_435, ImgReg1IN_434, ImgReg1IN_433, 
         ImgReg1IN_432, ImgReg1IN_431, ImgReg1IN_430, ImgReg1IN_429, 
         ImgReg1IN_428, ImgReg1IN_427, ImgReg1IN_426, ImgReg1IN_425, 
         ImgReg1IN_424, ImgReg1IN_423, ImgReg1IN_422, ImgReg1IN_421, 
         ImgReg1IN_420, ImgReg1IN_419, ImgReg1IN_418, ImgReg1IN_417, 
         ImgReg1IN_416, ImgReg1IN_415, ImgReg1IN_414, ImgReg1IN_413, 
         ImgReg1IN_412, ImgReg1IN_411, ImgReg1IN_410, ImgReg1IN_409, 
         ImgReg1IN_408, ImgReg1IN_407, ImgReg1IN_406, ImgReg1IN_405, 
         ImgReg1IN_404, ImgReg1IN_403, ImgReg1IN_402, ImgReg1IN_401, 
         ImgReg1IN_400, ImgReg1IN_399, ImgReg1IN_398, ImgReg1IN_397, 
         ImgReg1IN_396, ImgReg1IN_395, ImgReg1IN_394, ImgReg1IN_393, 
         ImgReg1IN_392, ImgReg1IN_391, ImgReg1IN_390, ImgReg1IN_389, 
         ImgReg1IN_388, ImgReg1IN_387, ImgReg1IN_386, ImgReg1IN_385, 
         ImgReg1IN_384, ImgReg1IN_383, ImgReg1IN_382, ImgReg1IN_381, 
         ImgReg1IN_380, ImgReg1IN_379, ImgReg1IN_378, ImgReg1IN_377, 
         ImgReg1IN_376, ImgReg1IN_375, ImgReg1IN_374, ImgReg1IN_373, 
         ImgReg1IN_372, ImgReg1IN_371, ImgReg1IN_370, ImgReg1IN_369, 
         ImgReg1IN_368, ImgReg1IN_367, ImgReg1IN_366, ImgReg1IN_365, 
         ImgReg1IN_364, ImgReg1IN_363, ImgReg1IN_362, ImgReg1IN_361, 
         ImgReg1IN_360, ImgReg1IN_359, ImgReg1IN_358, ImgReg1IN_357, 
         ImgReg1IN_356, ImgReg1IN_355, ImgReg1IN_354, ImgReg1IN_353, 
         ImgReg1IN_352, ImgReg1IN_351, ImgReg1IN_350, ImgReg1IN_349, 
         ImgReg1IN_348, ImgReg1IN_347, ImgReg1IN_346, ImgReg1IN_345, 
         ImgReg1IN_344, ImgReg1IN_343, ImgReg1IN_342, ImgReg1IN_341, 
         ImgReg1IN_340, ImgReg1IN_339, ImgReg1IN_338, ImgReg1IN_337, 
         ImgReg1IN_336, ImgReg1IN_335, ImgReg1IN_334, ImgReg1IN_333, 
         ImgReg1IN_332, ImgReg1IN_331, ImgReg1IN_330, ImgReg1IN_329, 
         ImgReg1IN_328, ImgReg1IN_327, ImgReg1IN_326, ImgReg1IN_325, 
         ImgReg1IN_324, ImgReg1IN_323, ImgReg1IN_322, ImgReg1IN_321, 
         ImgReg1IN_320, ImgReg1IN_319, ImgReg1IN_318, ImgReg1IN_317, 
         ImgReg1IN_316, ImgReg1IN_315, ImgReg1IN_314, ImgReg1IN_313, 
         ImgReg1IN_312, ImgReg1IN_311, ImgReg1IN_310, ImgReg1IN_309, 
         ImgReg1IN_308, ImgReg1IN_307, ImgReg1IN_306, ImgReg1IN_305, 
         ImgReg1IN_304, ImgReg1IN_303, ImgReg1IN_302, ImgReg1IN_301, 
         ImgReg1IN_300, ImgReg1IN_299, ImgReg1IN_298, ImgReg1IN_297, 
         ImgReg1IN_296, ImgReg1IN_295, ImgReg1IN_294, ImgReg1IN_293, 
         ImgReg1IN_292, ImgReg1IN_291, ImgReg1IN_290, ImgReg1IN_289, 
         ImgReg1IN_288, ImgReg1IN_287, ImgReg1IN_286, ImgReg1IN_285, 
         ImgReg1IN_284, ImgReg1IN_283, ImgReg1IN_282, ImgReg1IN_281, 
         ImgReg1IN_280, ImgReg1IN_279, ImgReg1IN_278, ImgReg1IN_277, 
         ImgReg1IN_276, ImgReg1IN_275, ImgReg1IN_274, ImgReg1IN_273, 
         ImgReg1IN_272, ImgReg1IN_271, ImgReg1IN_270, ImgReg1IN_269, 
         ImgReg1IN_268, ImgReg1IN_267, ImgReg1IN_266, ImgReg1IN_265, 
         ImgReg1IN_264, ImgReg1IN_263, ImgReg1IN_262, ImgReg1IN_261, 
         ImgReg1IN_260, ImgReg1IN_259, ImgReg1IN_258, ImgReg1IN_257, 
         ImgReg1IN_256, ImgReg1IN_255, ImgReg1IN_254, ImgReg1IN_253, 
         ImgReg1IN_252, ImgReg1IN_251, ImgReg1IN_250, ImgReg1IN_249, 
         ImgReg1IN_248, ImgReg1IN_247, ImgReg1IN_246, ImgReg1IN_245, 
         ImgReg1IN_244, ImgReg1IN_243, ImgReg1IN_242, ImgReg1IN_241, 
         ImgReg1IN_240, ImgReg1IN_239, ImgReg1IN_238, ImgReg1IN_237, 
         ImgReg1IN_236, ImgReg1IN_235, ImgReg1IN_234, ImgReg1IN_233, 
         ImgReg1IN_232, ImgReg1IN_231, ImgReg1IN_230, ImgReg1IN_229, 
         ImgReg1IN_228, ImgReg1IN_227, ImgReg1IN_226, ImgReg1IN_225, 
         ImgReg1IN_224, ImgReg1IN_223, ImgReg1IN_222, ImgReg1IN_221, 
         ImgReg1IN_220, ImgReg1IN_219, ImgReg1IN_218, ImgReg1IN_217, 
         ImgReg1IN_216, ImgReg1IN_215, ImgReg1IN_214, ImgReg1IN_213, 
         ImgReg1IN_212, ImgReg1IN_211, ImgReg1IN_210, ImgReg1IN_209, 
         ImgReg1IN_208, ImgReg1IN_207, ImgReg1IN_206, ImgReg1IN_205, 
         ImgReg1IN_204, ImgReg1IN_203, ImgReg1IN_202, ImgReg1IN_201, 
         ImgReg1IN_200, ImgReg1IN_199, ImgReg1IN_198, ImgReg1IN_197, 
         ImgReg1IN_196, ImgReg1IN_195, ImgReg1IN_194, ImgReg1IN_193, 
         ImgReg1IN_192, ImgReg1IN_191, ImgReg1IN_190, ImgReg1IN_189, 
         ImgReg1IN_188, ImgReg1IN_187, ImgReg1IN_186, ImgReg1IN_185, 
         ImgReg1IN_184, ImgReg1IN_183, ImgReg1IN_182, ImgReg1IN_181, 
         ImgReg1IN_180, ImgReg1IN_179, ImgReg1IN_178, ImgReg1IN_177, 
         ImgReg1IN_176, ImgReg1IN_175, ImgReg1IN_174, ImgReg1IN_173, 
         ImgReg1IN_172, ImgReg1IN_171, ImgReg1IN_170, ImgReg1IN_169, 
         ImgReg1IN_168, ImgReg1IN_167, ImgReg1IN_166, ImgReg1IN_165, 
         ImgReg1IN_164, ImgReg1IN_163, ImgReg1IN_162, ImgReg1IN_161, 
         ImgReg1IN_160, ImgReg1IN_159, ImgReg1IN_158, ImgReg1IN_157, 
         ImgReg1IN_156, ImgReg1IN_155, ImgReg1IN_154, ImgReg1IN_153, 
         ImgReg1IN_152, ImgReg1IN_151, ImgReg1IN_150, ImgReg1IN_149, 
         ImgReg1IN_148, ImgReg1IN_147, ImgReg1IN_146, ImgReg1IN_145, 
         ImgReg1IN_144, ImgReg1IN_143, ImgReg1IN_142, ImgReg1IN_141, 
         ImgReg1IN_140, ImgReg1IN_139, ImgReg1IN_138, ImgReg1IN_137, 
         ImgReg1IN_136, ImgReg1IN_135, ImgReg1IN_134, ImgReg1IN_133, 
         ImgReg1IN_132, ImgReg1IN_131, ImgReg1IN_130, ImgReg1IN_129, 
         ImgReg1IN_128, ImgReg1IN_127, ImgReg1IN_126, ImgReg1IN_125, 
         ImgReg1IN_124, ImgReg1IN_123, ImgReg1IN_122, ImgReg1IN_121, 
         ImgReg1IN_120, ImgReg1IN_119, ImgReg1IN_118, ImgReg1IN_117, 
         ImgReg1IN_116, ImgReg1IN_115, ImgReg1IN_114, ImgReg1IN_113, 
         ImgReg1IN_112, ImgReg1IN_111, ImgReg1IN_110, ImgReg1IN_109, 
         ImgReg1IN_108, ImgReg1IN_107, ImgReg1IN_106, ImgReg1IN_105, 
         ImgReg1IN_104, ImgReg1IN_103, ImgReg1IN_102, ImgReg1IN_101, 
         ImgReg1IN_100, ImgReg1IN_99, ImgReg1IN_98, ImgReg1IN_97, ImgReg1IN_96, 
         ImgReg1IN_95, ImgReg1IN_94, ImgReg1IN_93, ImgReg1IN_92, ImgReg1IN_91, 
         ImgReg1IN_90, ImgReg1IN_89, ImgReg1IN_88, ImgReg1IN_87, ImgReg1IN_86, 
         ImgReg1IN_85, ImgReg1IN_84, ImgReg1IN_83, ImgReg1IN_82, ImgReg1IN_81, 
         ImgReg1IN_80, ImgReg1IN_79, ImgReg1IN_78, ImgReg1IN_77, ImgReg1IN_76, 
         ImgReg1IN_75, ImgReg1IN_74, ImgReg1IN_73, ImgReg1IN_72, ImgReg1IN_71, 
         ImgReg1IN_70, ImgReg1IN_69, ImgReg1IN_68, ImgReg1IN_67, ImgReg1IN_66, 
         ImgReg1IN_65, ImgReg1IN_64, ImgReg1IN_63, ImgReg1IN_62, ImgReg1IN_61, 
         ImgReg1IN_60, ImgReg1IN_59, ImgReg1IN_58, ImgReg1IN_57, ImgReg1IN_56, 
         ImgReg1IN_55, ImgReg1IN_54, ImgReg1IN_53, ImgReg1IN_52, ImgReg1IN_51, 
         ImgReg1IN_50, ImgReg1IN_49, ImgReg1IN_48, ImgReg1IN_47, ImgReg1IN_46, 
         ImgReg1IN_45, ImgReg1IN_44, ImgReg1IN_43, ImgReg1IN_42, ImgReg1IN_41, 
         ImgReg1IN_40, ImgReg1IN_39, ImgReg1IN_38, ImgReg1IN_37, ImgReg1IN_36, 
         ImgReg1IN_35, ImgReg1IN_34, ImgReg1IN_33, ImgReg1IN_32, ImgReg1IN_31, 
         ImgReg1IN_30, ImgReg1IN_29, ImgReg1IN_28, ImgReg1IN_27, ImgReg1IN_26, 
         ImgReg1IN_25, ImgReg1IN_24, ImgReg1IN_23, ImgReg1IN_22, ImgReg1IN_21, 
         ImgReg1IN_20, ImgReg1IN_19, ImgReg1IN_18, ImgReg1IN_17, ImgReg1IN_16, 
         ImgReg1IN_15, ImgReg1IN_14, ImgReg1IN_13, ImgReg1IN_12, ImgReg1IN_11, 
         ImgReg1IN_10, ImgReg1IN_9, ImgReg1IN_8, ImgReg1IN_7, ImgReg1IN_6, 
         ImgReg1IN_5, ImgReg1IN_4, ImgReg1IN_3, ImgReg1IN_2, ImgReg1IN_1, 
         ImgReg1IN_0, ImgReg2IN_447, ImgReg2IN_446, ImgReg2IN_445, ImgReg2IN_444, 
         ImgReg2IN_443, ImgReg2IN_442, ImgReg2IN_441, ImgReg2IN_440, 
         ImgReg2IN_439, ImgReg2IN_438, ImgReg2IN_437, ImgReg2IN_436, 
         ImgReg2IN_435, ImgReg2IN_434, ImgReg2IN_433, ImgReg2IN_432, 
         ImgReg2IN_431, ImgReg2IN_430, ImgReg2IN_429, ImgReg2IN_428, 
         ImgReg2IN_427, ImgReg2IN_426, ImgReg2IN_425, ImgReg2IN_424, 
         ImgReg2IN_423, ImgReg2IN_422, ImgReg2IN_421, ImgReg2IN_420, 
         ImgReg2IN_419, ImgReg2IN_418, ImgReg2IN_417, ImgReg2IN_416, 
         ImgReg2IN_415, ImgReg2IN_414, ImgReg2IN_413, ImgReg2IN_412, 
         ImgReg2IN_411, ImgReg2IN_410, ImgReg2IN_409, ImgReg2IN_408, 
         ImgReg2IN_407, ImgReg2IN_406, ImgReg2IN_405, ImgReg2IN_404, 
         ImgReg2IN_403, ImgReg2IN_402, ImgReg2IN_401, ImgReg2IN_400, 
         ImgReg2IN_399, ImgReg2IN_398, ImgReg2IN_397, ImgReg2IN_396, 
         ImgReg2IN_395, ImgReg2IN_394, ImgReg2IN_393, ImgReg2IN_392, 
         ImgReg2IN_391, ImgReg2IN_390, ImgReg2IN_389, ImgReg2IN_388, 
         ImgReg2IN_387, ImgReg2IN_386, ImgReg2IN_385, ImgReg2IN_384, 
         ImgReg2IN_383, ImgReg2IN_382, ImgReg2IN_381, ImgReg2IN_380, 
         ImgReg2IN_379, ImgReg2IN_378, ImgReg2IN_377, ImgReg2IN_376, 
         ImgReg2IN_375, ImgReg2IN_374, ImgReg2IN_373, ImgReg2IN_372, 
         ImgReg2IN_371, ImgReg2IN_370, ImgReg2IN_369, ImgReg2IN_368, 
         ImgReg2IN_367, ImgReg2IN_366, ImgReg2IN_365, ImgReg2IN_364, 
         ImgReg2IN_363, ImgReg2IN_362, ImgReg2IN_361, ImgReg2IN_360, 
         ImgReg2IN_359, ImgReg2IN_358, ImgReg2IN_357, ImgReg2IN_356, 
         ImgReg2IN_355, ImgReg2IN_354, ImgReg2IN_353, ImgReg2IN_352, 
         ImgReg2IN_351, ImgReg2IN_350, ImgReg2IN_349, ImgReg2IN_348, 
         ImgReg2IN_347, ImgReg2IN_346, ImgReg2IN_345, ImgReg2IN_344, 
         ImgReg2IN_343, ImgReg2IN_342, ImgReg2IN_341, ImgReg2IN_340, 
         ImgReg2IN_339, ImgReg2IN_338, ImgReg2IN_337, ImgReg2IN_336, 
         ImgReg2IN_335, ImgReg2IN_334, ImgReg2IN_333, ImgReg2IN_332, 
         ImgReg2IN_331, ImgReg2IN_330, ImgReg2IN_329, ImgReg2IN_328, 
         ImgReg2IN_327, ImgReg2IN_326, ImgReg2IN_325, ImgReg2IN_324, 
         ImgReg2IN_323, ImgReg2IN_322, ImgReg2IN_321, ImgReg2IN_320, 
         ImgReg2IN_319, ImgReg2IN_318, ImgReg2IN_317, ImgReg2IN_316, 
         ImgReg2IN_315, ImgReg2IN_314, ImgReg2IN_313, ImgReg2IN_312, 
         ImgReg2IN_311, ImgReg2IN_310, ImgReg2IN_309, ImgReg2IN_308, 
         ImgReg2IN_307, ImgReg2IN_306, ImgReg2IN_305, ImgReg2IN_304, 
         ImgReg2IN_303, ImgReg2IN_302, ImgReg2IN_301, ImgReg2IN_300, 
         ImgReg2IN_299, ImgReg2IN_298, ImgReg2IN_297, ImgReg2IN_296, 
         ImgReg2IN_295, ImgReg2IN_294, ImgReg2IN_293, ImgReg2IN_292, 
         ImgReg2IN_291, ImgReg2IN_290, ImgReg2IN_289, ImgReg2IN_288, 
         ImgReg2IN_287, ImgReg2IN_286, ImgReg2IN_285, ImgReg2IN_284, 
         ImgReg2IN_283, ImgReg2IN_282, ImgReg2IN_281, ImgReg2IN_280, 
         ImgReg2IN_279, ImgReg2IN_278, ImgReg2IN_277, ImgReg2IN_276, 
         ImgReg2IN_275, ImgReg2IN_274, ImgReg2IN_273, ImgReg2IN_272, 
         ImgReg2IN_271, ImgReg2IN_270, ImgReg2IN_269, ImgReg2IN_268, 
         ImgReg2IN_267, ImgReg2IN_266, ImgReg2IN_265, ImgReg2IN_264, 
         ImgReg2IN_263, ImgReg2IN_262, ImgReg2IN_261, ImgReg2IN_260, 
         ImgReg2IN_259, ImgReg2IN_258, ImgReg2IN_257, ImgReg2IN_256, 
         ImgReg2IN_255, ImgReg2IN_254, ImgReg2IN_253, ImgReg2IN_252, 
         ImgReg2IN_251, ImgReg2IN_250, ImgReg2IN_249, ImgReg2IN_248, 
         ImgReg2IN_247, ImgReg2IN_246, ImgReg2IN_245, ImgReg2IN_244, 
         ImgReg2IN_243, ImgReg2IN_242, ImgReg2IN_241, ImgReg2IN_240, 
         ImgReg2IN_239, ImgReg2IN_238, ImgReg2IN_237, ImgReg2IN_236, 
         ImgReg2IN_235, ImgReg2IN_234, ImgReg2IN_233, ImgReg2IN_232, 
         ImgReg2IN_231, ImgReg2IN_230, ImgReg2IN_229, ImgReg2IN_228, 
         ImgReg2IN_227, ImgReg2IN_226, ImgReg2IN_225, ImgReg2IN_224, 
         ImgReg2IN_223, ImgReg2IN_222, ImgReg2IN_221, ImgReg2IN_220, 
         ImgReg2IN_219, ImgReg2IN_218, ImgReg2IN_217, ImgReg2IN_216, 
         ImgReg2IN_215, ImgReg2IN_214, ImgReg2IN_213, ImgReg2IN_212, 
         ImgReg2IN_211, ImgReg2IN_210, ImgReg2IN_209, ImgReg2IN_208, 
         ImgReg2IN_207, ImgReg2IN_206, ImgReg2IN_205, ImgReg2IN_204, 
         ImgReg2IN_203, ImgReg2IN_202, ImgReg2IN_201, ImgReg2IN_200, 
         ImgReg2IN_199, ImgReg2IN_198, ImgReg2IN_197, ImgReg2IN_196, 
         ImgReg2IN_195, ImgReg2IN_194, ImgReg2IN_193, ImgReg2IN_192, 
         ImgReg2IN_191, ImgReg2IN_190, ImgReg2IN_189, ImgReg2IN_188, 
         ImgReg2IN_187, ImgReg2IN_186, ImgReg2IN_185, ImgReg2IN_184, 
         ImgReg2IN_183, ImgReg2IN_182, ImgReg2IN_181, ImgReg2IN_180, 
         ImgReg2IN_179, ImgReg2IN_178, ImgReg2IN_177, ImgReg2IN_176, 
         ImgReg2IN_175, ImgReg2IN_174, ImgReg2IN_173, ImgReg2IN_172, 
         ImgReg2IN_171, ImgReg2IN_170, ImgReg2IN_169, ImgReg2IN_168, 
         ImgReg2IN_167, ImgReg2IN_166, ImgReg2IN_165, ImgReg2IN_164, 
         ImgReg2IN_163, ImgReg2IN_162, ImgReg2IN_161, ImgReg2IN_160, 
         ImgReg2IN_159, ImgReg2IN_158, ImgReg2IN_157, ImgReg2IN_156, 
         ImgReg2IN_155, ImgReg2IN_154, ImgReg2IN_153, ImgReg2IN_152, 
         ImgReg2IN_151, ImgReg2IN_150, ImgReg2IN_149, ImgReg2IN_148, 
         ImgReg2IN_147, ImgReg2IN_146, ImgReg2IN_145, ImgReg2IN_144, 
         ImgReg2IN_143, ImgReg2IN_142, ImgReg2IN_141, ImgReg2IN_140, 
         ImgReg2IN_139, ImgReg2IN_138, ImgReg2IN_137, ImgReg2IN_136, 
         ImgReg2IN_135, ImgReg2IN_134, ImgReg2IN_133, ImgReg2IN_132, 
         ImgReg2IN_131, ImgReg2IN_130, ImgReg2IN_129, ImgReg2IN_128, 
         ImgReg2IN_127, ImgReg2IN_126, ImgReg2IN_125, ImgReg2IN_124, 
         ImgReg2IN_123, ImgReg2IN_122, ImgReg2IN_121, ImgReg2IN_120, 
         ImgReg2IN_119, ImgReg2IN_118, ImgReg2IN_117, ImgReg2IN_116, 
         ImgReg2IN_115, ImgReg2IN_114, ImgReg2IN_113, ImgReg2IN_112, 
         ImgReg2IN_111, ImgReg2IN_110, ImgReg2IN_109, ImgReg2IN_108, 
         ImgReg2IN_107, ImgReg2IN_106, ImgReg2IN_105, ImgReg2IN_104, 
         ImgReg2IN_103, ImgReg2IN_102, ImgReg2IN_101, ImgReg2IN_100, 
         ImgReg2IN_99, ImgReg2IN_98, ImgReg2IN_97, ImgReg2IN_96, ImgReg2IN_95, 
         ImgReg2IN_94, ImgReg2IN_93, ImgReg2IN_92, ImgReg2IN_91, ImgReg2IN_90, 
         ImgReg2IN_89, ImgReg2IN_88, ImgReg2IN_87, ImgReg2IN_86, ImgReg2IN_85, 
         ImgReg2IN_84, ImgReg2IN_83, ImgReg2IN_82, ImgReg2IN_81, ImgReg2IN_80, 
         ImgReg2IN_79, ImgReg2IN_78, ImgReg2IN_77, ImgReg2IN_76, ImgReg2IN_75, 
         ImgReg2IN_74, ImgReg2IN_73, ImgReg2IN_72, ImgReg2IN_71, ImgReg2IN_70, 
         ImgReg2IN_69, ImgReg2IN_68, ImgReg2IN_67, ImgReg2IN_66, ImgReg2IN_65, 
         ImgReg2IN_64, ImgReg2IN_63, ImgReg2IN_62, ImgReg2IN_61, ImgReg2IN_60, 
         ImgReg2IN_59, ImgReg2IN_58, ImgReg2IN_57, ImgReg2IN_56, ImgReg2IN_55, 
         ImgReg2IN_54, ImgReg2IN_53, ImgReg2IN_52, ImgReg2IN_51, ImgReg2IN_50, 
         ImgReg2IN_49, ImgReg2IN_48, ImgReg2IN_47, ImgReg2IN_46, ImgReg2IN_45, 
         ImgReg2IN_44, ImgReg2IN_43, ImgReg2IN_42, ImgReg2IN_41, ImgReg2IN_40, 
         ImgReg2IN_39, ImgReg2IN_38, ImgReg2IN_37, ImgReg2IN_36, ImgReg2IN_35, 
         ImgReg2IN_34, ImgReg2IN_33, ImgReg2IN_32, ImgReg2IN_31, ImgReg2IN_30, 
         ImgReg2IN_29, ImgReg2IN_28, ImgReg2IN_27, ImgReg2IN_26, ImgReg2IN_25, 
         ImgReg2IN_24, ImgReg2IN_23, ImgReg2IN_22, ImgReg2IN_21, ImgReg2IN_20, 
         ImgReg2IN_19, ImgReg2IN_18, ImgReg2IN_17, ImgReg2IN_16, ImgReg2IN_15, 
         ImgReg2IN_14, ImgReg2IN_13, ImgReg2IN_12, ImgReg2IN_11, ImgReg2IN_10, 
         ImgReg2IN_9, ImgReg2IN_8, ImgReg2IN_7, ImgReg2IN_6, ImgReg2IN_5, 
         ImgReg2IN_4, ImgReg2IN_3, ImgReg2IN_2, ImgReg2IN_1, ImgReg2IN_0, 
         ImgReg3IN_447, ImgReg3IN_446, ImgReg3IN_445, ImgReg3IN_444, 
         ImgReg3IN_443, ImgReg3IN_442, ImgReg3IN_441, ImgReg3IN_440, 
         ImgReg3IN_439, ImgReg3IN_438, ImgReg3IN_437, ImgReg3IN_436, 
         ImgReg3IN_435, ImgReg3IN_434, ImgReg3IN_433, ImgReg3IN_432, 
         ImgReg3IN_431, ImgReg3IN_430, ImgReg3IN_429, ImgReg3IN_428, 
         ImgReg3IN_427, ImgReg3IN_426, ImgReg3IN_425, ImgReg3IN_424, 
         ImgReg3IN_423, ImgReg3IN_422, ImgReg3IN_421, ImgReg3IN_420, 
         ImgReg3IN_419, ImgReg3IN_418, ImgReg3IN_417, ImgReg3IN_416, 
         ImgReg3IN_415, ImgReg3IN_414, ImgReg3IN_413, ImgReg3IN_412, 
         ImgReg3IN_411, ImgReg3IN_410, ImgReg3IN_409, ImgReg3IN_408, 
         ImgReg3IN_407, ImgReg3IN_406, ImgReg3IN_405, ImgReg3IN_404, 
         ImgReg3IN_403, ImgReg3IN_402, ImgReg3IN_401, ImgReg3IN_400, 
         ImgReg3IN_399, ImgReg3IN_398, ImgReg3IN_397, ImgReg3IN_396, 
         ImgReg3IN_395, ImgReg3IN_394, ImgReg3IN_393, ImgReg3IN_392, 
         ImgReg3IN_391, ImgReg3IN_390, ImgReg3IN_389, ImgReg3IN_388, 
         ImgReg3IN_387, ImgReg3IN_386, ImgReg3IN_385, ImgReg3IN_384, 
         ImgReg3IN_383, ImgReg3IN_382, ImgReg3IN_381, ImgReg3IN_380, 
         ImgReg3IN_379, ImgReg3IN_378, ImgReg3IN_377, ImgReg3IN_376, 
         ImgReg3IN_375, ImgReg3IN_374, ImgReg3IN_373, ImgReg3IN_372, 
         ImgReg3IN_371, ImgReg3IN_370, ImgReg3IN_369, ImgReg3IN_368, 
         ImgReg3IN_367, ImgReg3IN_366, ImgReg3IN_365, ImgReg3IN_364, 
         ImgReg3IN_363, ImgReg3IN_362, ImgReg3IN_361, ImgReg3IN_360, 
         ImgReg3IN_359, ImgReg3IN_358, ImgReg3IN_357, ImgReg3IN_356, 
         ImgReg3IN_355, ImgReg3IN_354, ImgReg3IN_353, ImgReg3IN_352, 
         ImgReg3IN_351, ImgReg3IN_350, ImgReg3IN_349, ImgReg3IN_348, 
         ImgReg3IN_347, ImgReg3IN_346, ImgReg3IN_345, ImgReg3IN_344, 
         ImgReg3IN_343, ImgReg3IN_342, ImgReg3IN_341, ImgReg3IN_340, 
         ImgReg3IN_339, ImgReg3IN_338, ImgReg3IN_337, ImgReg3IN_336, 
         ImgReg3IN_335, ImgReg3IN_334, ImgReg3IN_333, ImgReg3IN_332, 
         ImgReg3IN_331, ImgReg3IN_330, ImgReg3IN_329, ImgReg3IN_328, 
         ImgReg3IN_327, ImgReg3IN_326, ImgReg3IN_325, ImgReg3IN_324, 
         ImgReg3IN_323, ImgReg3IN_322, ImgReg3IN_321, ImgReg3IN_320, 
         ImgReg3IN_319, ImgReg3IN_318, ImgReg3IN_317, ImgReg3IN_316, 
         ImgReg3IN_315, ImgReg3IN_314, ImgReg3IN_313, ImgReg3IN_312, 
         ImgReg3IN_311, ImgReg3IN_310, ImgReg3IN_309, ImgReg3IN_308, 
         ImgReg3IN_307, ImgReg3IN_306, ImgReg3IN_305, ImgReg3IN_304, 
         ImgReg3IN_303, ImgReg3IN_302, ImgReg3IN_301, ImgReg3IN_300, 
         ImgReg3IN_299, ImgReg3IN_298, ImgReg3IN_297, ImgReg3IN_296, 
         ImgReg3IN_295, ImgReg3IN_294, ImgReg3IN_293, ImgReg3IN_292, 
         ImgReg3IN_291, ImgReg3IN_290, ImgReg3IN_289, ImgReg3IN_288, 
         ImgReg3IN_287, ImgReg3IN_286, ImgReg3IN_285, ImgReg3IN_284, 
         ImgReg3IN_283, ImgReg3IN_282, ImgReg3IN_281, ImgReg3IN_280, 
         ImgReg3IN_279, ImgReg3IN_278, ImgReg3IN_277, ImgReg3IN_276, 
         ImgReg3IN_275, ImgReg3IN_274, ImgReg3IN_273, ImgReg3IN_272, 
         ImgReg3IN_271, ImgReg3IN_270, ImgReg3IN_269, ImgReg3IN_268, 
         ImgReg3IN_267, ImgReg3IN_266, ImgReg3IN_265, ImgReg3IN_264, 
         ImgReg3IN_263, ImgReg3IN_262, ImgReg3IN_261, ImgReg3IN_260, 
         ImgReg3IN_259, ImgReg3IN_258, ImgReg3IN_257, ImgReg3IN_256, 
         ImgReg3IN_255, ImgReg3IN_254, ImgReg3IN_253, ImgReg3IN_252, 
         ImgReg3IN_251, ImgReg3IN_250, ImgReg3IN_249, ImgReg3IN_248, 
         ImgReg3IN_247, ImgReg3IN_246, ImgReg3IN_245, ImgReg3IN_244, 
         ImgReg3IN_243, ImgReg3IN_242, ImgReg3IN_241, ImgReg3IN_240, 
         ImgReg3IN_239, ImgReg3IN_238, ImgReg3IN_237, ImgReg3IN_236, 
         ImgReg3IN_235, ImgReg3IN_234, ImgReg3IN_233, ImgReg3IN_232, 
         ImgReg3IN_231, ImgReg3IN_230, ImgReg3IN_229, ImgReg3IN_228, 
         ImgReg3IN_227, ImgReg3IN_226, ImgReg3IN_225, ImgReg3IN_224, 
         ImgReg3IN_223, ImgReg3IN_222, ImgReg3IN_221, ImgReg3IN_220, 
         ImgReg3IN_219, ImgReg3IN_218, ImgReg3IN_217, ImgReg3IN_216, 
         ImgReg3IN_215, ImgReg3IN_214, ImgReg3IN_213, ImgReg3IN_212, 
         ImgReg3IN_211, ImgReg3IN_210, ImgReg3IN_209, ImgReg3IN_208, 
         ImgReg3IN_207, ImgReg3IN_206, ImgReg3IN_205, ImgReg3IN_204, 
         ImgReg3IN_203, ImgReg3IN_202, ImgReg3IN_201, ImgReg3IN_200, 
         ImgReg3IN_199, ImgReg3IN_198, ImgReg3IN_197, ImgReg3IN_196, 
         ImgReg3IN_195, ImgReg3IN_194, ImgReg3IN_193, ImgReg3IN_192, 
         ImgReg3IN_191, ImgReg3IN_190, ImgReg3IN_189, ImgReg3IN_188, 
         ImgReg3IN_187, ImgReg3IN_186, ImgReg3IN_185, ImgReg3IN_184, 
         ImgReg3IN_183, ImgReg3IN_182, ImgReg3IN_181, ImgReg3IN_180, 
         ImgReg3IN_179, ImgReg3IN_178, ImgReg3IN_177, ImgReg3IN_176, 
         ImgReg3IN_175, ImgReg3IN_174, ImgReg3IN_173, ImgReg3IN_172, 
         ImgReg3IN_171, ImgReg3IN_170, ImgReg3IN_169, ImgReg3IN_168, 
         ImgReg3IN_167, ImgReg3IN_166, ImgReg3IN_165, ImgReg3IN_164, 
         ImgReg3IN_163, ImgReg3IN_162, ImgReg3IN_161, ImgReg3IN_160, 
         ImgReg3IN_159, ImgReg3IN_158, ImgReg3IN_157, ImgReg3IN_156, 
         ImgReg3IN_155, ImgReg3IN_154, ImgReg3IN_153, ImgReg3IN_152, 
         ImgReg3IN_151, ImgReg3IN_150, ImgReg3IN_149, ImgReg3IN_148, 
         ImgReg3IN_147, ImgReg3IN_146, ImgReg3IN_145, ImgReg3IN_144, 
         ImgReg3IN_143, ImgReg3IN_142, ImgReg3IN_141, ImgReg3IN_140, 
         ImgReg3IN_139, ImgReg3IN_138, ImgReg3IN_137, ImgReg3IN_136, 
         ImgReg3IN_135, ImgReg3IN_134, ImgReg3IN_133, ImgReg3IN_132, 
         ImgReg3IN_131, ImgReg3IN_130, ImgReg3IN_129, ImgReg3IN_128, 
         ImgReg3IN_127, ImgReg3IN_126, ImgReg3IN_125, ImgReg3IN_124, 
         ImgReg3IN_123, ImgReg3IN_122, ImgReg3IN_121, ImgReg3IN_120, 
         ImgReg3IN_119, ImgReg3IN_118, ImgReg3IN_117, ImgReg3IN_116, 
         ImgReg3IN_115, ImgReg3IN_114, ImgReg3IN_113, ImgReg3IN_112, 
         ImgReg3IN_111, ImgReg3IN_110, ImgReg3IN_109, ImgReg3IN_108, 
         ImgReg3IN_107, ImgReg3IN_106, ImgReg3IN_105, ImgReg3IN_104, 
         ImgReg3IN_103, ImgReg3IN_102, ImgReg3IN_101, ImgReg3IN_100, 
         ImgReg3IN_99, ImgReg3IN_98, ImgReg3IN_97, ImgReg3IN_96, ImgReg3IN_95, 
         ImgReg3IN_94, ImgReg3IN_93, ImgReg3IN_92, ImgReg3IN_91, ImgReg3IN_90, 
         ImgReg3IN_89, ImgReg3IN_88, ImgReg3IN_87, ImgReg3IN_86, ImgReg3IN_85, 
         ImgReg3IN_84, ImgReg3IN_83, ImgReg3IN_82, ImgReg3IN_81, ImgReg3IN_80, 
         ImgReg3IN_79, ImgReg3IN_78, ImgReg3IN_77, ImgReg3IN_76, ImgReg3IN_75, 
         ImgReg3IN_74, ImgReg3IN_73, ImgReg3IN_72, ImgReg3IN_71, ImgReg3IN_70, 
         ImgReg3IN_69, ImgReg3IN_68, ImgReg3IN_67, ImgReg3IN_66, ImgReg3IN_65, 
         ImgReg3IN_64, ImgReg3IN_63, ImgReg3IN_62, ImgReg3IN_61, ImgReg3IN_60, 
         ImgReg3IN_59, ImgReg3IN_58, ImgReg3IN_57, ImgReg3IN_56, ImgReg3IN_55, 
         ImgReg3IN_54, ImgReg3IN_53, ImgReg3IN_52, ImgReg3IN_51, ImgReg3IN_50, 
         ImgReg3IN_49, ImgReg3IN_48, ImgReg3IN_47, ImgReg3IN_46, ImgReg3IN_45, 
         ImgReg3IN_44, ImgReg3IN_43, ImgReg3IN_42, ImgReg3IN_41, ImgReg3IN_40, 
         ImgReg3IN_39, ImgReg3IN_38, ImgReg3IN_37, ImgReg3IN_36, ImgReg3IN_35, 
         ImgReg3IN_34, ImgReg3IN_33, ImgReg3IN_32, ImgReg3IN_31, ImgReg3IN_30, 
         ImgReg3IN_29, ImgReg3IN_28, ImgReg3IN_27, ImgReg3IN_26, ImgReg3IN_25, 
         ImgReg3IN_24, ImgReg3IN_23, ImgReg3IN_22, ImgReg3IN_21, ImgReg3IN_20, 
         ImgReg3IN_19, ImgReg3IN_18, ImgReg3IN_17, ImgReg3IN_16, ImgReg3IN_15, 
         ImgReg3IN_14, ImgReg3IN_13, ImgReg3IN_12, ImgReg3IN_11, ImgReg3IN_10, 
         ImgReg3IN_9, ImgReg3IN_8, ImgReg3IN_7, ImgReg3IN_6, ImgReg3IN_5, 
         ImgReg3IN_4, ImgReg3IN_3, ImgReg3IN_2, ImgReg3IN_1, ImgReg3IN_0, 
         ImgReg4IN_447, ImgReg4IN_446, ImgReg4IN_445, ImgReg4IN_444, 
         ImgReg4IN_443, ImgReg4IN_442, ImgReg4IN_441, ImgReg4IN_440, 
         ImgReg4IN_439, ImgReg4IN_438, ImgReg4IN_437, ImgReg4IN_436, 
         ImgReg4IN_435, ImgReg4IN_434, ImgReg4IN_433, ImgReg4IN_432, 
         ImgReg4IN_431, ImgReg4IN_430, ImgReg4IN_429, ImgReg4IN_428, 
         ImgReg4IN_427, ImgReg4IN_426, ImgReg4IN_425, ImgReg4IN_424, 
         ImgReg4IN_423, ImgReg4IN_422, ImgReg4IN_421, ImgReg4IN_420, 
         ImgReg4IN_419, ImgReg4IN_418, ImgReg4IN_417, ImgReg4IN_416, 
         ImgReg4IN_415, ImgReg4IN_414, ImgReg4IN_413, ImgReg4IN_412, 
         ImgReg4IN_411, ImgReg4IN_410, ImgReg4IN_409, ImgReg4IN_408, 
         ImgReg4IN_407, ImgReg4IN_406, ImgReg4IN_405, ImgReg4IN_404, 
         ImgReg4IN_403, ImgReg4IN_402, ImgReg4IN_401, ImgReg4IN_400, 
         ImgReg4IN_399, ImgReg4IN_398, ImgReg4IN_397, ImgReg4IN_396, 
         ImgReg4IN_395, ImgReg4IN_394, ImgReg4IN_393, ImgReg4IN_392, 
         ImgReg4IN_391, ImgReg4IN_390, ImgReg4IN_389, ImgReg4IN_388, 
         ImgReg4IN_387, ImgReg4IN_386, ImgReg4IN_385, ImgReg4IN_384, 
         ImgReg4IN_383, ImgReg4IN_382, ImgReg4IN_381, ImgReg4IN_380, 
         ImgReg4IN_379, ImgReg4IN_378, ImgReg4IN_377, ImgReg4IN_376, 
         ImgReg4IN_375, ImgReg4IN_374, ImgReg4IN_373, ImgReg4IN_372, 
         ImgReg4IN_371, ImgReg4IN_370, ImgReg4IN_369, ImgReg4IN_368, 
         ImgReg4IN_367, ImgReg4IN_366, ImgReg4IN_365, ImgReg4IN_364, 
         ImgReg4IN_363, ImgReg4IN_362, ImgReg4IN_361, ImgReg4IN_360, 
         ImgReg4IN_359, ImgReg4IN_358, ImgReg4IN_357, ImgReg4IN_356, 
         ImgReg4IN_355, ImgReg4IN_354, ImgReg4IN_353, ImgReg4IN_352, 
         ImgReg4IN_351, ImgReg4IN_350, ImgReg4IN_349, ImgReg4IN_348, 
         ImgReg4IN_347, ImgReg4IN_346, ImgReg4IN_345, ImgReg4IN_344, 
         ImgReg4IN_343, ImgReg4IN_342, ImgReg4IN_341, ImgReg4IN_340, 
         ImgReg4IN_339, ImgReg4IN_338, ImgReg4IN_337, ImgReg4IN_336, 
         ImgReg4IN_335, ImgReg4IN_334, ImgReg4IN_333, ImgReg4IN_332, 
         ImgReg4IN_331, ImgReg4IN_330, ImgReg4IN_329, ImgReg4IN_328, 
         ImgReg4IN_327, ImgReg4IN_326, ImgReg4IN_325, ImgReg4IN_324, 
         ImgReg4IN_323, ImgReg4IN_322, ImgReg4IN_321, ImgReg4IN_320, 
         ImgReg4IN_319, ImgReg4IN_318, ImgReg4IN_317, ImgReg4IN_316, 
         ImgReg4IN_315, ImgReg4IN_314, ImgReg4IN_313, ImgReg4IN_312, 
         ImgReg4IN_311, ImgReg4IN_310, ImgReg4IN_309, ImgReg4IN_308, 
         ImgReg4IN_307, ImgReg4IN_306, ImgReg4IN_305, ImgReg4IN_304, 
         ImgReg4IN_303, ImgReg4IN_302, ImgReg4IN_301, ImgReg4IN_300, 
         ImgReg4IN_299, ImgReg4IN_298, ImgReg4IN_297, ImgReg4IN_296, 
         ImgReg4IN_295, ImgReg4IN_294, ImgReg4IN_293, ImgReg4IN_292, 
         ImgReg4IN_291, ImgReg4IN_290, ImgReg4IN_289, ImgReg4IN_288, 
         ImgReg4IN_287, ImgReg4IN_286, ImgReg4IN_285, ImgReg4IN_284, 
         ImgReg4IN_283, ImgReg4IN_282, ImgReg4IN_281, ImgReg4IN_280, 
         ImgReg4IN_279, ImgReg4IN_278, ImgReg4IN_277, ImgReg4IN_276, 
         ImgReg4IN_275, ImgReg4IN_274, ImgReg4IN_273, ImgReg4IN_272, 
         ImgReg4IN_271, ImgReg4IN_270, ImgReg4IN_269, ImgReg4IN_268, 
         ImgReg4IN_267, ImgReg4IN_266, ImgReg4IN_265, ImgReg4IN_264, 
         ImgReg4IN_263, ImgReg4IN_262, ImgReg4IN_261, ImgReg4IN_260, 
         ImgReg4IN_259, ImgReg4IN_258, ImgReg4IN_257, ImgReg4IN_256, 
         ImgReg4IN_255, ImgReg4IN_254, ImgReg4IN_253, ImgReg4IN_252, 
         ImgReg4IN_251, ImgReg4IN_250, ImgReg4IN_249, ImgReg4IN_248, 
         ImgReg4IN_247, ImgReg4IN_246, ImgReg4IN_245, ImgReg4IN_244, 
         ImgReg4IN_243, ImgReg4IN_242, ImgReg4IN_241, ImgReg4IN_240, 
         ImgReg4IN_239, ImgReg4IN_238, ImgReg4IN_237, ImgReg4IN_236, 
         ImgReg4IN_235, ImgReg4IN_234, ImgReg4IN_233, ImgReg4IN_232, 
         ImgReg4IN_231, ImgReg4IN_230, ImgReg4IN_229, ImgReg4IN_228, 
         ImgReg4IN_227, ImgReg4IN_226, ImgReg4IN_225, ImgReg4IN_224, 
         ImgReg4IN_223, ImgReg4IN_222, ImgReg4IN_221, ImgReg4IN_220, 
         ImgReg4IN_219, ImgReg4IN_218, ImgReg4IN_217, ImgReg4IN_216, 
         ImgReg4IN_215, ImgReg4IN_214, ImgReg4IN_213, ImgReg4IN_212, 
         ImgReg4IN_211, ImgReg4IN_210, ImgReg4IN_209, ImgReg4IN_208, 
         ImgReg4IN_207, ImgReg4IN_206, ImgReg4IN_205, ImgReg4IN_204, 
         ImgReg4IN_203, ImgReg4IN_202, ImgReg4IN_201, ImgReg4IN_200, 
         ImgReg4IN_199, ImgReg4IN_198, ImgReg4IN_197, ImgReg4IN_196, 
         ImgReg4IN_195, ImgReg4IN_194, ImgReg4IN_193, ImgReg4IN_192, 
         ImgReg4IN_191, ImgReg4IN_190, ImgReg4IN_189, ImgReg4IN_188, 
         ImgReg4IN_187, ImgReg4IN_186, ImgReg4IN_185, ImgReg4IN_184, 
         ImgReg4IN_183, ImgReg4IN_182, ImgReg4IN_181, ImgReg4IN_180, 
         ImgReg4IN_179, ImgReg4IN_178, ImgReg4IN_177, ImgReg4IN_176, 
         ImgReg4IN_175, ImgReg4IN_174, ImgReg4IN_173, ImgReg4IN_172, 
         ImgReg4IN_171, ImgReg4IN_170, ImgReg4IN_169, ImgReg4IN_168, 
         ImgReg4IN_167, ImgReg4IN_166, ImgReg4IN_165, ImgReg4IN_164, 
         ImgReg4IN_163, ImgReg4IN_162, ImgReg4IN_161, ImgReg4IN_160, 
         ImgReg4IN_159, ImgReg4IN_158, ImgReg4IN_157, ImgReg4IN_156, 
         ImgReg4IN_155, ImgReg4IN_154, ImgReg4IN_153, ImgReg4IN_152, 
         ImgReg4IN_151, ImgReg4IN_150, ImgReg4IN_149, ImgReg4IN_148, 
         ImgReg4IN_147, ImgReg4IN_146, ImgReg4IN_145, ImgReg4IN_144, 
         ImgReg4IN_143, ImgReg4IN_142, ImgReg4IN_141, ImgReg4IN_140, 
         ImgReg4IN_139, ImgReg4IN_138, ImgReg4IN_137, ImgReg4IN_136, 
         ImgReg4IN_135, ImgReg4IN_134, ImgReg4IN_133, ImgReg4IN_132, 
         ImgReg4IN_131, ImgReg4IN_130, ImgReg4IN_129, ImgReg4IN_128, 
         ImgReg4IN_127, ImgReg4IN_126, ImgReg4IN_125, ImgReg4IN_124, 
         ImgReg4IN_123, ImgReg4IN_122, ImgReg4IN_121, ImgReg4IN_120, 
         ImgReg4IN_119, ImgReg4IN_118, ImgReg4IN_117, ImgReg4IN_116, 
         ImgReg4IN_115, ImgReg4IN_114, ImgReg4IN_113, ImgReg4IN_112, 
         ImgReg4IN_111, ImgReg4IN_110, ImgReg4IN_109, ImgReg4IN_108, 
         ImgReg4IN_107, ImgReg4IN_106, ImgReg4IN_105, ImgReg4IN_104, 
         ImgReg4IN_103, ImgReg4IN_102, ImgReg4IN_101, ImgReg4IN_100, 
         ImgReg4IN_99, ImgReg4IN_98, ImgReg4IN_97, ImgReg4IN_96, ImgReg4IN_95, 
         ImgReg4IN_94, ImgReg4IN_93, ImgReg4IN_92, ImgReg4IN_91, ImgReg4IN_90, 
         ImgReg4IN_89, ImgReg4IN_88, ImgReg4IN_87, ImgReg4IN_86, ImgReg4IN_85, 
         ImgReg4IN_84, ImgReg4IN_83, ImgReg4IN_82, ImgReg4IN_81, ImgReg4IN_80, 
         ImgReg4IN_79, ImgReg4IN_78, ImgReg4IN_77, ImgReg4IN_76, ImgReg4IN_75, 
         ImgReg4IN_74, ImgReg4IN_73, ImgReg4IN_72, ImgReg4IN_71, ImgReg4IN_70, 
         ImgReg4IN_69, ImgReg4IN_68, ImgReg4IN_67, ImgReg4IN_66, ImgReg4IN_65, 
         ImgReg4IN_64, ImgReg4IN_63, ImgReg4IN_62, ImgReg4IN_61, ImgReg4IN_60, 
         ImgReg4IN_59, ImgReg4IN_58, ImgReg4IN_57, ImgReg4IN_56, ImgReg4IN_55, 
         ImgReg4IN_54, ImgReg4IN_53, ImgReg4IN_52, ImgReg4IN_51, ImgReg4IN_50, 
         ImgReg4IN_49, ImgReg4IN_48, ImgReg4IN_47, ImgReg4IN_46, ImgReg4IN_45, 
         ImgReg4IN_44, ImgReg4IN_43, ImgReg4IN_42, ImgReg4IN_41, ImgReg4IN_40, 
         ImgReg4IN_39, ImgReg4IN_38, ImgReg4IN_37, ImgReg4IN_36, ImgReg4IN_35, 
         ImgReg4IN_34, ImgReg4IN_33, ImgReg4IN_32, ImgReg4IN_31, ImgReg4IN_30, 
         ImgReg4IN_29, ImgReg4IN_28, ImgReg4IN_27, ImgReg4IN_26, ImgReg4IN_25, 
         ImgReg4IN_24, ImgReg4IN_23, ImgReg4IN_22, ImgReg4IN_21, ImgReg4IN_20, 
         ImgReg4IN_19, ImgReg4IN_18, ImgReg4IN_17, ImgReg4IN_16, ImgReg4IN_15, 
         ImgReg4IN_14, ImgReg4IN_13, ImgReg4IN_12, ImgReg4IN_11, ImgReg4IN_10, 
         ImgReg4IN_9, ImgReg4IN_8, ImgReg4IN_7, ImgReg4IN_6, ImgReg4IN_5, 
         ImgReg4IN_4, ImgReg4IN_3, ImgReg4IN_2, ImgReg4IN_1, ImgReg4IN_0, 
         ImgReg5IN_447, ImgReg5IN_446, ImgReg5IN_445, ImgReg5IN_444, 
         ImgReg5IN_443, ImgReg5IN_442, ImgReg5IN_441, ImgReg5IN_440, 
         ImgReg5IN_439, ImgReg5IN_438, ImgReg5IN_437, ImgReg5IN_436, 
         ImgReg5IN_435, ImgReg5IN_434, ImgReg5IN_433, ImgReg5IN_432, 
         ImgReg5IN_431, ImgReg5IN_430, ImgReg5IN_429, ImgReg5IN_428, 
         ImgReg5IN_427, ImgReg5IN_426, ImgReg5IN_425, ImgReg5IN_424, 
         ImgReg5IN_423, ImgReg5IN_422, ImgReg5IN_421, ImgReg5IN_420, 
         ImgReg5IN_419, ImgReg5IN_418, ImgReg5IN_417, ImgReg5IN_416, 
         ImgReg5IN_415, ImgReg5IN_414, ImgReg5IN_413, ImgReg5IN_412, 
         ImgReg5IN_411, ImgReg5IN_410, ImgReg5IN_409, ImgReg5IN_408, 
         ImgReg5IN_407, ImgReg5IN_406, ImgReg5IN_405, ImgReg5IN_404, 
         ImgReg5IN_403, ImgReg5IN_402, ImgReg5IN_401, ImgReg5IN_400, 
         ImgReg5IN_399, ImgReg5IN_398, ImgReg5IN_397, ImgReg5IN_396, 
         ImgReg5IN_395, ImgReg5IN_394, ImgReg5IN_393, ImgReg5IN_392, 
         ImgReg5IN_391, ImgReg5IN_390, ImgReg5IN_389, ImgReg5IN_388, 
         ImgReg5IN_387, ImgReg5IN_386, ImgReg5IN_385, ImgReg5IN_384, 
         ImgReg5IN_383, ImgReg5IN_382, ImgReg5IN_381, ImgReg5IN_380, 
         ImgReg5IN_379, ImgReg5IN_378, ImgReg5IN_377, ImgReg5IN_376, 
         ImgReg5IN_375, ImgReg5IN_374, ImgReg5IN_373, ImgReg5IN_372, 
         ImgReg5IN_371, ImgReg5IN_370, ImgReg5IN_369, ImgReg5IN_368, 
         ImgReg5IN_367, ImgReg5IN_366, ImgReg5IN_365, ImgReg5IN_364, 
         ImgReg5IN_363, ImgReg5IN_362, ImgReg5IN_361, ImgReg5IN_360, 
         ImgReg5IN_359, ImgReg5IN_358, ImgReg5IN_357, ImgReg5IN_356, 
         ImgReg5IN_355, ImgReg5IN_354, ImgReg5IN_353, ImgReg5IN_352, 
         ImgReg5IN_351, ImgReg5IN_350, ImgReg5IN_349, ImgReg5IN_348, 
         ImgReg5IN_347, ImgReg5IN_346, ImgReg5IN_345, ImgReg5IN_344, 
         ImgReg5IN_343, ImgReg5IN_342, ImgReg5IN_341, ImgReg5IN_340, 
         ImgReg5IN_339, ImgReg5IN_338, ImgReg5IN_337, ImgReg5IN_336, 
         ImgReg5IN_335, ImgReg5IN_334, ImgReg5IN_333, ImgReg5IN_332, 
         ImgReg5IN_331, ImgReg5IN_330, ImgReg5IN_329, ImgReg5IN_328, 
         ImgReg5IN_327, ImgReg5IN_326, ImgReg5IN_325, ImgReg5IN_324, 
         ImgReg5IN_323, ImgReg5IN_322, ImgReg5IN_321, ImgReg5IN_320, 
         ImgReg5IN_319, ImgReg5IN_318, ImgReg5IN_317, ImgReg5IN_316, 
         ImgReg5IN_315, ImgReg5IN_314, ImgReg5IN_313, ImgReg5IN_312, 
         ImgReg5IN_311, ImgReg5IN_310, ImgReg5IN_309, ImgReg5IN_308, 
         ImgReg5IN_307, ImgReg5IN_306, ImgReg5IN_305, ImgReg5IN_304, 
         ImgReg5IN_303, ImgReg5IN_302, ImgReg5IN_301, ImgReg5IN_300, 
         ImgReg5IN_299, ImgReg5IN_298, ImgReg5IN_297, ImgReg5IN_296, 
         ImgReg5IN_295, ImgReg5IN_294, ImgReg5IN_293, ImgReg5IN_292, 
         ImgReg5IN_291, ImgReg5IN_290, ImgReg5IN_289, ImgReg5IN_288, 
         ImgReg5IN_287, ImgReg5IN_286, ImgReg5IN_285, ImgReg5IN_284, 
         ImgReg5IN_283, ImgReg5IN_282, ImgReg5IN_281, ImgReg5IN_280, 
         ImgReg5IN_279, ImgReg5IN_278, ImgReg5IN_277, ImgReg5IN_276, 
         ImgReg5IN_275, ImgReg5IN_274, ImgReg5IN_273, ImgReg5IN_272, 
         ImgReg5IN_271, ImgReg5IN_270, ImgReg5IN_269, ImgReg5IN_268, 
         ImgReg5IN_267, ImgReg5IN_266, ImgReg5IN_265, ImgReg5IN_264, 
         ImgReg5IN_263, ImgReg5IN_262, ImgReg5IN_261, ImgReg5IN_260, 
         ImgReg5IN_259, ImgReg5IN_258, ImgReg5IN_257, ImgReg5IN_256, 
         ImgReg5IN_255, ImgReg5IN_254, ImgReg5IN_253, ImgReg5IN_252, 
         ImgReg5IN_251, ImgReg5IN_250, ImgReg5IN_249, ImgReg5IN_248, 
         ImgReg5IN_247, ImgReg5IN_246, ImgReg5IN_245, ImgReg5IN_244, 
         ImgReg5IN_243, ImgReg5IN_242, ImgReg5IN_241, ImgReg5IN_240, 
         ImgReg5IN_239, ImgReg5IN_238, ImgReg5IN_237, ImgReg5IN_236, 
         ImgReg5IN_235, ImgReg5IN_234, ImgReg5IN_233, ImgReg5IN_232, 
         ImgReg5IN_231, ImgReg5IN_230, ImgReg5IN_229, ImgReg5IN_228, 
         ImgReg5IN_227, ImgReg5IN_226, ImgReg5IN_225, ImgReg5IN_224, 
         ImgReg5IN_223, ImgReg5IN_222, ImgReg5IN_221, ImgReg5IN_220, 
         ImgReg5IN_219, ImgReg5IN_218, ImgReg5IN_217, ImgReg5IN_216, 
         ImgReg5IN_215, ImgReg5IN_214, ImgReg5IN_213, ImgReg5IN_212, 
         ImgReg5IN_211, ImgReg5IN_210, ImgReg5IN_209, ImgReg5IN_208, 
         ImgReg5IN_207, ImgReg5IN_206, ImgReg5IN_205, ImgReg5IN_204, 
         ImgReg5IN_203, ImgReg5IN_202, ImgReg5IN_201, ImgReg5IN_200, 
         ImgReg5IN_199, ImgReg5IN_198, ImgReg5IN_197, ImgReg5IN_196, 
         ImgReg5IN_195, ImgReg5IN_194, ImgReg5IN_193, ImgReg5IN_192, 
         ImgReg5IN_191, ImgReg5IN_190, ImgReg5IN_189, ImgReg5IN_188, 
         ImgReg5IN_187, ImgReg5IN_186, ImgReg5IN_185, ImgReg5IN_184, 
         ImgReg5IN_183, ImgReg5IN_182, ImgReg5IN_181, ImgReg5IN_180, 
         ImgReg5IN_179, ImgReg5IN_178, ImgReg5IN_177, ImgReg5IN_176, 
         ImgReg5IN_175, ImgReg5IN_174, ImgReg5IN_173, ImgReg5IN_172, 
         ImgReg5IN_171, ImgReg5IN_170, ImgReg5IN_169, ImgReg5IN_168, 
         ImgReg5IN_167, ImgReg5IN_166, ImgReg5IN_165, ImgReg5IN_164, 
         ImgReg5IN_163, ImgReg5IN_162, ImgReg5IN_161, ImgReg5IN_160, 
         ImgReg5IN_159, ImgReg5IN_158, ImgReg5IN_157, ImgReg5IN_156, 
         ImgReg5IN_155, ImgReg5IN_154, ImgReg5IN_153, ImgReg5IN_152, 
         ImgReg5IN_151, ImgReg5IN_150, ImgReg5IN_149, ImgReg5IN_148, 
         ImgReg5IN_147, ImgReg5IN_146, ImgReg5IN_145, ImgReg5IN_144, 
         ImgReg5IN_143, ImgReg5IN_142, ImgReg5IN_141, ImgReg5IN_140, 
         ImgReg5IN_139, ImgReg5IN_138, ImgReg5IN_137, ImgReg5IN_136, 
         ImgReg5IN_135, ImgReg5IN_134, ImgReg5IN_133, ImgReg5IN_132, 
         ImgReg5IN_131, ImgReg5IN_130, ImgReg5IN_129, ImgReg5IN_128, 
         ImgReg5IN_127, ImgReg5IN_126, ImgReg5IN_125, ImgReg5IN_124, 
         ImgReg5IN_123, ImgReg5IN_122, ImgReg5IN_121, ImgReg5IN_120, 
         ImgReg5IN_119, ImgReg5IN_118, ImgReg5IN_117, ImgReg5IN_116, 
         ImgReg5IN_115, ImgReg5IN_114, ImgReg5IN_113, ImgReg5IN_112, 
         ImgReg5IN_111, ImgReg5IN_110, ImgReg5IN_109, ImgReg5IN_108, 
         ImgReg5IN_107, ImgReg5IN_106, ImgReg5IN_105, ImgReg5IN_104, 
         ImgReg5IN_103, ImgReg5IN_102, ImgReg5IN_101, ImgReg5IN_100, 
         ImgReg5IN_99, ImgReg5IN_98, ImgReg5IN_97, ImgReg5IN_96, ImgReg5IN_95, 
         ImgReg5IN_94, ImgReg5IN_93, ImgReg5IN_92, ImgReg5IN_91, ImgReg5IN_90, 
         ImgReg5IN_89, ImgReg5IN_88, ImgReg5IN_87, ImgReg5IN_86, ImgReg5IN_85, 
         ImgReg5IN_84, ImgReg5IN_83, ImgReg5IN_82, ImgReg5IN_81, ImgReg5IN_80, 
         ImgReg5IN_79, ImgReg5IN_78, ImgReg5IN_77, ImgReg5IN_76, ImgReg5IN_75, 
         ImgReg5IN_74, ImgReg5IN_73, ImgReg5IN_72, ImgReg5IN_71, ImgReg5IN_70, 
         ImgReg5IN_69, ImgReg5IN_68, ImgReg5IN_67, ImgReg5IN_66, ImgReg5IN_65, 
         ImgReg5IN_64, ImgReg5IN_63, ImgReg5IN_62, ImgReg5IN_61, ImgReg5IN_60, 
         ImgReg5IN_59, ImgReg5IN_58, ImgReg5IN_57, ImgReg5IN_56, ImgReg5IN_55, 
         ImgReg5IN_54, ImgReg5IN_53, ImgReg5IN_52, ImgReg5IN_51, ImgReg5IN_50, 
         ImgReg5IN_49, ImgReg5IN_48, ImgReg5IN_47, ImgReg5IN_46, ImgReg5IN_45, 
         ImgReg5IN_44, ImgReg5IN_43, ImgReg5IN_42, ImgReg5IN_41, ImgReg5IN_40, 
         ImgReg5IN_39, ImgReg5IN_38, ImgReg5IN_37, ImgReg5IN_36, ImgReg5IN_35, 
         ImgReg5IN_34, ImgReg5IN_33, ImgReg5IN_32, ImgReg5IN_31, ImgReg5IN_30, 
         ImgReg5IN_29, ImgReg5IN_28, ImgReg5IN_27, ImgReg5IN_26, ImgReg5IN_25, 
         ImgReg5IN_24, ImgReg5IN_23, ImgReg5IN_22, ImgReg5IN_21, ImgReg5IN_20, 
         ImgReg5IN_19, ImgReg5IN_18, ImgReg5IN_17, ImgReg5IN_16, ImgReg5IN_15, 
         ImgReg5IN_14, ImgReg5IN_13, ImgReg5IN_12, ImgReg5IN_11, ImgReg5IN_10, 
         ImgReg5IN_9, ImgReg5IN_8, ImgReg5IN_7, ImgReg5IN_6, ImgReg5IN_5, 
         ImgReg5IN_4, ImgReg5IN_3, ImgReg5IN_2, ImgReg5IN_1, ImgReg5IN_0, 
         TriAddEn, IndRst, cReset, cEnable, TriImgRegEn, TriImgLeftEn, PWR, 
         firstOperand_15, nx2, nx20, nx34, NOT_ImgIndic_0, nx23568, nx23573, 
         nx23580, nx23583, nx23592, nx23594, nx23596, nx23598, nx23600, nx23604, 
         nx23606, nx23608, nx23610, nx23612, nx23616, nx23618, nx23620, nx23622, 
         nx23624, nx23628, nx23630, nx23632, nx23634, nx23636, nx23640, nx23642, 
         nx23644, nx23646, nx23648, nx23652, nx23654, nx23656, nx23658, nx23660, 
         nx23664, nx23666, nx23668, nx23670, nx23672, nx23674, nx23676, nx23678, 
         nx23680, nx23682, nx23684, nx23686, nx23688, nx23690, nx23692, nx23694, 
         nx23696, nx23698, nx23700, nx23702, nx23704, nx23706, nx23708, nx23710, 
         nx23712, nx23716, nx23718, nx23720, nx23722, nx23724, nx23726, nx23728, 
         nx23730, nx23732, nx23734, nx23736, nx23738, nx23740, nx23742, nx23744, 
         nx23746, nx23748, nx23750, nx23752, nx23754, nx23756, nx23758, nx23760, 
         nx23762, nx23764, nx23766, nx23768, nx23770, nx23772, nx23774, nx23776, 
         nx23778, nx23780, nx23786, nx23788, nx23790, nx23792, nx23794, nx23796, 
         nx23798, nx23800, nx23802, nx23804, nx23806, nx23808, nx23810, nx23812, 
         nx23814, nx23816, nx23818, nx23820, nx23822, nx23824, nx23828, nx23830, 
         nx23832, nx23834, nx23836, nx23838, nx23840, nx23842, nx23844, nx23846, 
         nx23848, nx23850, nx23852, nx23854, nx23856, nx23858, nx23860, nx23862, 
         nx23864, nx23866, nx23868, nx23870, nx23872, nx23874, nx23876, nx23878, 
         nx23880, nx23882, nx23884, nx23886, nx23888, nx23890, nx23892, nx23894, 
         nx23896, nx23898, nx23900, nx23902, nx23904, nx23906, nx23908, nx23910, 
         nx23912, nx23914, nx23916, nx23918, nx23920, nx23922, nx23924, nx23926, 
         nx23928, nx23930, nx23932, nx23934, nx23936, nx23938, nx23940, nx23942, 
         nx23944, nx23946, nx23948, nx23950, nx23952, nx23954, nx23956, nx23958, 
         nx23960, nx23962, nx23964, nx23966, nx23968, nx23970, nx23972, nx23974, 
         nx23976, nx23978, nx23980, nx23982, nx23984, nx23986, nx23988, nx23990, 
         nx23992, nx23994, nx23996, nx23998, nx24000, nx24002, nx24004, nx24006, 
         nx24008, nx24010, nx24012, nx24014, nx24016, nx24018, nx24020, nx24022, 
         nx24024, nx24026, nx24028, nx24030, nx24032, nx24038, nx24040;
    wire [4:0] \$dummy ;




    my_nadder_16 adder0 (.a ({firstOperand_15,firstOperand_15,firstOperand_15,
                 ImgAddress[12],ImgAddress[11],ImgAddress[10],ImgAddress[9],
                 ImgAddress[8],ImgAddress[7],ImgAddress[6],ImgAddress[5],
                 ImgAddress[4],ImgAddress[3],ImgAddress[2],ImgAddress[1],
                 ImgAddress[0]}), .b ({ImgWidth[15],ImgWidth[14],ImgWidth[13],
                 ImgWidth[12],ImgWidth[11],ImgWidth[10],ImgWidth[9],ImgWidth[8],
                 ImgWidth[7],ImgWidth[6],ImgWidth[5],ImgWidth[4],ImgWidth[3],
                 ImgWidth[2],ImgWidth[1],ImgWidth[0]}), .cin (firstOperand_15), 
                 .s ({\$dummy [0],\$dummy [1],\$dummy [2],newAdd16_12,
                 newAdd16_11,newAdd16_10,newAdd16_9,newAdd16_8,newAdd16_7,
                 newAdd16_6,newAdd16_5,newAdd16_4,newAdd16_3,newAdd16_2,
                 newAdd16_1,newAdd16_0}), .cout (\$dummy [3])) ;
    triStateBuffer_13 triStateAdd (.D ({newAdd16_12,newAdd16_11,newAdd16_10,
                      newAdd16_9,newAdd16_8,newAdd16_7,newAdd16_6,newAdd16_5,
                      newAdd16_4,newAdd16_3,newAdd16_2,newAdd16_1,newAdd16_0}), 
                      .EN (TriAddEn), .F ({UpdatedAddress[12],UpdatedAddress[11]
                      ,UpdatedAddress[10],UpdatedAddress[9],UpdatedAddress[8],
                      UpdatedAddress[7],UpdatedAddress[6],UpdatedAddress[5],
                      UpdatedAddress[4],UpdatedAddress[3],UpdatedAddress[2],
                      UpdatedAddress[1],UpdatedAddress[0]})) ;
    triStateBuffer_13 TriStateAddToDma (.D ({ImgAddress[12],ImgAddress[11],
                      ImgAddress[10],ImgAddress[9],ImgAddress[8],ImgAddress[7],
                      ImgAddress[6],ImgAddress[5],ImgAddress[4],ImgAddress[3],
                      ImgAddress[2],ImgAddress[1],ImgAddress[0]}), .EN (TriAddEn
                      ), .F ({ImgAddToDma[12],ImgAddToDma[11],ImgAddToDma[10],
                      ImgAddToDma[9],ImgAddToDma[8],ImgAddToDma[7],
                      ImgAddToDma[6],ImgAddToDma[5],ImgAddToDma[4],
                      ImgAddToDma[3],ImgAddToDma[2],ImgAddToDma[1],
                      ImgAddToDma[0]})) ;
    nBitRegister_1 DDF0 (.D ({NOT_ImgIndic_0}), .CLK (DFFCLK), .RST (IndRst), .EN (
                   PWR), .Q ({ImgIndic[0]})) ;
    Counter_3 RegCounter0 (.enable (cEnable), .reset (cReset), .clk (nx23828), .load (
              firstOperand_15), .\output  ({ImgCounterOuput[2],
              ImgCounterOuput[1],ImgCounterOuput[0]}), .\input  ({
              firstOperand_15,firstOperand_15,PWR})) ;
    Decoder dec (.\input  ({ImgCounterOuput[2],ImgCounterOuput[1],
            ImgCounterOuput[0]}), .\output  ({DecOutput_5,DecOutput_4,
            DecOutput_3,DecOutput_2,DecOutput_1,DecOutput_0})) ;
    triStateBuffer_6 TriImgReg (.D ({DecOutput_5,DecOutput_4,DecOutput_3,
                     DecOutput_2,DecOutput_1,DecOutput_0}), .EN (TriImgRegEn), .F (
                     {ImgEn[5],ImgEn[4],ImgEn[3],ImgEn[2],ImgEn[1],ImgEn[0]})) ;
    triStateBuffer_16 loop3_0_TriState0L (.D ({OutputImg0[31],OutputImg0[30],
                      OutputImg0[29],OutputImg0[28],OutputImg0[27],
                      OutputImg0[26],OutputImg0[25],OutputImg0[24],
                      OutputImg0[23],OutputImg0[22],OutputImg0[21],
                      OutputImg0[20],OutputImg0[19],OutputImg0[18],
                      OutputImg0[17],OutputImg0[16]}), .EN (nx23666), .F ({
                      ImgReg0IN_15,ImgReg0IN_14,ImgReg0IN_13,ImgReg0IN_12,
                      ImgReg0IN_11,ImgReg0IN_10,ImgReg0IN_9,ImgReg0IN_8,
                      ImgReg0IN_7,ImgReg0IN_6,ImgReg0IN_5,ImgReg0IN_4,
                      ImgReg0IN_3,ImgReg0IN_2,ImgReg0IN_1,ImgReg0IN_0})) ;
    triStateBuffer_16 loop3_0_TriState1L (.D ({OutputImg1[31],OutputImg1[30],
                      OutputImg1[29],OutputImg1[28],OutputImg1[27],
                      OutputImg1[26],OutputImg1[25],OutputImg1[24],
                      OutputImg1[23],OutputImg1[22],OutputImg1[21],
                      OutputImg1[20],OutputImg1[19],OutputImg1[18],
                      OutputImg1[17],OutputImg1[16]}), .EN (nx23666), .F ({
                      ImgReg1IN_15,ImgReg1IN_14,ImgReg1IN_13,ImgReg1IN_12,
                      ImgReg1IN_11,ImgReg1IN_10,ImgReg1IN_9,ImgReg1IN_8,
                      ImgReg1IN_7,ImgReg1IN_6,ImgReg1IN_5,ImgReg1IN_4,
                      ImgReg1IN_3,ImgReg1IN_2,ImgReg1IN_1,ImgReg1IN_0})) ;
    triStateBuffer_16 loop3_0_TriState2L (.D ({OutputImg2[31],OutputImg2[30],
                      OutputImg2[29],OutputImg2[28],OutputImg2[27],
                      OutputImg2[26],OutputImg2[25],OutputImg2[24],
                      OutputImg2[23],OutputImg2[22],OutputImg2[21],
                      OutputImg2[20],OutputImg2[19],OutputImg2[18],
                      OutputImg2[17],OutputImg2[16]}), .EN (nx23666), .F ({
                      ImgReg2IN_15,ImgReg2IN_14,ImgReg2IN_13,ImgReg2IN_12,
                      ImgReg2IN_11,ImgReg2IN_10,ImgReg2IN_9,ImgReg2IN_8,
                      ImgReg2IN_7,ImgReg2IN_6,ImgReg2IN_5,ImgReg2IN_4,
                      ImgReg2IN_3,ImgReg2IN_2,ImgReg2IN_1,ImgReg2IN_0})) ;
    triStateBuffer_16 loop3_0_TriState3L (.D ({OutputImg3[31],OutputImg3[30],
                      OutputImg3[29],OutputImg3[28],OutputImg3[27],
                      OutputImg3[26],OutputImg3[25],OutputImg3[24],
                      OutputImg3[23],OutputImg3[22],OutputImg3[21],
                      OutputImg3[20],OutputImg3[19],OutputImg3[18],
                      OutputImg3[17],OutputImg3[16]}), .EN (nx23666), .F ({
                      ImgReg3IN_15,ImgReg3IN_14,ImgReg3IN_13,ImgReg3IN_12,
                      ImgReg3IN_11,ImgReg3IN_10,ImgReg3IN_9,ImgReg3IN_8,
                      ImgReg3IN_7,ImgReg3IN_6,ImgReg3IN_5,ImgReg3IN_4,
                      ImgReg3IN_3,ImgReg3IN_2,ImgReg3IN_1,ImgReg3IN_0})) ;
    triStateBuffer_16 loop3_0_TriState4L (.D ({OutputImg4[31],OutputImg4[30],
                      OutputImg4[29],OutputImg4[28],OutputImg4[27],
                      OutputImg4[26],OutputImg4[25],OutputImg4[24],
                      OutputImg4[23],OutputImg4[22],OutputImg4[21],
                      OutputImg4[20],OutputImg4[19],OutputImg4[18],
                      OutputImg4[17],OutputImg4[16]}), .EN (nx23666), .F ({
                      ImgReg4IN_15,ImgReg4IN_14,ImgReg4IN_13,ImgReg4IN_12,
                      ImgReg4IN_11,ImgReg4IN_10,ImgReg4IN_9,ImgReg4IN_8,
                      ImgReg4IN_7,ImgReg4IN_6,ImgReg4IN_5,ImgReg4IN_4,
                      ImgReg4IN_3,ImgReg4IN_2,ImgReg4IN_1,ImgReg4IN_0})) ;
    triStateBuffer_16 loop3_0_TriState5L (.D ({OutputImg5[31],OutputImg5[30],
                      OutputImg5[29],OutputImg5[28],OutputImg5[27],
                      OutputImg5[26],OutputImg5[25],OutputImg5[24],
                      OutputImg5[23],OutputImg5[22],OutputImg5[21],
                      OutputImg5[20],OutputImg5[19],OutputImg5[18],
                      OutputImg5[17],OutputImg5[16]}), .EN (nx23666), .F ({
                      ImgReg5IN_15,ImgReg5IN_14,ImgReg5IN_13,ImgReg5IN_12,
                      ImgReg5IN_11,ImgReg5IN_10,ImgReg5IN_9,ImgReg5IN_8,
                      ImgReg5IN_7,ImgReg5IN_6,ImgReg5IN_5,ImgReg5IN_4,
                      ImgReg5IN_3,ImgReg5IN_2,ImgReg5IN_1,ImgReg5IN_0})) ;
    triStateBuffer_16 loop3_0_TriState0N (.D ({DATA[15],DATA[14],DATA[13],
                      DATA[12],DATA[11],DATA[10],DATA[9],DATA[8],DATA[7],DATA[6]
                      ,DATA[5],DATA[4],DATA[3],DATA[2],DATA[1],DATA[0]}), .EN (
                      nx23654), .F ({ImgReg0IN_15,ImgReg0IN_14,ImgReg0IN_13,
                      ImgReg0IN_12,ImgReg0IN_11,ImgReg0IN_10,ImgReg0IN_9,
                      ImgReg0IN_8,ImgReg0IN_7,ImgReg0IN_6,ImgReg0IN_5,
                      ImgReg0IN_4,ImgReg0IN_3,ImgReg0IN_2,ImgReg0IN_1,
                      ImgReg0IN_0})) ;
    triStateBuffer_16 loop3_0_TriState1N (.D ({DATA[15],DATA[14],DATA[13],
                      DATA[12],DATA[11],DATA[10],DATA[9],DATA[8],DATA[7],DATA[6]
                      ,DATA[5],DATA[4],DATA[3],DATA[2],DATA[1],DATA[0]}), .EN (
                      nx23642), .F ({ImgReg1IN_15,ImgReg1IN_14,ImgReg1IN_13,
                      ImgReg1IN_12,ImgReg1IN_11,ImgReg1IN_10,ImgReg1IN_9,
                      ImgReg1IN_8,ImgReg1IN_7,ImgReg1IN_6,ImgReg1IN_5,
                      ImgReg1IN_4,ImgReg1IN_3,ImgReg1IN_2,ImgReg1IN_1,
                      ImgReg1IN_0})) ;
    triStateBuffer_16 loop3_0_TriState2N (.D ({DATA[15],DATA[14],DATA[13],
                      DATA[12],DATA[11],DATA[10],DATA[9],DATA[8],DATA[7],DATA[6]
                      ,DATA[5],DATA[4],DATA[3],DATA[2],DATA[1],DATA[0]}), .EN (
                      nx23630), .F ({ImgReg2IN_15,ImgReg2IN_14,ImgReg2IN_13,
                      ImgReg2IN_12,ImgReg2IN_11,ImgReg2IN_10,ImgReg2IN_9,
                      ImgReg2IN_8,ImgReg2IN_7,ImgReg2IN_6,ImgReg2IN_5,
                      ImgReg2IN_4,ImgReg2IN_3,ImgReg2IN_2,ImgReg2IN_1,
                      ImgReg2IN_0})) ;
    triStateBuffer_16 loop3_0_TriState3N (.D ({DATA[15],DATA[14],DATA[13],
                      DATA[12],DATA[11],DATA[10],DATA[9],DATA[8],DATA[7],DATA[6]
                      ,DATA[5],DATA[4],DATA[3],DATA[2],DATA[1],DATA[0]}), .EN (
                      nx23618), .F ({ImgReg3IN_15,ImgReg3IN_14,ImgReg3IN_13,
                      ImgReg3IN_12,ImgReg3IN_11,ImgReg3IN_10,ImgReg3IN_9,
                      ImgReg3IN_8,ImgReg3IN_7,ImgReg3IN_6,ImgReg3IN_5,
                      ImgReg3IN_4,ImgReg3IN_3,ImgReg3IN_2,ImgReg3IN_1,
                      ImgReg3IN_0})) ;
    triStateBuffer_16 loop3_0_TriState4N (.D ({DATA[15],DATA[14],DATA[13],
                      DATA[12],DATA[11],DATA[10],DATA[9],DATA[8],DATA[7],DATA[6]
                      ,DATA[5],DATA[4],DATA[3],DATA[2],DATA[1],DATA[0]}), .EN (
                      nx23606), .F ({ImgReg4IN_15,ImgReg4IN_14,ImgReg4IN_13,
                      ImgReg4IN_12,ImgReg4IN_11,ImgReg4IN_10,ImgReg4IN_9,
                      ImgReg4IN_8,ImgReg4IN_7,ImgReg4IN_6,ImgReg4IN_5,
                      ImgReg4IN_4,ImgReg4IN_3,ImgReg4IN_2,ImgReg4IN_1,
                      ImgReg4IN_0})) ;
    triStateBuffer_16 loop3_0_TriState5N (.D ({DATA[15],DATA[14],DATA[13],
                      DATA[12],DATA[11],DATA[10],DATA[9],DATA[8],DATA[7],DATA[6]
                      ,DATA[5],DATA[4],DATA[3],DATA[2],DATA[1],DATA[0]}), .EN (
                      nx23594), .F ({ImgReg5IN_15,ImgReg5IN_14,ImgReg5IN_13,
                      ImgReg5IN_12,ImgReg5IN_11,ImgReg5IN_10,ImgReg5IN_9,
                      ImgReg5IN_8,ImgReg5IN_7,ImgReg5IN_6,ImgReg5IN_5,
                      ImgReg5IN_4,ImgReg5IN_3,ImgReg5IN_2,ImgReg5IN_1,
                      ImgReg5IN_0})) ;
    triStateBuffer_16 loop3_0_TriState0U (.D ({OutputImg1[15],OutputImg1[14],
                      OutputImg1[13],OutputImg1[12],OutputImg1[11],
                      OutputImg1[10],OutputImg1[9],OutputImg1[8],OutputImg1[7],
                      OutputImg1[6],OutputImg1[5],OutputImg1[4],OutputImg1[3],
                      OutputImg1[2],OutputImg1[1],OutputImg1[0]}), .EN (nx23786)
                      , .F ({ImgReg0IN_15,ImgReg0IN_14,ImgReg0IN_13,ImgReg0IN_12
                      ,ImgReg0IN_11,ImgReg0IN_10,ImgReg0IN_9,ImgReg0IN_8,
                      ImgReg0IN_7,ImgReg0IN_6,ImgReg0IN_5,ImgReg0IN_4,
                      ImgReg0IN_3,ImgReg0IN_2,ImgReg0IN_1,ImgReg0IN_0})) ;
    triStateBuffer_16 loop3_0_TriState1U (.D ({OutputImg2[15],OutputImg2[14],
                      OutputImg2[13],OutputImg2[12],OutputImg2[11],
                      OutputImg2[10],OutputImg2[9],OutputImg2[8],OutputImg2[7],
                      OutputImg2[6],OutputImg2[5],OutputImg2[4],OutputImg2[3],
                      OutputImg2[2],OutputImg2[1],OutputImg2[0]}), .EN (nx23786)
                      , .F ({ImgReg1IN_15,ImgReg1IN_14,ImgReg1IN_13,ImgReg1IN_12
                      ,ImgReg1IN_11,ImgReg1IN_10,ImgReg1IN_9,ImgReg1IN_8,
                      ImgReg1IN_7,ImgReg1IN_6,ImgReg1IN_5,ImgReg1IN_4,
                      ImgReg1IN_3,ImgReg1IN_2,ImgReg1IN_1,ImgReg1IN_0})) ;
    triStateBuffer_16 loop3_0_TriState2U (.D ({OutputImg3[15],OutputImg3[14],
                      OutputImg3[13],OutputImg3[12],OutputImg3[11],
                      OutputImg3[10],OutputImg3[9],OutputImg3[8],OutputImg3[7],
                      OutputImg3[6],OutputImg3[5],OutputImg3[4],OutputImg3[3],
                      OutputImg3[2],OutputImg3[1],OutputImg3[0]}), .EN (nx23786)
                      , .F ({ImgReg2IN_15,ImgReg2IN_14,ImgReg2IN_13,ImgReg2IN_12
                      ,ImgReg2IN_11,ImgReg2IN_10,ImgReg2IN_9,ImgReg2IN_8,
                      ImgReg2IN_7,ImgReg2IN_6,ImgReg2IN_5,ImgReg2IN_4,
                      ImgReg2IN_3,ImgReg2IN_2,ImgReg2IN_1,ImgReg2IN_0})) ;
    triStateBuffer_16 loop3_0_TriState3U (.D ({OutputImg4[15],OutputImg4[14],
                      OutputImg4[13],OutputImg4[12],OutputImg4[11],
                      OutputImg4[10],OutputImg4[9],OutputImg4[8],OutputImg4[7],
                      OutputImg4[6],OutputImg4[5],OutputImg4[4],OutputImg4[3],
                      OutputImg4[2],OutputImg4[1],OutputImg4[0]}), .EN (nx23786)
                      , .F ({ImgReg3IN_15,ImgReg3IN_14,ImgReg3IN_13,ImgReg3IN_12
                      ,ImgReg3IN_11,ImgReg3IN_10,ImgReg3IN_9,ImgReg3IN_8,
                      ImgReg3IN_7,ImgReg3IN_6,ImgReg3IN_5,ImgReg3IN_4,
                      ImgReg3IN_3,ImgReg3IN_2,ImgReg3IN_1,ImgReg3IN_0})) ;
    triStateBuffer_16 loop3_0_TriState4U (.D ({OutputImg5[15],OutputImg5[14],
                      OutputImg5[13],OutputImg5[12],OutputImg5[11],
                      OutputImg5[10],OutputImg5[9],OutputImg5[8],OutputImg5[7],
                      OutputImg5[6],OutputImg5[5],OutputImg5[4],OutputImg5[3],
                      OutputImg5[2],OutputImg5[1],OutputImg5[0]}), .EN (nx23786)
                      , .F ({ImgReg4IN_15,ImgReg4IN_14,ImgReg4IN_13,ImgReg4IN_12
                      ,ImgReg4IN_11,ImgReg4IN_10,ImgReg4IN_9,ImgReg4IN_8,
                      ImgReg4IN_7,ImgReg4IN_6,ImgReg4IN_5,ImgReg4IN_4,
                      ImgReg4IN_3,ImgReg4IN_2,ImgReg4IN_1,ImgReg4IN_0})) ;
    nBitRegister_16 loop3_0_reg1 (.D ({ImgReg0IN_15,ImgReg0IN_14,ImgReg0IN_13,
                    ImgReg0IN_12,ImgReg0IN_11,ImgReg0IN_10,ImgReg0IN_9,
                    ImgReg0IN_8,ImgReg0IN_7,ImgReg0IN_6,ImgReg0IN_5,ImgReg0IN_4,
                    ImgReg0IN_3,ImgReg0IN_2,ImgReg0IN_1,ImgReg0IN_0}), .CLK (
                    nx23828), .RST (RST), .EN (nx23718), .Q ({OutputImg0[15],
                    OutputImg0[14],OutputImg0[13],OutputImg0[12],OutputImg0[11],
                    OutputImg0[10],OutputImg0[9],OutputImg0[8],OutputImg0[7],
                    OutputImg0[6],OutputImg0[5],OutputImg0[4],OutputImg0[3],
                    OutputImg0[2],OutputImg0[1],OutputImg0[0]})) ;
    nBitRegister_16 loop3_0_reg2 (.D ({ImgReg1IN_15,ImgReg1IN_14,ImgReg1IN_13,
                    ImgReg1IN_12,ImgReg1IN_11,ImgReg1IN_10,ImgReg1IN_9,
                    ImgReg1IN_8,ImgReg1IN_7,ImgReg1IN_6,ImgReg1IN_5,ImgReg1IN_4,
                    ImgReg1IN_3,ImgReg1IN_2,ImgReg1IN_1,ImgReg1IN_0}), .CLK (
                    nx23830), .RST (RST), .EN (nx23728), .Q ({OutputImg1[15],
                    OutputImg1[14],OutputImg1[13],OutputImg1[12],OutputImg1[11],
                    OutputImg1[10],OutputImg1[9],OutputImg1[8],OutputImg1[7],
                    OutputImg1[6],OutputImg1[5],OutputImg1[4],OutputImg1[3],
                    OutputImg1[2],OutputImg1[1],OutputImg1[0]})) ;
    nBitRegister_16 loop3_0_reg3 (.D ({ImgReg2IN_15,ImgReg2IN_14,ImgReg2IN_13,
                    ImgReg2IN_12,ImgReg2IN_11,ImgReg2IN_10,ImgReg2IN_9,
                    ImgReg2IN_8,ImgReg2IN_7,ImgReg2IN_6,ImgReg2IN_5,ImgReg2IN_4,
                    ImgReg2IN_3,ImgReg2IN_2,ImgReg2IN_1,ImgReg2IN_0}), .CLK (
                    nx23830), .RST (RST), .EN (nx23738), .Q ({OutputImg2[15],
                    OutputImg2[14],OutputImg2[13],OutputImg2[12],OutputImg2[11],
                    OutputImg2[10],OutputImg2[9],OutputImg2[8],OutputImg2[7],
                    OutputImg2[6],OutputImg2[5],OutputImg2[4],OutputImg2[3],
                    OutputImg2[2],OutputImg2[1],OutputImg2[0]})) ;
    nBitRegister_16 loop3_0_reg4 (.D ({ImgReg3IN_15,ImgReg3IN_14,ImgReg3IN_13,
                    ImgReg3IN_12,ImgReg3IN_11,ImgReg3IN_10,ImgReg3IN_9,
                    ImgReg3IN_8,ImgReg3IN_7,ImgReg3IN_6,ImgReg3IN_5,ImgReg3IN_4,
                    ImgReg3IN_3,ImgReg3IN_2,ImgReg3IN_1,ImgReg3IN_0}), .CLK (
                    nx23832), .RST (RST), .EN (nx23748), .Q ({OutputImg3[15],
                    OutputImg3[14],OutputImg3[13],OutputImg3[12],OutputImg3[11],
                    OutputImg3[10],OutputImg3[9],OutputImg3[8],OutputImg3[7],
                    OutputImg3[6],OutputImg3[5],OutputImg3[4],OutputImg3[3],
                    OutputImg3[2],OutputImg3[1],OutputImg3[0]})) ;
    nBitRegister_16 loop3_0_reg5 (.D ({ImgReg4IN_15,ImgReg4IN_14,ImgReg4IN_13,
                    ImgReg4IN_12,ImgReg4IN_11,ImgReg4IN_10,ImgReg4IN_9,
                    ImgReg4IN_8,ImgReg4IN_7,ImgReg4IN_6,ImgReg4IN_5,ImgReg4IN_4,
                    ImgReg4IN_3,ImgReg4IN_2,ImgReg4IN_1,ImgReg4IN_0}), .CLK (
                    nx23832), .RST (RST), .EN (nx23758), .Q ({OutputImg4[15],
                    OutputImg4[14],OutputImg4[13],OutputImg4[12],OutputImg4[11],
                    OutputImg4[10],OutputImg4[9],OutputImg4[8],OutputImg4[7],
                    OutputImg4[6],OutputImg4[5],OutputImg4[4],OutputImg4[3],
                    OutputImg4[2],OutputImg4[1],OutputImg4[0]})) ;
    nBitRegister_16 loop3_0_reg6 (.D ({ImgReg5IN_15,ImgReg5IN_14,ImgReg5IN_13,
                    ImgReg5IN_12,ImgReg5IN_11,ImgReg5IN_10,ImgReg5IN_9,
                    ImgReg5IN_8,ImgReg5IN_7,ImgReg5IN_6,ImgReg5IN_5,ImgReg5IN_4,
                    ImgReg5IN_3,ImgReg5IN_2,ImgReg5IN_1,ImgReg5IN_0}), .CLK (
                    nx23834), .RST (RST), .EN (nx23768), .Q ({OutputImg5[15],
                    OutputImg5[14],OutputImg5[13],OutputImg5[12],OutputImg5[11],
                    OutputImg5[10],OutputImg5[9],OutputImg5[8],OutputImg5[7],
                    OutputImg5[6],OutputImg5[5],OutputImg5[4],OutputImg5[3],
                    OutputImg5[2],OutputImg5[1],OutputImg5[0]})) ;
    triStateBuffer_16 loop3_1_TriState0L (.D ({OutputImg0[47],OutputImg0[46],
                      OutputImg0[45],OutputImg0[44],OutputImg0[43],
                      OutputImg0[42],OutputImg0[41],OutputImg0[40],
                      OutputImg0[39],OutputImg0[38],OutputImg0[37],
                      OutputImg0[36],OutputImg0[35],OutputImg0[34],
                      OutputImg0[33],OutputImg0[32]}), .EN (nx23666), .F ({
                      ImgReg0IN_31,ImgReg0IN_30,ImgReg0IN_29,ImgReg0IN_28,
                      ImgReg0IN_27,ImgReg0IN_26,ImgReg0IN_25,ImgReg0IN_24,
                      ImgReg0IN_23,ImgReg0IN_22,ImgReg0IN_21,ImgReg0IN_20,
                      ImgReg0IN_19,ImgReg0IN_18,ImgReg0IN_17,ImgReg0IN_16})) ;
    triStateBuffer_16 loop3_1_TriState1L (.D ({OutputImg1[47],OutputImg1[46],
                      OutputImg1[45],OutputImg1[44],OutputImg1[43],
                      OutputImg1[42],OutputImg1[41],OutputImg1[40],
                      OutputImg1[39],OutputImg1[38],OutputImg1[37],
                      OutputImg1[36],OutputImg1[35],OutputImg1[34],
                      OutputImg1[33],OutputImg1[32]}), .EN (nx23668), .F ({
                      ImgReg1IN_31,ImgReg1IN_30,ImgReg1IN_29,ImgReg1IN_28,
                      ImgReg1IN_27,ImgReg1IN_26,ImgReg1IN_25,ImgReg1IN_24,
                      ImgReg1IN_23,ImgReg1IN_22,ImgReg1IN_21,ImgReg1IN_20,
                      ImgReg1IN_19,ImgReg1IN_18,ImgReg1IN_17,ImgReg1IN_16})) ;
    triStateBuffer_16 loop3_1_TriState2L (.D ({OutputImg2[47],OutputImg2[46],
                      OutputImg2[45],OutputImg2[44],OutputImg2[43],
                      OutputImg2[42],OutputImg2[41],OutputImg2[40],
                      OutputImg2[39],OutputImg2[38],OutputImg2[37],
                      OutputImg2[36],OutputImg2[35],OutputImg2[34],
                      OutputImg2[33],OutputImg2[32]}), .EN (nx23668), .F ({
                      ImgReg2IN_31,ImgReg2IN_30,ImgReg2IN_29,ImgReg2IN_28,
                      ImgReg2IN_27,ImgReg2IN_26,ImgReg2IN_25,ImgReg2IN_24,
                      ImgReg2IN_23,ImgReg2IN_22,ImgReg2IN_21,ImgReg2IN_20,
                      ImgReg2IN_19,ImgReg2IN_18,ImgReg2IN_17,ImgReg2IN_16})) ;
    triStateBuffer_16 loop3_1_TriState3L (.D ({OutputImg3[47],OutputImg3[46],
                      OutputImg3[45],OutputImg3[44],OutputImg3[43],
                      OutputImg3[42],OutputImg3[41],OutputImg3[40],
                      OutputImg3[39],OutputImg3[38],OutputImg3[37],
                      OutputImg3[36],OutputImg3[35],OutputImg3[34],
                      OutputImg3[33],OutputImg3[32]}), .EN (nx23668), .F ({
                      ImgReg3IN_31,ImgReg3IN_30,ImgReg3IN_29,ImgReg3IN_28,
                      ImgReg3IN_27,ImgReg3IN_26,ImgReg3IN_25,ImgReg3IN_24,
                      ImgReg3IN_23,ImgReg3IN_22,ImgReg3IN_21,ImgReg3IN_20,
                      ImgReg3IN_19,ImgReg3IN_18,ImgReg3IN_17,ImgReg3IN_16})) ;
    triStateBuffer_16 loop3_1_TriState4L (.D ({OutputImg4[47],OutputImg4[46],
                      OutputImg4[45],OutputImg4[44],OutputImg4[43],
                      OutputImg4[42],OutputImg4[41],OutputImg4[40],
                      OutputImg4[39],OutputImg4[38],OutputImg4[37],
                      OutputImg4[36],OutputImg4[35],OutputImg4[34],
                      OutputImg4[33],OutputImg4[32]}), .EN (nx23668), .F ({
                      ImgReg4IN_31,ImgReg4IN_30,ImgReg4IN_29,ImgReg4IN_28,
                      ImgReg4IN_27,ImgReg4IN_26,ImgReg4IN_25,ImgReg4IN_24,
                      ImgReg4IN_23,ImgReg4IN_22,ImgReg4IN_21,ImgReg4IN_20,
                      ImgReg4IN_19,ImgReg4IN_18,ImgReg4IN_17,ImgReg4IN_16})) ;
    triStateBuffer_16 loop3_1_TriState5L (.D ({OutputImg5[47],OutputImg5[46],
                      OutputImg5[45],OutputImg5[44],OutputImg5[43],
                      OutputImg5[42],OutputImg5[41],OutputImg5[40],
                      OutputImg5[39],OutputImg5[38],OutputImg5[37],
                      OutputImg5[36],OutputImg5[35],OutputImg5[34],
                      OutputImg5[33],OutputImg5[32]}), .EN (nx23668), .F ({
                      ImgReg5IN_31,ImgReg5IN_30,ImgReg5IN_29,ImgReg5IN_28,
                      ImgReg5IN_27,ImgReg5IN_26,ImgReg5IN_25,ImgReg5IN_24,
                      ImgReg5IN_23,ImgReg5IN_22,ImgReg5IN_21,ImgReg5IN_20,
                      ImgReg5IN_19,ImgReg5IN_18,ImgReg5IN_17,ImgReg5IN_16})) ;
    triStateBuffer_16 loop3_1_TriState0N (.D ({DATA[31],DATA[30],DATA[29],
                      DATA[28],DATA[27],DATA[26],DATA[25],DATA[24],DATA[23],
                      DATA[22],DATA[21],DATA[20],DATA[19],DATA[18],DATA[17],
                      DATA[16]}), .EN (nx23654), .F ({ImgReg0IN_31,ImgReg0IN_30,
                      ImgReg0IN_29,ImgReg0IN_28,ImgReg0IN_27,ImgReg0IN_26,
                      ImgReg0IN_25,ImgReg0IN_24,ImgReg0IN_23,ImgReg0IN_22,
                      ImgReg0IN_21,ImgReg0IN_20,ImgReg0IN_19,ImgReg0IN_18,
                      ImgReg0IN_17,ImgReg0IN_16})) ;
    triStateBuffer_16 loop3_1_TriState1N (.D ({DATA[31],DATA[30],DATA[29],
                      DATA[28],DATA[27],DATA[26],DATA[25],DATA[24],DATA[23],
                      DATA[22],DATA[21],DATA[20],DATA[19],DATA[18],DATA[17],
                      DATA[16]}), .EN (nx23642), .F ({ImgReg1IN_31,ImgReg1IN_30,
                      ImgReg1IN_29,ImgReg1IN_28,ImgReg1IN_27,ImgReg1IN_26,
                      ImgReg1IN_25,ImgReg1IN_24,ImgReg1IN_23,ImgReg1IN_22,
                      ImgReg1IN_21,ImgReg1IN_20,ImgReg1IN_19,ImgReg1IN_18,
                      ImgReg1IN_17,ImgReg1IN_16})) ;
    triStateBuffer_16 loop3_1_TriState2N (.D ({DATA[31],DATA[30],DATA[29],
                      DATA[28],DATA[27],DATA[26],DATA[25],DATA[24],DATA[23],
                      DATA[22],DATA[21],DATA[20],DATA[19],DATA[18],DATA[17],
                      DATA[16]}), .EN (nx23630), .F ({ImgReg2IN_31,ImgReg2IN_30,
                      ImgReg2IN_29,ImgReg2IN_28,ImgReg2IN_27,ImgReg2IN_26,
                      ImgReg2IN_25,ImgReg2IN_24,ImgReg2IN_23,ImgReg2IN_22,
                      ImgReg2IN_21,ImgReg2IN_20,ImgReg2IN_19,ImgReg2IN_18,
                      ImgReg2IN_17,ImgReg2IN_16})) ;
    triStateBuffer_16 loop3_1_TriState3N (.D ({DATA[31],DATA[30],DATA[29],
                      DATA[28],DATA[27],DATA[26],DATA[25],DATA[24],DATA[23],
                      DATA[22],DATA[21],DATA[20],DATA[19],DATA[18],DATA[17],
                      DATA[16]}), .EN (nx23618), .F ({ImgReg3IN_31,ImgReg3IN_30,
                      ImgReg3IN_29,ImgReg3IN_28,ImgReg3IN_27,ImgReg3IN_26,
                      ImgReg3IN_25,ImgReg3IN_24,ImgReg3IN_23,ImgReg3IN_22,
                      ImgReg3IN_21,ImgReg3IN_20,ImgReg3IN_19,ImgReg3IN_18,
                      ImgReg3IN_17,ImgReg3IN_16})) ;
    triStateBuffer_16 loop3_1_TriState4N (.D ({DATA[31],DATA[30],DATA[29],
                      DATA[28],DATA[27],DATA[26],DATA[25],DATA[24],DATA[23],
                      DATA[22],DATA[21],DATA[20],DATA[19],DATA[18],DATA[17],
                      DATA[16]}), .EN (nx23606), .F ({ImgReg4IN_31,ImgReg4IN_30,
                      ImgReg4IN_29,ImgReg4IN_28,ImgReg4IN_27,ImgReg4IN_26,
                      ImgReg4IN_25,ImgReg4IN_24,ImgReg4IN_23,ImgReg4IN_22,
                      ImgReg4IN_21,ImgReg4IN_20,ImgReg4IN_19,ImgReg4IN_18,
                      ImgReg4IN_17,ImgReg4IN_16})) ;
    triStateBuffer_16 loop3_1_TriState5N (.D ({DATA[31],DATA[30],DATA[29],
                      DATA[28],DATA[27],DATA[26],DATA[25],DATA[24],DATA[23],
                      DATA[22],DATA[21],DATA[20],DATA[19],DATA[18],DATA[17],
                      DATA[16]}), .EN (nx23594), .F ({ImgReg5IN_31,ImgReg5IN_30,
                      ImgReg5IN_29,ImgReg5IN_28,ImgReg5IN_27,ImgReg5IN_26,
                      ImgReg5IN_25,ImgReg5IN_24,ImgReg5IN_23,ImgReg5IN_22,
                      ImgReg5IN_21,ImgReg5IN_20,ImgReg5IN_19,ImgReg5IN_18,
                      ImgReg5IN_17,ImgReg5IN_16})) ;
    triStateBuffer_16 loop3_1_TriState0U (.D ({OutputImg1[31],OutputImg1[30],
                      OutputImg1[29],OutputImg1[28],OutputImg1[27],
                      OutputImg1[26],OutputImg1[25],OutputImg1[24],
                      OutputImg1[23],OutputImg1[22],OutputImg1[21],
                      OutputImg1[20],OutputImg1[19],OutputImg1[18],
                      OutputImg1[17],OutputImg1[16]}), .EN (nx23786), .F ({
                      ImgReg0IN_31,ImgReg0IN_30,ImgReg0IN_29,ImgReg0IN_28,
                      ImgReg0IN_27,ImgReg0IN_26,ImgReg0IN_25,ImgReg0IN_24,
                      ImgReg0IN_23,ImgReg0IN_22,ImgReg0IN_21,ImgReg0IN_20,
                      ImgReg0IN_19,ImgReg0IN_18,ImgReg0IN_17,ImgReg0IN_16})) ;
    triStateBuffer_16 loop3_1_TriState1U (.D ({OutputImg2[31],OutputImg2[30],
                      OutputImg2[29],OutputImg2[28],OutputImg2[27],
                      OutputImg2[26],OutputImg2[25],OutputImg2[24],
                      OutputImg2[23],OutputImg2[22],OutputImg2[21],
                      OutputImg2[20],OutputImg2[19],OutputImg2[18],
                      OutputImg2[17],OutputImg2[16]}), .EN (nx23786), .F ({
                      ImgReg1IN_31,ImgReg1IN_30,ImgReg1IN_29,ImgReg1IN_28,
                      ImgReg1IN_27,ImgReg1IN_26,ImgReg1IN_25,ImgReg1IN_24,
                      ImgReg1IN_23,ImgReg1IN_22,ImgReg1IN_21,ImgReg1IN_20,
                      ImgReg1IN_19,ImgReg1IN_18,ImgReg1IN_17,ImgReg1IN_16})) ;
    triStateBuffer_16 loop3_1_TriState2U (.D ({OutputImg3[31],OutputImg3[30],
                      OutputImg3[29],OutputImg3[28],OutputImg3[27],
                      OutputImg3[26],OutputImg3[25],OutputImg3[24],
                      OutputImg3[23],OutputImg3[22],OutputImg3[21],
                      OutputImg3[20],OutputImg3[19],OutputImg3[18],
                      OutputImg3[17],OutputImg3[16]}), .EN (nx23788), .F ({
                      ImgReg2IN_31,ImgReg2IN_30,ImgReg2IN_29,ImgReg2IN_28,
                      ImgReg2IN_27,ImgReg2IN_26,ImgReg2IN_25,ImgReg2IN_24,
                      ImgReg2IN_23,ImgReg2IN_22,ImgReg2IN_21,ImgReg2IN_20,
                      ImgReg2IN_19,ImgReg2IN_18,ImgReg2IN_17,ImgReg2IN_16})) ;
    triStateBuffer_16 loop3_1_TriState3U (.D ({OutputImg4[31],OutputImg4[30],
                      OutputImg4[29],OutputImg4[28],OutputImg4[27],
                      OutputImg4[26],OutputImg4[25],OutputImg4[24],
                      OutputImg4[23],OutputImg4[22],OutputImg4[21],
                      OutputImg4[20],OutputImg4[19],OutputImg4[18],
                      OutputImg4[17],OutputImg4[16]}), .EN (nx23788), .F ({
                      ImgReg3IN_31,ImgReg3IN_30,ImgReg3IN_29,ImgReg3IN_28,
                      ImgReg3IN_27,ImgReg3IN_26,ImgReg3IN_25,ImgReg3IN_24,
                      ImgReg3IN_23,ImgReg3IN_22,ImgReg3IN_21,ImgReg3IN_20,
                      ImgReg3IN_19,ImgReg3IN_18,ImgReg3IN_17,ImgReg3IN_16})) ;
    triStateBuffer_16 loop3_1_TriState4U (.D ({OutputImg5[31],OutputImg5[30],
                      OutputImg5[29],OutputImg5[28],OutputImg5[27],
                      OutputImg5[26],OutputImg5[25],OutputImg5[24],
                      OutputImg5[23],OutputImg5[22],OutputImg5[21],
                      OutputImg5[20],OutputImg5[19],OutputImg5[18],
                      OutputImg5[17],OutputImg5[16]}), .EN (nx23788), .F ({
                      ImgReg4IN_31,ImgReg4IN_30,ImgReg4IN_29,ImgReg4IN_28,
                      ImgReg4IN_27,ImgReg4IN_26,ImgReg4IN_25,ImgReg4IN_24,
                      ImgReg4IN_23,ImgReg4IN_22,ImgReg4IN_21,ImgReg4IN_20,
                      ImgReg4IN_19,ImgReg4IN_18,ImgReg4IN_17,ImgReg4IN_16})) ;
    nBitRegister_16 loop3_1_reg1 (.D ({ImgReg0IN_31,ImgReg0IN_30,ImgReg0IN_29,
                    ImgReg0IN_28,ImgReg0IN_27,ImgReg0IN_26,ImgReg0IN_25,
                    ImgReg0IN_24,ImgReg0IN_23,ImgReg0IN_22,ImgReg0IN_21,
                    ImgReg0IN_20,ImgReg0IN_19,ImgReg0IN_18,ImgReg0IN_17,
                    ImgReg0IN_16}), .CLK (nx23834), .RST (RST), .EN (nx23718), .Q (
                    {OutputImg0[31],OutputImg0[30],OutputImg0[29],OutputImg0[28]
                    ,OutputImg0[27],OutputImg0[26],OutputImg0[25],OutputImg0[24]
                    ,OutputImg0[23],OutputImg0[22],OutputImg0[21],OutputImg0[20]
                    ,OutputImg0[19],OutputImg0[18],OutputImg0[17],OutputImg0[16]
                    })) ;
    nBitRegister_16 loop3_1_reg2 (.D ({ImgReg1IN_31,ImgReg1IN_30,ImgReg1IN_29,
                    ImgReg1IN_28,ImgReg1IN_27,ImgReg1IN_26,ImgReg1IN_25,
                    ImgReg1IN_24,ImgReg1IN_23,ImgReg1IN_22,ImgReg1IN_21,
                    ImgReg1IN_20,ImgReg1IN_19,ImgReg1IN_18,ImgReg1IN_17,
                    ImgReg1IN_16}), .CLK (nx23836), .RST (RST), .EN (nx23728), .Q (
                    {OutputImg1[31],OutputImg1[30],OutputImg1[29],OutputImg1[28]
                    ,OutputImg1[27],OutputImg1[26],OutputImg1[25],OutputImg1[24]
                    ,OutputImg1[23],OutputImg1[22],OutputImg1[21],OutputImg1[20]
                    ,OutputImg1[19],OutputImg1[18],OutputImg1[17],OutputImg1[16]
                    })) ;
    nBitRegister_16 loop3_1_reg3 (.D ({ImgReg2IN_31,ImgReg2IN_30,ImgReg2IN_29,
                    ImgReg2IN_28,ImgReg2IN_27,ImgReg2IN_26,ImgReg2IN_25,
                    ImgReg2IN_24,ImgReg2IN_23,ImgReg2IN_22,ImgReg2IN_21,
                    ImgReg2IN_20,ImgReg2IN_19,ImgReg2IN_18,ImgReg2IN_17,
                    ImgReg2IN_16}), .CLK (nx23836), .RST (RST), .EN (nx23738), .Q (
                    {OutputImg2[31],OutputImg2[30],OutputImg2[29],OutputImg2[28]
                    ,OutputImg2[27],OutputImg2[26],OutputImg2[25],OutputImg2[24]
                    ,OutputImg2[23],OutputImg2[22],OutputImg2[21],OutputImg2[20]
                    ,OutputImg2[19],OutputImg2[18],OutputImg2[17],OutputImg2[16]
                    })) ;
    nBitRegister_16 loop3_1_reg4 (.D ({ImgReg3IN_31,ImgReg3IN_30,ImgReg3IN_29,
                    ImgReg3IN_28,ImgReg3IN_27,ImgReg3IN_26,ImgReg3IN_25,
                    ImgReg3IN_24,ImgReg3IN_23,ImgReg3IN_22,ImgReg3IN_21,
                    ImgReg3IN_20,ImgReg3IN_19,ImgReg3IN_18,ImgReg3IN_17,
                    ImgReg3IN_16}), .CLK (nx23838), .RST (RST), .EN (nx23748), .Q (
                    {OutputImg3[31],OutputImg3[30],OutputImg3[29],OutputImg3[28]
                    ,OutputImg3[27],OutputImg3[26],OutputImg3[25],OutputImg3[24]
                    ,OutputImg3[23],OutputImg3[22],OutputImg3[21],OutputImg3[20]
                    ,OutputImg3[19],OutputImg3[18],OutputImg3[17],OutputImg3[16]
                    })) ;
    nBitRegister_16 loop3_1_reg5 (.D ({ImgReg4IN_31,ImgReg4IN_30,ImgReg4IN_29,
                    ImgReg4IN_28,ImgReg4IN_27,ImgReg4IN_26,ImgReg4IN_25,
                    ImgReg4IN_24,ImgReg4IN_23,ImgReg4IN_22,ImgReg4IN_21,
                    ImgReg4IN_20,ImgReg4IN_19,ImgReg4IN_18,ImgReg4IN_17,
                    ImgReg4IN_16}), .CLK (nx23838), .RST (RST), .EN (nx23758), .Q (
                    {OutputImg4[31],OutputImg4[30],OutputImg4[29],OutputImg4[28]
                    ,OutputImg4[27],OutputImg4[26],OutputImg4[25],OutputImg4[24]
                    ,OutputImg4[23],OutputImg4[22],OutputImg4[21],OutputImg4[20]
                    ,OutputImg4[19],OutputImg4[18],OutputImg4[17],OutputImg4[16]
                    })) ;
    nBitRegister_16 loop3_1_reg6 (.D ({ImgReg5IN_31,ImgReg5IN_30,ImgReg5IN_29,
                    ImgReg5IN_28,ImgReg5IN_27,ImgReg5IN_26,ImgReg5IN_25,
                    ImgReg5IN_24,ImgReg5IN_23,ImgReg5IN_22,ImgReg5IN_21,
                    ImgReg5IN_20,ImgReg5IN_19,ImgReg5IN_18,ImgReg5IN_17,
                    ImgReg5IN_16}), .CLK (nx23840), .RST (RST), .EN (nx23768), .Q (
                    {OutputImg5[31],OutputImg5[30],OutputImg5[29],OutputImg5[28]
                    ,OutputImg5[27],OutputImg5[26],OutputImg5[25],OutputImg5[24]
                    ,OutputImg5[23],OutputImg5[22],OutputImg5[21],OutputImg5[20]
                    ,OutputImg5[19],OutputImg5[18],OutputImg5[17],OutputImg5[16]
                    })) ;
    triStateBuffer_16 loop3_2_TriState0L (.D ({OutputImg0[63],OutputImg0[62],
                      OutputImg0[61],OutputImg0[60],OutputImg0[59],
                      OutputImg0[58],OutputImg0[57],OutputImg0[56],
                      OutputImg0[55],OutputImg0[54],OutputImg0[53],
                      OutputImg0[52],OutputImg0[51],OutputImg0[50],
                      OutputImg0[49],OutputImg0[48]}), .EN (nx23668), .F ({
                      ImgReg0IN_47,ImgReg0IN_46,ImgReg0IN_45,ImgReg0IN_44,
                      ImgReg0IN_43,ImgReg0IN_42,ImgReg0IN_41,ImgReg0IN_40,
                      ImgReg0IN_39,ImgReg0IN_38,ImgReg0IN_37,ImgReg0IN_36,
                      ImgReg0IN_35,ImgReg0IN_34,ImgReg0IN_33,ImgReg0IN_32})) ;
    triStateBuffer_16 loop3_2_TriState1L (.D ({OutputImg1[63],OutputImg1[62],
                      OutputImg1[61],OutputImg1[60],OutputImg1[59],
                      OutputImg1[58],OutputImg1[57],OutputImg1[56],
                      OutputImg1[55],OutputImg1[54],OutputImg1[53],
                      OutputImg1[52],OutputImg1[51],OutputImg1[50],
                      OutputImg1[49],OutputImg1[48]}), .EN (nx23668), .F ({
                      ImgReg1IN_47,ImgReg1IN_46,ImgReg1IN_45,ImgReg1IN_44,
                      ImgReg1IN_43,ImgReg1IN_42,ImgReg1IN_41,ImgReg1IN_40,
                      ImgReg1IN_39,ImgReg1IN_38,ImgReg1IN_37,ImgReg1IN_36,
                      ImgReg1IN_35,ImgReg1IN_34,ImgReg1IN_33,ImgReg1IN_32})) ;
    triStateBuffer_16 loop3_2_TriState2L (.D ({OutputImg2[63],OutputImg2[62],
                      OutputImg2[61],OutputImg2[60],OutputImg2[59],
                      OutputImg2[58],OutputImg2[57],OutputImg2[56],
                      OutputImg2[55],OutputImg2[54],OutputImg2[53],
                      OutputImg2[52],OutputImg2[51],OutputImg2[50],
                      OutputImg2[49],OutputImg2[48]}), .EN (nx23670), .F ({
                      ImgReg2IN_47,ImgReg2IN_46,ImgReg2IN_45,ImgReg2IN_44,
                      ImgReg2IN_43,ImgReg2IN_42,ImgReg2IN_41,ImgReg2IN_40,
                      ImgReg2IN_39,ImgReg2IN_38,ImgReg2IN_37,ImgReg2IN_36,
                      ImgReg2IN_35,ImgReg2IN_34,ImgReg2IN_33,ImgReg2IN_32})) ;
    triStateBuffer_16 loop3_2_TriState3L (.D ({OutputImg3[63],OutputImg3[62],
                      OutputImg3[61],OutputImg3[60],OutputImg3[59],
                      OutputImg3[58],OutputImg3[57],OutputImg3[56],
                      OutputImg3[55],OutputImg3[54],OutputImg3[53],
                      OutputImg3[52],OutputImg3[51],OutputImg3[50],
                      OutputImg3[49],OutputImg3[48]}), .EN (nx23670), .F ({
                      ImgReg3IN_47,ImgReg3IN_46,ImgReg3IN_45,ImgReg3IN_44,
                      ImgReg3IN_43,ImgReg3IN_42,ImgReg3IN_41,ImgReg3IN_40,
                      ImgReg3IN_39,ImgReg3IN_38,ImgReg3IN_37,ImgReg3IN_36,
                      ImgReg3IN_35,ImgReg3IN_34,ImgReg3IN_33,ImgReg3IN_32})) ;
    triStateBuffer_16 loop3_2_TriState4L (.D ({OutputImg4[63],OutputImg4[62],
                      OutputImg4[61],OutputImg4[60],OutputImg4[59],
                      OutputImg4[58],OutputImg4[57],OutputImg4[56],
                      OutputImg4[55],OutputImg4[54],OutputImg4[53],
                      OutputImg4[52],OutputImg4[51],OutputImg4[50],
                      OutputImg4[49],OutputImg4[48]}), .EN (nx23670), .F ({
                      ImgReg4IN_47,ImgReg4IN_46,ImgReg4IN_45,ImgReg4IN_44,
                      ImgReg4IN_43,ImgReg4IN_42,ImgReg4IN_41,ImgReg4IN_40,
                      ImgReg4IN_39,ImgReg4IN_38,ImgReg4IN_37,ImgReg4IN_36,
                      ImgReg4IN_35,ImgReg4IN_34,ImgReg4IN_33,ImgReg4IN_32})) ;
    triStateBuffer_16 loop3_2_TriState5L (.D ({OutputImg5[63],OutputImg5[62],
                      OutputImg5[61],OutputImg5[60],OutputImg5[59],
                      OutputImg5[58],OutputImg5[57],OutputImg5[56],
                      OutputImg5[55],OutputImg5[54],OutputImg5[53],
                      OutputImg5[52],OutputImg5[51],OutputImg5[50],
                      OutputImg5[49],OutputImg5[48]}), .EN (nx23670), .F ({
                      ImgReg5IN_47,ImgReg5IN_46,ImgReg5IN_45,ImgReg5IN_44,
                      ImgReg5IN_43,ImgReg5IN_42,ImgReg5IN_41,ImgReg5IN_40,
                      ImgReg5IN_39,ImgReg5IN_38,ImgReg5IN_37,ImgReg5IN_36,
                      ImgReg5IN_35,ImgReg5IN_34,ImgReg5IN_33,ImgReg5IN_32})) ;
    triStateBuffer_16 loop3_2_TriState0N (.D ({DATA[47],DATA[46],DATA[45],
                      DATA[44],DATA[43],DATA[42],DATA[41],DATA[40],DATA[39],
                      DATA[38],DATA[37],DATA[36],DATA[35],DATA[34],DATA[33],
                      DATA[32]}), .EN (nx23654), .F ({ImgReg0IN_47,ImgReg0IN_46,
                      ImgReg0IN_45,ImgReg0IN_44,ImgReg0IN_43,ImgReg0IN_42,
                      ImgReg0IN_41,ImgReg0IN_40,ImgReg0IN_39,ImgReg0IN_38,
                      ImgReg0IN_37,ImgReg0IN_36,ImgReg0IN_35,ImgReg0IN_34,
                      ImgReg0IN_33,ImgReg0IN_32})) ;
    triStateBuffer_16 loop3_2_TriState1N (.D ({DATA[47],DATA[46],DATA[45],
                      DATA[44],DATA[43],DATA[42],DATA[41],DATA[40],DATA[39],
                      DATA[38],DATA[37],DATA[36],DATA[35],DATA[34],DATA[33],
                      DATA[32]}), .EN (nx23642), .F ({ImgReg1IN_47,ImgReg1IN_46,
                      ImgReg1IN_45,ImgReg1IN_44,ImgReg1IN_43,ImgReg1IN_42,
                      ImgReg1IN_41,ImgReg1IN_40,ImgReg1IN_39,ImgReg1IN_38,
                      ImgReg1IN_37,ImgReg1IN_36,ImgReg1IN_35,ImgReg1IN_34,
                      ImgReg1IN_33,ImgReg1IN_32})) ;
    triStateBuffer_16 loop3_2_TriState2N (.D ({DATA[47],DATA[46],DATA[45],
                      DATA[44],DATA[43],DATA[42],DATA[41],DATA[40],DATA[39],
                      DATA[38],DATA[37],DATA[36],DATA[35],DATA[34],DATA[33],
                      DATA[32]}), .EN (nx23630), .F ({ImgReg2IN_47,ImgReg2IN_46,
                      ImgReg2IN_45,ImgReg2IN_44,ImgReg2IN_43,ImgReg2IN_42,
                      ImgReg2IN_41,ImgReg2IN_40,ImgReg2IN_39,ImgReg2IN_38,
                      ImgReg2IN_37,ImgReg2IN_36,ImgReg2IN_35,ImgReg2IN_34,
                      ImgReg2IN_33,ImgReg2IN_32})) ;
    triStateBuffer_16 loop3_2_TriState3N (.D ({DATA[47],DATA[46],DATA[45],
                      DATA[44],DATA[43],DATA[42],DATA[41],DATA[40],DATA[39],
                      DATA[38],DATA[37],DATA[36],DATA[35],DATA[34],DATA[33],
                      DATA[32]}), .EN (nx23618), .F ({ImgReg3IN_47,ImgReg3IN_46,
                      ImgReg3IN_45,ImgReg3IN_44,ImgReg3IN_43,ImgReg3IN_42,
                      ImgReg3IN_41,ImgReg3IN_40,ImgReg3IN_39,ImgReg3IN_38,
                      ImgReg3IN_37,ImgReg3IN_36,ImgReg3IN_35,ImgReg3IN_34,
                      ImgReg3IN_33,ImgReg3IN_32})) ;
    triStateBuffer_16 loop3_2_TriState4N (.D ({DATA[47],DATA[46],DATA[45],
                      DATA[44],DATA[43],DATA[42],DATA[41],DATA[40],DATA[39],
                      DATA[38],DATA[37],DATA[36],DATA[35],DATA[34],DATA[33],
                      DATA[32]}), .EN (nx23606), .F ({ImgReg4IN_47,ImgReg4IN_46,
                      ImgReg4IN_45,ImgReg4IN_44,ImgReg4IN_43,ImgReg4IN_42,
                      ImgReg4IN_41,ImgReg4IN_40,ImgReg4IN_39,ImgReg4IN_38,
                      ImgReg4IN_37,ImgReg4IN_36,ImgReg4IN_35,ImgReg4IN_34,
                      ImgReg4IN_33,ImgReg4IN_32})) ;
    triStateBuffer_16 loop3_2_TriState5N (.D ({DATA[47],DATA[46],DATA[45],
                      DATA[44],DATA[43],DATA[42],DATA[41],DATA[40],DATA[39],
                      DATA[38],DATA[37],DATA[36],DATA[35],DATA[34],DATA[33],
                      DATA[32]}), .EN (nx23594), .F ({ImgReg5IN_47,ImgReg5IN_46,
                      ImgReg5IN_45,ImgReg5IN_44,ImgReg5IN_43,ImgReg5IN_42,
                      ImgReg5IN_41,ImgReg5IN_40,ImgReg5IN_39,ImgReg5IN_38,
                      ImgReg5IN_37,ImgReg5IN_36,ImgReg5IN_35,ImgReg5IN_34,
                      ImgReg5IN_33,ImgReg5IN_32})) ;
    triStateBuffer_16 loop3_2_TriState0U (.D ({OutputImg1[47],OutputImg1[46],
                      OutputImg1[45],OutputImg1[44],OutputImg1[43],
                      OutputImg1[42],OutputImg1[41],OutputImg1[40],
                      OutputImg1[39],OutputImg1[38],OutputImg1[37],
                      OutputImg1[36],OutputImg1[35],OutputImg1[34],
                      OutputImg1[33],OutputImg1[32]}), .EN (nx23788), .F ({
                      ImgReg0IN_47,ImgReg0IN_46,ImgReg0IN_45,ImgReg0IN_44,
                      ImgReg0IN_43,ImgReg0IN_42,ImgReg0IN_41,ImgReg0IN_40,
                      ImgReg0IN_39,ImgReg0IN_38,ImgReg0IN_37,ImgReg0IN_36,
                      ImgReg0IN_35,ImgReg0IN_34,ImgReg0IN_33,ImgReg0IN_32})) ;
    triStateBuffer_16 loop3_2_TriState1U (.D ({OutputImg2[47],OutputImg2[46],
                      OutputImg2[45],OutputImg2[44],OutputImg2[43],
                      OutputImg2[42],OutputImg2[41],OutputImg2[40],
                      OutputImg2[39],OutputImg2[38],OutputImg2[37],
                      OutputImg2[36],OutputImg2[35],OutputImg2[34],
                      OutputImg2[33],OutputImg2[32]}), .EN (nx23788), .F ({
                      ImgReg1IN_47,ImgReg1IN_46,ImgReg1IN_45,ImgReg1IN_44,
                      ImgReg1IN_43,ImgReg1IN_42,ImgReg1IN_41,ImgReg1IN_40,
                      ImgReg1IN_39,ImgReg1IN_38,ImgReg1IN_37,ImgReg1IN_36,
                      ImgReg1IN_35,ImgReg1IN_34,ImgReg1IN_33,ImgReg1IN_32})) ;
    triStateBuffer_16 loop3_2_TriState2U (.D ({OutputImg3[47],OutputImg3[46],
                      OutputImg3[45],OutputImg3[44],OutputImg3[43],
                      OutputImg3[42],OutputImg3[41],OutputImg3[40],
                      OutputImg3[39],OutputImg3[38],OutputImg3[37],
                      OutputImg3[36],OutputImg3[35],OutputImg3[34],
                      OutputImg3[33],OutputImg3[32]}), .EN (nx23788), .F ({
                      ImgReg2IN_47,ImgReg2IN_46,ImgReg2IN_45,ImgReg2IN_44,
                      ImgReg2IN_43,ImgReg2IN_42,ImgReg2IN_41,ImgReg2IN_40,
                      ImgReg2IN_39,ImgReg2IN_38,ImgReg2IN_37,ImgReg2IN_36,
                      ImgReg2IN_35,ImgReg2IN_34,ImgReg2IN_33,ImgReg2IN_32})) ;
    triStateBuffer_16 loop3_2_TriState3U (.D ({OutputImg4[47],OutputImg4[46],
                      OutputImg4[45],OutputImg4[44],OutputImg4[43],
                      OutputImg4[42],OutputImg4[41],OutputImg4[40],
                      OutputImg4[39],OutputImg4[38],OutputImg4[37],
                      OutputImg4[36],OutputImg4[35],OutputImg4[34],
                      OutputImg4[33],OutputImg4[32]}), .EN (nx23788), .F ({
                      ImgReg3IN_47,ImgReg3IN_46,ImgReg3IN_45,ImgReg3IN_44,
                      ImgReg3IN_43,ImgReg3IN_42,ImgReg3IN_41,ImgReg3IN_40,
                      ImgReg3IN_39,ImgReg3IN_38,ImgReg3IN_37,ImgReg3IN_36,
                      ImgReg3IN_35,ImgReg3IN_34,ImgReg3IN_33,ImgReg3IN_32})) ;
    triStateBuffer_16 loop3_2_TriState4U (.D ({OutputImg5[47],OutputImg5[46],
                      OutputImg5[45],OutputImg5[44],OutputImg5[43],
                      OutputImg5[42],OutputImg5[41],OutputImg5[40],
                      OutputImg5[39],OutputImg5[38],OutputImg5[37],
                      OutputImg5[36],OutputImg5[35],OutputImg5[34],
                      OutputImg5[33],OutputImg5[32]}), .EN (nx23790), .F ({
                      ImgReg4IN_47,ImgReg4IN_46,ImgReg4IN_45,ImgReg4IN_44,
                      ImgReg4IN_43,ImgReg4IN_42,ImgReg4IN_41,ImgReg4IN_40,
                      ImgReg4IN_39,ImgReg4IN_38,ImgReg4IN_37,ImgReg4IN_36,
                      ImgReg4IN_35,ImgReg4IN_34,ImgReg4IN_33,ImgReg4IN_32})) ;
    nBitRegister_16 loop3_2_reg1 (.D ({ImgReg0IN_47,ImgReg0IN_46,ImgReg0IN_45,
                    ImgReg0IN_44,ImgReg0IN_43,ImgReg0IN_42,ImgReg0IN_41,
                    ImgReg0IN_40,ImgReg0IN_39,ImgReg0IN_38,ImgReg0IN_37,
                    ImgReg0IN_36,ImgReg0IN_35,ImgReg0IN_34,ImgReg0IN_33,
                    ImgReg0IN_32}), .CLK (nx23840), .RST (RST), .EN (nx23718), .Q (
                    {OutputImg0[47],OutputImg0[46],OutputImg0[45],OutputImg0[44]
                    ,OutputImg0[43],OutputImg0[42],OutputImg0[41],OutputImg0[40]
                    ,OutputImg0[39],OutputImg0[38],OutputImg0[37],OutputImg0[36]
                    ,OutputImg0[35],OutputImg0[34],OutputImg0[33],OutputImg0[32]
                    })) ;
    nBitRegister_16 loop3_2_reg2 (.D ({ImgReg1IN_47,ImgReg1IN_46,ImgReg1IN_45,
                    ImgReg1IN_44,ImgReg1IN_43,ImgReg1IN_42,ImgReg1IN_41,
                    ImgReg1IN_40,ImgReg1IN_39,ImgReg1IN_38,ImgReg1IN_37,
                    ImgReg1IN_36,ImgReg1IN_35,ImgReg1IN_34,ImgReg1IN_33,
                    ImgReg1IN_32}), .CLK (nx23842), .RST (RST), .EN (nx23728), .Q (
                    {OutputImg1[47],OutputImg1[46],OutputImg1[45],OutputImg1[44]
                    ,OutputImg1[43],OutputImg1[42],OutputImg1[41],OutputImg1[40]
                    ,OutputImg1[39],OutputImg1[38],OutputImg1[37],OutputImg1[36]
                    ,OutputImg1[35],OutputImg1[34],OutputImg1[33],OutputImg1[32]
                    })) ;
    nBitRegister_16 loop3_2_reg3 (.D ({ImgReg2IN_47,ImgReg2IN_46,ImgReg2IN_45,
                    ImgReg2IN_44,ImgReg2IN_43,ImgReg2IN_42,ImgReg2IN_41,
                    ImgReg2IN_40,ImgReg2IN_39,ImgReg2IN_38,ImgReg2IN_37,
                    ImgReg2IN_36,ImgReg2IN_35,ImgReg2IN_34,ImgReg2IN_33,
                    ImgReg2IN_32}), .CLK (nx23842), .RST (RST), .EN (nx23738), .Q (
                    {OutputImg2[47],OutputImg2[46],OutputImg2[45],OutputImg2[44]
                    ,OutputImg2[43],OutputImg2[42],OutputImg2[41],OutputImg2[40]
                    ,OutputImg2[39],OutputImg2[38],OutputImg2[37],OutputImg2[36]
                    ,OutputImg2[35],OutputImg2[34],OutputImg2[33],OutputImg2[32]
                    })) ;
    nBitRegister_16 loop3_2_reg4 (.D ({ImgReg3IN_47,ImgReg3IN_46,ImgReg3IN_45,
                    ImgReg3IN_44,ImgReg3IN_43,ImgReg3IN_42,ImgReg3IN_41,
                    ImgReg3IN_40,ImgReg3IN_39,ImgReg3IN_38,ImgReg3IN_37,
                    ImgReg3IN_36,ImgReg3IN_35,ImgReg3IN_34,ImgReg3IN_33,
                    ImgReg3IN_32}), .CLK (nx23844), .RST (RST), .EN (nx23748), .Q (
                    {OutputImg3[47],OutputImg3[46],OutputImg3[45],OutputImg3[44]
                    ,OutputImg3[43],OutputImg3[42],OutputImg3[41],OutputImg3[40]
                    ,OutputImg3[39],OutputImg3[38],OutputImg3[37],OutputImg3[36]
                    ,OutputImg3[35],OutputImg3[34],OutputImg3[33],OutputImg3[32]
                    })) ;
    nBitRegister_16 loop3_2_reg5 (.D ({ImgReg4IN_47,ImgReg4IN_46,ImgReg4IN_45,
                    ImgReg4IN_44,ImgReg4IN_43,ImgReg4IN_42,ImgReg4IN_41,
                    ImgReg4IN_40,ImgReg4IN_39,ImgReg4IN_38,ImgReg4IN_37,
                    ImgReg4IN_36,ImgReg4IN_35,ImgReg4IN_34,ImgReg4IN_33,
                    ImgReg4IN_32}), .CLK (nx23844), .RST (RST), .EN (nx23758), .Q (
                    {OutputImg4[47],OutputImg4[46],OutputImg4[45],OutputImg4[44]
                    ,OutputImg4[43],OutputImg4[42],OutputImg4[41],OutputImg4[40]
                    ,OutputImg4[39],OutputImg4[38],OutputImg4[37],OutputImg4[36]
                    ,OutputImg4[35],OutputImg4[34],OutputImg4[33],OutputImg4[32]
                    })) ;
    nBitRegister_16 loop3_2_reg6 (.D ({ImgReg5IN_47,ImgReg5IN_46,ImgReg5IN_45,
                    ImgReg5IN_44,ImgReg5IN_43,ImgReg5IN_42,ImgReg5IN_41,
                    ImgReg5IN_40,ImgReg5IN_39,ImgReg5IN_38,ImgReg5IN_37,
                    ImgReg5IN_36,ImgReg5IN_35,ImgReg5IN_34,ImgReg5IN_33,
                    ImgReg5IN_32}), .CLK (nx23846), .RST (RST), .EN (nx23768), .Q (
                    {OutputImg5[47],OutputImg5[46],OutputImg5[45],OutputImg5[44]
                    ,OutputImg5[43],OutputImg5[42],OutputImg5[41],OutputImg5[40]
                    ,OutputImg5[39],OutputImg5[38],OutputImg5[37],OutputImg5[36]
                    ,OutputImg5[35],OutputImg5[34],OutputImg5[33],OutputImg5[32]
                    })) ;
    triStateBuffer_16 loop3_3_TriState0L (.D ({OutputImg0[79],OutputImg0[78],
                      OutputImg0[77],OutputImg0[76],OutputImg0[75],
                      OutputImg0[74],OutputImg0[73],OutputImg0[72],
                      OutputImg0[71],OutputImg0[70],OutputImg0[69],
                      OutputImg0[68],OutputImg0[67],OutputImg0[66],
                      OutputImg0[65],OutputImg0[64]}), .EN (nx23670), .F ({
                      ImgReg0IN_63,ImgReg0IN_62,ImgReg0IN_61,ImgReg0IN_60,
                      ImgReg0IN_59,ImgReg0IN_58,ImgReg0IN_57,ImgReg0IN_56,
                      ImgReg0IN_55,ImgReg0IN_54,ImgReg0IN_53,ImgReg0IN_52,
                      ImgReg0IN_51,ImgReg0IN_50,ImgReg0IN_49,ImgReg0IN_48})) ;
    triStateBuffer_16 loop3_3_TriState1L (.D ({OutputImg1[79],OutputImg1[78],
                      OutputImg1[77],OutputImg1[76],OutputImg1[75],
                      OutputImg1[74],OutputImg1[73],OutputImg1[72],
                      OutputImg1[71],OutputImg1[70],OutputImg1[69],
                      OutputImg1[68],OutputImg1[67],OutputImg1[66],
                      OutputImg1[65],OutputImg1[64]}), .EN (nx23670), .F ({
                      ImgReg1IN_63,ImgReg1IN_62,ImgReg1IN_61,ImgReg1IN_60,
                      ImgReg1IN_59,ImgReg1IN_58,ImgReg1IN_57,ImgReg1IN_56,
                      ImgReg1IN_55,ImgReg1IN_54,ImgReg1IN_53,ImgReg1IN_52,
                      ImgReg1IN_51,ImgReg1IN_50,ImgReg1IN_49,ImgReg1IN_48})) ;
    triStateBuffer_16 loop3_3_TriState2L (.D ({OutputImg2[79],OutputImg2[78],
                      OutputImg2[77],OutputImg2[76],OutputImg2[75],
                      OutputImg2[74],OutputImg2[73],OutputImg2[72],
                      OutputImg2[71],OutputImg2[70],OutputImg2[69],
                      OutputImg2[68],OutputImg2[67],OutputImg2[66],
                      OutputImg2[65],OutputImg2[64]}), .EN (nx23670), .F ({
                      ImgReg2IN_63,ImgReg2IN_62,ImgReg2IN_61,ImgReg2IN_60,
                      ImgReg2IN_59,ImgReg2IN_58,ImgReg2IN_57,ImgReg2IN_56,
                      ImgReg2IN_55,ImgReg2IN_54,ImgReg2IN_53,ImgReg2IN_52,
                      ImgReg2IN_51,ImgReg2IN_50,ImgReg2IN_49,ImgReg2IN_48})) ;
    triStateBuffer_16 loop3_3_TriState3L (.D ({OutputImg3[79],OutputImg3[78],
                      OutputImg3[77],OutputImg3[76],OutputImg3[75],
                      OutputImg3[74],OutputImg3[73],OutputImg3[72],
                      OutputImg3[71],OutputImg3[70],OutputImg3[69],
                      OutputImg3[68],OutputImg3[67],OutputImg3[66],
                      OutputImg3[65],OutputImg3[64]}), .EN (nx23672), .F ({
                      ImgReg3IN_63,ImgReg3IN_62,ImgReg3IN_61,ImgReg3IN_60,
                      ImgReg3IN_59,ImgReg3IN_58,ImgReg3IN_57,ImgReg3IN_56,
                      ImgReg3IN_55,ImgReg3IN_54,ImgReg3IN_53,ImgReg3IN_52,
                      ImgReg3IN_51,ImgReg3IN_50,ImgReg3IN_49,ImgReg3IN_48})) ;
    triStateBuffer_16 loop3_3_TriState4L (.D ({OutputImg4[79],OutputImg4[78],
                      OutputImg4[77],OutputImg4[76],OutputImg4[75],
                      OutputImg4[74],OutputImg4[73],OutputImg4[72],
                      OutputImg4[71],OutputImg4[70],OutputImg4[69],
                      OutputImg4[68],OutputImg4[67],OutputImg4[66],
                      OutputImg4[65],OutputImg4[64]}), .EN (nx23672), .F ({
                      ImgReg4IN_63,ImgReg4IN_62,ImgReg4IN_61,ImgReg4IN_60,
                      ImgReg4IN_59,ImgReg4IN_58,ImgReg4IN_57,ImgReg4IN_56,
                      ImgReg4IN_55,ImgReg4IN_54,ImgReg4IN_53,ImgReg4IN_52,
                      ImgReg4IN_51,ImgReg4IN_50,ImgReg4IN_49,ImgReg4IN_48})) ;
    triStateBuffer_16 loop3_3_TriState5L (.D ({OutputImg5[79],OutputImg5[78],
                      OutputImg5[77],OutputImg5[76],OutputImg5[75],
                      OutputImg5[74],OutputImg5[73],OutputImg5[72],
                      OutputImg5[71],OutputImg5[70],OutputImg5[69],
                      OutputImg5[68],OutputImg5[67],OutputImg5[66],
                      OutputImg5[65],OutputImg5[64]}), .EN (nx23672), .F ({
                      ImgReg5IN_63,ImgReg5IN_62,ImgReg5IN_61,ImgReg5IN_60,
                      ImgReg5IN_59,ImgReg5IN_58,ImgReg5IN_57,ImgReg5IN_56,
                      ImgReg5IN_55,ImgReg5IN_54,ImgReg5IN_53,ImgReg5IN_52,
                      ImgReg5IN_51,ImgReg5IN_50,ImgReg5IN_49,ImgReg5IN_48})) ;
    triStateBuffer_16 loop3_3_TriState0N (.D ({DATA[63],DATA[62],DATA[61],
                      DATA[60],DATA[59],DATA[58],DATA[57],DATA[56],DATA[55],
                      DATA[54],DATA[53],DATA[52],DATA[51],DATA[50],DATA[49],
                      DATA[48]}), .EN (nx23654), .F ({ImgReg0IN_63,ImgReg0IN_62,
                      ImgReg0IN_61,ImgReg0IN_60,ImgReg0IN_59,ImgReg0IN_58,
                      ImgReg0IN_57,ImgReg0IN_56,ImgReg0IN_55,ImgReg0IN_54,
                      ImgReg0IN_53,ImgReg0IN_52,ImgReg0IN_51,ImgReg0IN_50,
                      ImgReg0IN_49,ImgReg0IN_48})) ;
    triStateBuffer_16 loop3_3_TriState1N (.D ({DATA[63],DATA[62],DATA[61],
                      DATA[60],DATA[59],DATA[58],DATA[57],DATA[56],DATA[55],
                      DATA[54],DATA[53],DATA[52],DATA[51],DATA[50],DATA[49],
                      DATA[48]}), .EN (nx23642), .F ({ImgReg1IN_63,ImgReg1IN_62,
                      ImgReg1IN_61,ImgReg1IN_60,ImgReg1IN_59,ImgReg1IN_58,
                      ImgReg1IN_57,ImgReg1IN_56,ImgReg1IN_55,ImgReg1IN_54,
                      ImgReg1IN_53,ImgReg1IN_52,ImgReg1IN_51,ImgReg1IN_50,
                      ImgReg1IN_49,ImgReg1IN_48})) ;
    triStateBuffer_16 loop3_3_TriState2N (.D ({DATA[63],DATA[62],DATA[61],
                      DATA[60],DATA[59],DATA[58],DATA[57],DATA[56],DATA[55],
                      DATA[54],DATA[53],DATA[52],DATA[51],DATA[50],DATA[49],
                      DATA[48]}), .EN (nx23630), .F ({ImgReg2IN_63,ImgReg2IN_62,
                      ImgReg2IN_61,ImgReg2IN_60,ImgReg2IN_59,ImgReg2IN_58,
                      ImgReg2IN_57,ImgReg2IN_56,ImgReg2IN_55,ImgReg2IN_54,
                      ImgReg2IN_53,ImgReg2IN_52,ImgReg2IN_51,ImgReg2IN_50,
                      ImgReg2IN_49,ImgReg2IN_48})) ;
    triStateBuffer_16 loop3_3_TriState3N (.D ({DATA[63],DATA[62],DATA[61],
                      DATA[60],DATA[59],DATA[58],DATA[57],DATA[56],DATA[55],
                      DATA[54],DATA[53],DATA[52],DATA[51],DATA[50],DATA[49],
                      DATA[48]}), .EN (nx23618), .F ({ImgReg3IN_63,ImgReg3IN_62,
                      ImgReg3IN_61,ImgReg3IN_60,ImgReg3IN_59,ImgReg3IN_58,
                      ImgReg3IN_57,ImgReg3IN_56,ImgReg3IN_55,ImgReg3IN_54,
                      ImgReg3IN_53,ImgReg3IN_52,ImgReg3IN_51,ImgReg3IN_50,
                      ImgReg3IN_49,ImgReg3IN_48})) ;
    triStateBuffer_16 loop3_3_TriState4N (.D ({DATA[63],DATA[62],DATA[61],
                      DATA[60],DATA[59],DATA[58],DATA[57],DATA[56],DATA[55],
                      DATA[54],DATA[53],DATA[52],DATA[51],DATA[50],DATA[49],
                      DATA[48]}), .EN (nx23606), .F ({ImgReg4IN_63,ImgReg4IN_62,
                      ImgReg4IN_61,ImgReg4IN_60,ImgReg4IN_59,ImgReg4IN_58,
                      ImgReg4IN_57,ImgReg4IN_56,ImgReg4IN_55,ImgReg4IN_54,
                      ImgReg4IN_53,ImgReg4IN_52,ImgReg4IN_51,ImgReg4IN_50,
                      ImgReg4IN_49,ImgReg4IN_48})) ;
    triStateBuffer_16 loop3_3_TriState5N (.D ({DATA[63],DATA[62],DATA[61],
                      DATA[60],DATA[59],DATA[58],DATA[57],DATA[56],DATA[55],
                      DATA[54],DATA[53],DATA[52],DATA[51],DATA[50],DATA[49],
                      DATA[48]}), .EN (nx23594), .F ({ImgReg5IN_63,ImgReg5IN_62,
                      ImgReg5IN_61,ImgReg5IN_60,ImgReg5IN_59,ImgReg5IN_58,
                      ImgReg5IN_57,ImgReg5IN_56,ImgReg5IN_55,ImgReg5IN_54,
                      ImgReg5IN_53,ImgReg5IN_52,ImgReg5IN_51,ImgReg5IN_50,
                      ImgReg5IN_49,ImgReg5IN_48})) ;
    triStateBuffer_16 loop3_3_TriState0U (.D ({OutputImg1[63],OutputImg1[62],
                      OutputImg1[61],OutputImg1[60],OutputImg1[59],
                      OutputImg1[58],OutputImg1[57],OutputImg1[56],
                      OutputImg1[55],OutputImg1[54],OutputImg1[53],
                      OutputImg1[52],OutputImg1[51],OutputImg1[50],
                      OutputImg1[49],OutputImg1[48]}), .EN (nx23790), .F ({
                      ImgReg0IN_63,ImgReg0IN_62,ImgReg0IN_61,ImgReg0IN_60,
                      ImgReg0IN_59,ImgReg0IN_58,ImgReg0IN_57,ImgReg0IN_56,
                      ImgReg0IN_55,ImgReg0IN_54,ImgReg0IN_53,ImgReg0IN_52,
                      ImgReg0IN_51,ImgReg0IN_50,ImgReg0IN_49,ImgReg0IN_48})) ;
    triStateBuffer_16 loop3_3_TriState1U (.D ({OutputImg2[63],OutputImg2[62],
                      OutputImg2[61],OutputImg2[60],OutputImg2[59],
                      OutputImg2[58],OutputImg2[57],OutputImg2[56],
                      OutputImg2[55],OutputImg2[54],OutputImg2[53],
                      OutputImg2[52],OutputImg2[51],OutputImg2[50],
                      OutputImg2[49],OutputImg2[48]}), .EN (nx23790), .F ({
                      ImgReg1IN_63,ImgReg1IN_62,ImgReg1IN_61,ImgReg1IN_60,
                      ImgReg1IN_59,ImgReg1IN_58,ImgReg1IN_57,ImgReg1IN_56,
                      ImgReg1IN_55,ImgReg1IN_54,ImgReg1IN_53,ImgReg1IN_52,
                      ImgReg1IN_51,ImgReg1IN_50,ImgReg1IN_49,ImgReg1IN_48})) ;
    triStateBuffer_16 loop3_3_TriState2U (.D ({OutputImg3[63],OutputImg3[62],
                      OutputImg3[61],OutputImg3[60],OutputImg3[59],
                      OutputImg3[58],OutputImg3[57],OutputImg3[56],
                      OutputImg3[55],OutputImg3[54],OutputImg3[53],
                      OutputImg3[52],OutputImg3[51],OutputImg3[50],
                      OutputImg3[49],OutputImg3[48]}), .EN (nx23790), .F ({
                      ImgReg2IN_63,ImgReg2IN_62,ImgReg2IN_61,ImgReg2IN_60,
                      ImgReg2IN_59,ImgReg2IN_58,ImgReg2IN_57,ImgReg2IN_56,
                      ImgReg2IN_55,ImgReg2IN_54,ImgReg2IN_53,ImgReg2IN_52,
                      ImgReg2IN_51,ImgReg2IN_50,ImgReg2IN_49,ImgReg2IN_48})) ;
    triStateBuffer_16 loop3_3_TriState3U (.D ({OutputImg4[63],OutputImg4[62],
                      OutputImg4[61],OutputImg4[60],OutputImg4[59],
                      OutputImg4[58],OutputImg4[57],OutputImg4[56],
                      OutputImg4[55],OutputImg4[54],OutputImg4[53],
                      OutputImg4[52],OutputImg4[51],OutputImg4[50],
                      OutputImg4[49],OutputImg4[48]}), .EN (nx23790), .F ({
                      ImgReg3IN_63,ImgReg3IN_62,ImgReg3IN_61,ImgReg3IN_60,
                      ImgReg3IN_59,ImgReg3IN_58,ImgReg3IN_57,ImgReg3IN_56,
                      ImgReg3IN_55,ImgReg3IN_54,ImgReg3IN_53,ImgReg3IN_52,
                      ImgReg3IN_51,ImgReg3IN_50,ImgReg3IN_49,ImgReg3IN_48})) ;
    triStateBuffer_16 loop3_3_TriState4U (.D ({OutputImg5[63],OutputImg5[62],
                      OutputImg5[61],OutputImg5[60],OutputImg5[59],
                      OutputImg5[58],OutputImg5[57],OutputImg5[56],
                      OutputImg5[55],OutputImg5[54],OutputImg5[53],
                      OutputImg5[52],OutputImg5[51],OutputImg5[50],
                      OutputImg5[49],OutputImg5[48]}), .EN (nx23790), .F ({
                      ImgReg4IN_63,ImgReg4IN_62,ImgReg4IN_61,ImgReg4IN_60,
                      ImgReg4IN_59,ImgReg4IN_58,ImgReg4IN_57,ImgReg4IN_56,
                      ImgReg4IN_55,ImgReg4IN_54,ImgReg4IN_53,ImgReg4IN_52,
                      ImgReg4IN_51,ImgReg4IN_50,ImgReg4IN_49,ImgReg4IN_48})) ;
    nBitRegister_16 loop3_3_reg1 (.D ({ImgReg0IN_63,ImgReg0IN_62,ImgReg0IN_61,
                    ImgReg0IN_60,ImgReg0IN_59,ImgReg0IN_58,ImgReg0IN_57,
                    ImgReg0IN_56,ImgReg0IN_55,ImgReg0IN_54,ImgReg0IN_53,
                    ImgReg0IN_52,ImgReg0IN_51,ImgReg0IN_50,ImgReg0IN_49,
                    ImgReg0IN_48}), .CLK (nx23846), .RST (RST), .EN (nx23718), .Q (
                    {OutputImg0[63],OutputImg0[62],OutputImg0[61],OutputImg0[60]
                    ,OutputImg0[59],OutputImg0[58],OutputImg0[57],OutputImg0[56]
                    ,OutputImg0[55],OutputImg0[54],OutputImg0[53],OutputImg0[52]
                    ,OutputImg0[51],OutputImg0[50],OutputImg0[49],OutputImg0[48]
                    })) ;
    nBitRegister_16 loop3_3_reg2 (.D ({ImgReg1IN_63,ImgReg1IN_62,ImgReg1IN_61,
                    ImgReg1IN_60,ImgReg1IN_59,ImgReg1IN_58,ImgReg1IN_57,
                    ImgReg1IN_56,ImgReg1IN_55,ImgReg1IN_54,ImgReg1IN_53,
                    ImgReg1IN_52,ImgReg1IN_51,ImgReg1IN_50,ImgReg1IN_49,
                    ImgReg1IN_48}), .CLK (nx23848), .RST (RST), .EN (nx23728), .Q (
                    {OutputImg1[63],OutputImg1[62],OutputImg1[61],OutputImg1[60]
                    ,OutputImg1[59],OutputImg1[58],OutputImg1[57],OutputImg1[56]
                    ,OutputImg1[55],OutputImg1[54],OutputImg1[53],OutputImg1[52]
                    ,OutputImg1[51],OutputImg1[50],OutputImg1[49],OutputImg1[48]
                    })) ;
    nBitRegister_16 loop3_3_reg3 (.D ({ImgReg2IN_63,ImgReg2IN_62,ImgReg2IN_61,
                    ImgReg2IN_60,ImgReg2IN_59,ImgReg2IN_58,ImgReg2IN_57,
                    ImgReg2IN_56,ImgReg2IN_55,ImgReg2IN_54,ImgReg2IN_53,
                    ImgReg2IN_52,ImgReg2IN_51,ImgReg2IN_50,ImgReg2IN_49,
                    ImgReg2IN_48}), .CLK (nx23848), .RST (RST), .EN (nx23738), .Q (
                    {OutputImg2[63],OutputImg2[62],OutputImg2[61],OutputImg2[60]
                    ,OutputImg2[59],OutputImg2[58],OutputImg2[57],OutputImg2[56]
                    ,OutputImg2[55],OutputImg2[54],OutputImg2[53],OutputImg2[52]
                    ,OutputImg2[51],OutputImg2[50],OutputImg2[49],OutputImg2[48]
                    })) ;
    nBitRegister_16 loop3_3_reg4 (.D ({ImgReg3IN_63,ImgReg3IN_62,ImgReg3IN_61,
                    ImgReg3IN_60,ImgReg3IN_59,ImgReg3IN_58,ImgReg3IN_57,
                    ImgReg3IN_56,ImgReg3IN_55,ImgReg3IN_54,ImgReg3IN_53,
                    ImgReg3IN_52,ImgReg3IN_51,ImgReg3IN_50,ImgReg3IN_49,
                    ImgReg3IN_48}), .CLK (nx23850), .RST (RST), .EN (nx23748), .Q (
                    {OutputImg3[63],OutputImg3[62],OutputImg3[61],OutputImg3[60]
                    ,OutputImg3[59],OutputImg3[58],OutputImg3[57],OutputImg3[56]
                    ,OutputImg3[55],OutputImg3[54],OutputImg3[53],OutputImg3[52]
                    ,OutputImg3[51],OutputImg3[50],OutputImg3[49],OutputImg3[48]
                    })) ;
    nBitRegister_16 loop3_3_reg5 (.D ({ImgReg4IN_63,ImgReg4IN_62,ImgReg4IN_61,
                    ImgReg4IN_60,ImgReg4IN_59,ImgReg4IN_58,ImgReg4IN_57,
                    ImgReg4IN_56,ImgReg4IN_55,ImgReg4IN_54,ImgReg4IN_53,
                    ImgReg4IN_52,ImgReg4IN_51,ImgReg4IN_50,ImgReg4IN_49,
                    ImgReg4IN_48}), .CLK (nx23850), .RST (RST), .EN (nx23758), .Q (
                    {OutputImg4[63],OutputImg4[62],OutputImg4[61],OutputImg4[60]
                    ,OutputImg4[59],OutputImg4[58],OutputImg4[57],OutputImg4[56]
                    ,OutputImg4[55],OutputImg4[54],OutputImg4[53],OutputImg4[52]
                    ,OutputImg4[51],OutputImg4[50],OutputImg4[49],OutputImg4[48]
                    })) ;
    nBitRegister_16 loop3_3_reg6 (.D ({ImgReg5IN_63,ImgReg5IN_62,ImgReg5IN_61,
                    ImgReg5IN_60,ImgReg5IN_59,ImgReg5IN_58,ImgReg5IN_57,
                    ImgReg5IN_56,ImgReg5IN_55,ImgReg5IN_54,ImgReg5IN_53,
                    ImgReg5IN_52,ImgReg5IN_51,ImgReg5IN_50,ImgReg5IN_49,
                    ImgReg5IN_48}), .CLK (nx23852), .RST (RST), .EN (nx23768), .Q (
                    {OutputImg5[63],OutputImg5[62],OutputImg5[61],OutputImg5[60]
                    ,OutputImg5[59],OutputImg5[58],OutputImg5[57],OutputImg5[56]
                    ,OutputImg5[55],OutputImg5[54],OutputImg5[53],OutputImg5[52]
                    ,OutputImg5[51],OutputImg5[50],OutputImg5[49],OutputImg5[48]
                    })) ;
    triStateBuffer_16 loop3_4_TriState0L (.D ({OutputImg0[95],OutputImg0[94],
                      OutputImg0[93],OutputImg0[92],OutputImg0[91],
                      OutputImg0[90],OutputImg0[89],OutputImg0[88],
                      OutputImg0[87],OutputImg0[86],OutputImg0[85],
                      OutputImg0[84],OutputImg0[83],OutputImg0[82],
                      OutputImg0[81],OutputImg0[80]}), .EN (nx23672), .F ({
                      ImgReg0IN_79,ImgReg0IN_78,ImgReg0IN_77,ImgReg0IN_76,
                      ImgReg0IN_75,ImgReg0IN_74,ImgReg0IN_73,ImgReg0IN_72,
                      ImgReg0IN_71,ImgReg0IN_70,ImgReg0IN_69,ImgReg0IN_68,
                      ImgReg0IN_67,ImgReg0IN_66,ImgReg0IN_65,ImgReg0IN_64})) ;
    triStateBuffer_16 loop3_4_TriState1L (.D ({OutputImg1[95],OutputImg1[94],
                      OutputImg1[93],OutputImg1[92],OutputImg1[91],
                      OutputImg1[90],OutputImg1[89],OutputImg1[88],
                      OutputImg1[87],OutputImg1[86],OutputImg1[85],
                      OutputImg1[84],OutputImg1[83],OutputImg1[82],
                      OutputImg1[81],OutputImg1[80]}), .EN (nx23672), .F ({
                      ImgReg1IN_79,ImgReg1IN_78,ImgReg1IN_77,ImgReg1IN_76,
                      ImgReg1IN_75,ImgReg1IN_74,ImgReg1IN_73,ImgReg1IN_72,
                      ImgReg1IN_71,ImgReg1IN_70,ImgReg1IN_69,ImgReg1IN_68,
                      ImgReg1IN_67,ImgReg1IN_66,ImgReg1IN_65,ImgReg1IN_64})) ;
    triStateBuffer_16 loop3_4_TriState2L (.D ({OutputImg2[95],OutputImg2[94],
                      OutputImg2[93],OutputImg2[92],OutputImg2[91],
                      OutputImg2[90],OutputImg2[89],OutputImg2[88],
                      OutputImg2[87],OutputImg2[86],OutputImg2[85],
                      OutputImg2[84],OutputImg2[83],OutputImg2[82],
                      OutputImg2[81],OutputImg2[80]}), .EN (nx23672), .F ({
                      ImgReg2IN_79,ImgReg2IN_78,ImgReg2IN_77,ImgReg2IN_76,
                      ImgReg2IN_75,ImgReg2IN_74,ImgReg2IN_73,ImgReg2IN_72,
                      ImgReg2IN_71,ImgReg2IN_70,ImgReg2IN_69,ImgReg2IN_68,
                      ImgReg2IN_67,ImgReg2IN_66,ImgReg2IN_65,ImgReg2IN_64})) ;
    triStateBuffer_16 loop3_4_TriState3L (.D ({OutputImg3[95],OutputImg3[94],
                      OutputImg3[93],OutputImg3[92],OutputImg3[91],
                      OutputImg3[90],OutputImg3[89],OutputImg3[88],
                      OutputImg3[87],OutputImg3[86],OutputImg3[85],
                      OutputImg3[84],OutputImg3[83],OutputImg3[82],
                      OutputImg3[81],OutputImg3[80]}), .EN (nx23672), .F ({
                      ImgReg3IN_79,ImgReg3IN_78,ImgReg3IN_77,ImgReg3IN_76,
                      ImgReg3IN_75,ImgReg3IN_74,ImgReg3IN_73,ImgReg3IN_72,
                      ImgReg3IN_71,ImgReg3IN_70,ImgReg3IN_69,ImgReg3IN_68,
                      ImgReg3IN_67,ImgReg3IN_66,ImgReg3IN_65,ImgReg3IN_64})) ;
    triStateBuffer_16 loop3_4_TriState4L (.D ({OutputImg4[95],OutputImg4[94],
                      OutputImg4[93],OutputImg4[92],OutputImg4[91],
                      OutputImg4[90],OutputImg4[89],OutputImg4[88],
                      OutputImg4[87],OutputImg4[86],OutputImg4[85],
                      OutputImg4[84],OutputImg4[83],OutputImg4[82],
                      OutputImg4[81],OutputImg4[80]}), .EN (nx23674), .F ({
                      ImgReg4IN_79,ImgReg4IN_78,ImgReg4IN_77,ImgReg4IN_76,
                      ImgReg4IN_75,ImgReg4IN_74,ImgReg4IN_73,ImgReg4IN_72,
                      ImgReg4IN_71,ImgReg4IN_70,ImgReg4IN_69,ImgReg4IN_68,
                      ImgReg4IN_67,ImgReg4IN_66,ImgReg4IN_65,ImgReg4IN_64})) ;
    triStateBuffer_16 loop3_4_TriState5L (.D ({OutputImg5[95],OutputImg5[94],
                      OutputImg5[93],OutputImg5[92],OutputImg5[91],
                      OutputImg5[90],OutputImg5[89],OutputImg5[88],
                      OutputImg5[87],OutputImg5[86],OutputImg5[85],
                      OutputImg5[84],OutputImg5[83],OutputImg5[82],
                      OutputImg5[81],OutputImg5[80]}), .EN (nx23674), .F ({
                      ImgReg5IN_79,ImgReg5IN_78,ImgReg5IN_77,ImgReg5IN_76,
                      ImgReg5IN_75,ImgReg5IN_74,ImgReg5IN_73,ImgReg5IN_72,
                      ImgReg5IN_71,ImgReg5IN_70,ImgReg5IN_69,ImgReg5IN_68,
                      ImgReg5IN_67,ImgReg5IN_66,ImgReg5IN_65,ImgReg5IN_64})) ;
    triStateBuffer_16 loop3_4_TriState0N (.D ({DATA[79],DATA[78],DATA[77],
                      DATA[76],DATA[75],DATA[74],DATA[73],DATA[72],DATA[71],
                      DATA[70],DATA[69],DATA[68],DATA[67],DATA[66],DATA[65],
                      DATA[64]}), .EN (nx23654), .F ({ImgReg0IN_79,ImgReg0IN_78,
                      ImgReg0IN_77,ImgReg0IN_76,ImgReg0IN_75,ImgReg0IN_74,
                      ImgReg0IN_73,ImgReg0IN_72,ImgReg0IN_71,ImgReg0IN_70,
                      ImgReg0IN_69,ImgReg0IN_68,ImgReg0IN_67,ImgReg0IN_66,
                      ImgReg0IN_65,ImgReg0IN_64})) ;
    triStateBuffer_16 loop3_4_TriState1N (.D ({DATA[79],DATA[78],DATA[77],
                      DATA[76],DATA[75],DATA[74],DATA[73],DATA[72],DATA[71],
                      DATA[70],DATA[69],DATA[68],DATA[67],DATA[66],DATA[65],
                      DATA[64]}), .EN (nx23642), .F ({ImgReg1IN_79,ImgReg1IN_78,
                      ImgReg1IN_77,ImgReg1IN_76,ImgReg1IN_75,ImgReg1IN_74,
                      ImgReg1IN_73,ImgReg1IN_72,ImgReg1IN_71,ImgReg1IN_70,
                      ImgReg1IN_69,ImgReg1IN_68,ImgReg1IN_67,ImgReg1IN_66,
                      ImgReg1IN_65,ImgReg1IN_64})) ;
    triStateBuffer_16 loop3_4_TriState2N (.D ({DATA[79],DATA[78],DATA[77],
                      DATA[76],DATA[75],DATA[74],DATA[73],DATA[72],DATA[71],
                      DATA[70],DATA[69],DATA[68],DATA[67],DATA[66],DATA[65],
                      DATA[64]}), .EN (nx23630), .F ({ImgReg2IN_79,ImgReg2IN_78,
                      ImgReg2IN_77,ImgReg2IN_76,ImgReg2IN_75,ImgReg2IN_74,
                      ImgReg2IN_73,ImgReg2IN_72,ImgReg2IN_71,ImgReg2IN_70,
                      ImgReg2IN_69,ImgReg2IN_68,ImgReg2IN_67,ImgReg2IN_66,
                      ImgReg2IN_65,ImgReg2IN_64})) ;
    triStateBuffer_16 loop3_4_TriState3N (.D ({DATA[79],DATA[78],DATA[77],
                      DATA[76],DATA[75],DATA[74],DATA[73],DATA[72],DATA[71],
                      DATA[70],DATA[69],DATA[68],DATA[67],DATA[66],DATA[65],
                      DATA[64]}), .EN (nx23618), .F ({ImgReg3IN_79,ImgReg3IN_78,
                      ImgReg3IN_77,ImgReg3IN_76,ImgReg3IN_75,ImgReg3IN_74,
                      ImgReg3IN_73,ImgReg3IN_72,ImgReg3IN_71,ImgReg3IN_70,
                      ImgReg3IN_69,ImgReg3IN_68,ImgReg3IN_67,ImgReg3IN_66,
                      ImgReg3IN_65,ImgReg3IN_64})) ;
    triStateBuffer_16 loop3_4_TriState4N (.D ({DATA[79],DATA[78],DATA[77],
                      DATA[76],DATA[75],DATA[74],DATA[73],DATA[72],DATA[71],
                      DATA[70],DATA[69],DATA[68],DATA[67],DATA[66],DATA[65],
                      DATA[64]}), .EN (nx23606), .F ({ImgReg4IN_79,ImgReg4IN_78,
                      ImgReg4IN_77,ImgReg4IN_76,ImgReg4IN_75,ImgReg4IN_74,
                      ImgReg4IN_73,ImgReg4IN_72,ImgReg4IN_71,ImgReg4IN_70,
                      ImgReg4IN_69,ImgReg4IN_68,ImgReg4IN_67,ImgReg4IN_66,
                      ImgReg4IN_65,ImgReg4IN_64})) ;
    triStateBuffer_16 loop3_4_TriState5N (.D ({DATA[79],DATA[78],DATA[77],
                      DATA[76],DATA[75],DATA[74],DATA[73],DATA[72],DATA[71],
                      DATA[70],DATA[69],DATA[68],DATA[67],DATA[66],DATA[65],
                      DATA[64]}), .EN (nx23594), .F ({ImgReg5IN_79,ImgReg5IN_78,
                      ImgReg5IN_77,ImgReg5IN_76,ImgReg5IN_75,ImgReg5IN_74,
                      ImgReg5IN_73,ImgReg5IN_72,ImgReg5IN_71,ImgReg5IN_70,
                      ImgReg5IN_69,ImgReg5IN_68,ImgReg5IN_67,ImgReg5IN_66,
                      ImgReg5IN_65,ImgReg5IN_64})) ;
    triStateBuffer_16 loop3_4_TriState0U (.D ({OutputImg1[79],OutputImg1[78],
                      OutputImg1[77],OutputImg1[76],OutputImg1[75],
                      OutputImg1[74],OutputImg1[73],OutputImg1[72],
                      OutputImg1[71],OutputImg1[70],OutputImg1[69],
                      OutputImg1[68],OutputImg1[67],OutputImg1[66],
                      OutputImg1[65],OutputImg1[64]}), .EN (nx23790), .F ({
                      ImgReg0IN_79,ImgReg0IN_78,ImgReg0IN_77,ImgReg0IN_76,
                      ImgReg0IN_75,ImgReg0IN_74,ImgReg0IN_73,ImgReg0IN_72,
                      ImgReg0IN_71,ImgReg0IN_70,ImgReg0IN_69,ImgReg0IN_68,
                      ImgReg0IN_67,ImgReg0IN_66,ImgReg0IN_65,ImgReg0IN_64})) ;
    triStateBuffer_16 loop3_4_TriState1U (.D ({OutputImg2[79],OutputImg2[78],
                      OutputImg2[77],OutputImg2[76],OutputImg2[75],
                      OutputImg2[74],OutputImg2[73],OutputImg2[72],
                      OutputImg2[71],OutputImg2[70],OutputImg2[69],
                      OutputImg2[68],OutputImg2[67],OutputImg2[66],
                      OutputImg2[65],OutputImg2[64]}), .EN (nx23792), .F ({
                      ImgReg1IN_79,ImgReg1IN_78,ImgReg1IN_77,ImgReg1IN_76,
                      ImgReg1IN_75,ImgReg1IN_74,ImgReg1IN_73,ImgReg1IN_72,
                      ImgReg1IN_71,ImgReg1IN_70,ImgReg1IN_69,ImgReg1IN_68,
                      ImgReg1IN_67,ImgReg1IN_66,ImgReg1IN_65,ImgReg1IN_64})) ;
    triStateBuffer_16 loop3_4_TriState2U (.D ({OutputImg3[79],OutputImg3[78],
                      OutputImg3[77],OutputImg3[76],OutputImg3[75],
                      OutputImg3[74],OutputImg3[73],OutputImg3[72],
                      OutputImg3[71],OutputImg3[70],OutputImg3[69],
                      OutputImg3[68],OutputImg3[67],OutputImg3[66],
                      OutputImg3[65],OutputImg3[64]}), .EN (nx23792), .F ({
                      ImgReg2IN_79,ImgReg2IN_78,ImgReg2IN_77,ImgReg2IN_76,
                      ImgReg2IN_75,ImgReg2IN_74,ImgReg2IN_73,ImgReg2IN_72,
                      ImgReg2IN_71,ImgReg2IN_70,ImgReg2IN_69,ImgReg2IN_68,
                      ImgReg2IN_67,ImgReg2IN_66,ImgReg2IN_65,ImgReg2IN_64})) ;
    triStateBuffer_16 loop3_4_TriState3U (.D ({OutputImg4[79],OutputImg4[78],
                      OutputImg4[77],OutputImg4[76],OutputImg4[75],
                      OutputImg4[74],OutputImg4[73],OutputImg4[72],
                      OutputImg4[71],OutputImg4[70],OutputImg4[69],
                      OutputImg4[68],OutputImg4[67],OutputImg4[66],
                      OutputImg4[65],OutputImg4[64]}), .EN (nx23792), .F ({
                      ImgReg3IN_79,ImgReg3IN_78,ImgReg3IN_77,ImgReg3IN_76,
                      ImgReg3IN_75,ImgReg3IN_74,ImgReg3IN_73,ImgReg3IN_72,
                      ImgReg3IN_71,ImgReg3IN_70,ImgReg3IN_69,ImgReg3IN_68,
                      ImgReg3IN_67,ImgReg3IN_66,ImgReg3IN_65,ImgReg3IN_64})) ;
    triStateBuffer_16 loop3_4_TriState4U (.D ({OutputImg5[79],OutputImg5[78],
                      OutputImg5[77],OutputImg5[76],OutputImg5[75],
                      OutputImg5[74],OutputImg5[73],OutputImg5[72],
                      OutputImg5[71],OutputImg5[70],OutputImg5[69],
                      OutputImg5[68],OutputImg5[67],OutputImg5[66],
                      OutputImg5[65],OutputImg5[64]}), .EN (nx23792), .F ({
                      ImgReg4IN_79,ImgReg4IN_78,ImgReg4IN_77,ImgReg4IN_76,
                      ImgReg4IN_75,ImgReg4IN_74,ImgReg4IN_73,ImgReg4IN_72,
                      ImgReg4IN_71,ImgReg4IN_70,ImgReg4IN_69,ImgReg4IN_68,
                      ImgReg4IN_67,ImgReg4IN_66,ImgReg4IN_65,ImgReg4IN_64})) ;
    nBitRegister_16 loop3_4_reg1 (.D ({ImgReg0IN_79,ImgReg0IN_78,ImgReg0IN_77,
                    ImgReg0IN_76,ImgReg0IN_75,ImgReg0IN_74,ImgReg0IN_73,
                    ImgReg0IN_72,ImgReg0IN_71,ImgReg0IN_70,ImgReg0IN_69,
                    ImgReg0IN_68,ImgReg0IN_67,ImgReg0IN_66,ImgReg0IN_65,
                    ImgReg0IN_64}), .CLK (nx23852), .RST (RST), .EN (nx23718), .Q (
                    {OutputImg0[79],OutputImg0[78],OutputImg0[77],OutputImg0[76]
                    ,OutputImg0[75],OutputImg0[74],OutputImg0[73],OutputImg0[72]
                    ,OutputImg0[71],OutputImg0[70],OutputImg0[69],OutputImg0[68]
                    ,OutputImg0[67],OutputImg0[66],OutputImg0[65],OutputImg0[64]
                    })) ;
    nBitRegister_16 loop3_4_reg2 (.D ({ImgReg1IN_79,ImgReg1IN_78,ImgReg1IN_77,
                    ImgReg1IN_76,ImgReg1IN_75,ImgReg1IN_74,ImgReg1IN_73,
                    ImgReg1IN_72,ImgReg1IN_71,ImgReg1IN_70,ImgReg1IN_69,
                    ImgReg1IN_68,ImgReg1IN_67,ImgReg1IN_66,ImgReg1IN_65,
                    ImgReg1IN_64}), .CLK (nx23854), .RST (RST), .EN (nx23728), .Q (
                    {OutputImg1[79],OutputImg1[78],OutputImg1[77],OutputImg1[76]
                    ,OutputImg1[75],OutputImg1[74],OutputImg1[73],OutputImg1[72]
                    ,OutputImg1[71],OutputImg1[70],OutputImg1[69],OutputImg1[68]
                    ,OutputImg1[67],OutputImg1[66],OutputImg1[65],OutputImg1[64]
                    })) ;
    nBitRegister_16 loop3_4_reg3 (.D ({ImgReg2IN_79,ImgReg2IN_78,ImgReg2IN_77,
                    ImgReg2IN_76,ImgReg2IN_75,ImgReg2IN_74,ImgReg2IN_73,
                    ImgReg2IN_72,ImgReg2IN_71,ImgReg2IN_70,ImgReg2IN_69,
                    ImgReg2IN_68,ImgReg2IN_67,ImgReg2IN_66,ImgReg2IN_65,
                    ImgReg2IN_64}), .CLK (nx23854), .RST (RST), .EN (nx23738), .Q (
                    {OutputImg2[79],OutputImg2[78],OutputImg2[77],OutputImg2[76]
                    ,OutputImg2[75],OutputImg2[74],OutputImg2[73],OutputImg2[72]
                    ,OutputImg2[71],OutputImg2[70],OutputImg2[69],OutputImg2[68]
                    ,OutputImg2[67],OutputImg2[66],OutputImg2[65],OutputImg2[64]
                    })) ;
    nBitRegister_16 loop3_4_reg4 (.D ({ImgReg3IN_79,ImgReg3IN_78,ImgReg3IN_77,
                    ImgReg3IN_76,ImgReg3IN_75,ImgReg3IN_74,ImgReg3IN_73,
                    ImgReg3IN_72,ImgReg3IN_71,ImgReg3IN_70,ImgReg3IN_69,
                    ImgReg3IN_68,ImgReg3IN_67,ImgReg3IN_66,ImgReg3IN_65,
                    ImgReg3IN_64}), .CLK (nx23856), .RST (RST), .EN (nx23748), .Q (
                    {OutputImg3[79],OutputImg3[78],OutputImg3[77],OutputImg3[76]
                    ,OutputImg3[75],OutputImg3[74],OutputImg3[73],OutputImg3[72]
                    ,OutputImg3[71],OutputImg3[70],OutputImg3[69],OutputImg3[68]
                    ,OutputImg3[67],OutputImg3[66],OutputImg3[65],OutputImg3[64]
                    })) ;
    nBitRegister_16 loop3_4_reg5 (.D ({ImgReg4IN_79,ImgReg4IN_78,ImgReg4IN_77,
                    ImgReg4IN_76,ImgReg4IN_75,ImgReg4IN_74,ImgReg4IN_73,
                    ImgReg4IN_72,ImgReg4IN_71,ImgReg4IN_70,ImgReg4IN_69,
                    ImgReg4IN_68,ImgReg4IN_67,ImgReg4IN_66,ImgReg4IN_65,
                    ImgReg4IN_64}), .CLK (nx23856), .RST (RST), .EN (nx23758), .Q (
                    {OutputImg4[79],OutputImg4[78],OutputImg4[77],OutputImg4[76]
                    ,OutputImg4[75],OutputImg4[74],OutputImg4[73],OutputImg4[72]
                    ,OutputImg4[71],OutputImg4[70],OutputImg4[69],OutputImg4[68]
                    ,OutputImg4[67],OutputImg4[66],OutputImg4[65],OutputImg4[64]
                    })) ;
    nBitRegister_16 loop3_4_reg6 (.D ({ImgReg5IN_79,ImgReg5IN_78,ImgReg5IN_77,
                    ImgReg5IN_76,ImgReg5IN_75,ImgReg5IN_74,ImgReg5IN_73,
                    ImgReg5IN_72,ImgReg5IN_71,ImgReg5IN_70,ImgReg5IN_69,
                    ImgReg5IN_68,ImgReg5IN_67,ImgReg5IN_66,ImgReg5IN_65,
                    ImgReg5IN_64}), .CLK (nx23858), .RST (RST), .EN (nx23768), .Q (
                    {OutputImg5[79],OutputImg5[78],OutputImg5[77],OutputImg5[76]
                    ,OutputImg5[75],OutputImg5[74],OutputImg5[73],OutputImg5[72]
                    ,OutputImg5[71],OutputImg5[70],OutputImg5[69],OutputImg5[68]
                    ,OutputImg5[67],OutputImg5[66],OutputImg5[65],OutputImg5[64]
                    })) ;
    triStateBuffer_16 loop3_5_TriState0L (.D ({OutputImg0[111],OutputImg0[110],
                      OutputImg0[109],OutputImg0[108],OutputImg0[107],
                      OutputImg0[106],OutputImg0[105],OutputImg0[104],
                      OutputImg0[103],OutputImg0[102],OutputImg0[101],
                      OutputImg0[100],OutputImg0[99],OutputImg0[98],
                      OutputImg0[97],OutputImg0[96]}), .EN (nx23674), .F ({
                      ImgReg0IN_95,ImgReg0IN_94,ImgReg0IN_93,ImgReg0IN_92,
                      ImgReg0IN_91,ImgReg0IN_90,ImgReg0IN_89,ImgReg0IN_88,
                      ImgReg0IN_87,ImgReg0IN_86,ImgReg0IN_85,ImgReg0IN_84,
                      ImgReg0IN_83,ImgReg0IN_82,ImgReg0IN_81,ImgReg0IN_80})) ;
    triStateBuffer_16 loop3_5_TriState1L (.D ({OutputImg1[111],OutputImg1[110],
                      OutputImg1[109],OutputImg1[108],OutputImg1[107],
                      OutputImg1[106],OutputImg1[105],OutputImg1[104],
                      OutputImg1[103],OutputImg1[102],OutputImg1[101],
                      OutputImg1[100],OutputImg1[99],OutputImg1[98],
                      OutputImg1[97],OutputImg1[96]}), .EN (nx23674), .F ({
                      ImgReg1IN_95,ImgReg1IN_94,ImgReg1IN_93,ImgReg1IN_92,
                      ImgReg1IN_91,ImgReg1IN_90,ImgReg1IN_89,ImgReg1IN_88,
                      ImgReg1IN_87,ImgReg1IN_86,ImgReg1IN_85,ImgReg1IN_84,
                      ImgReg1IN_83,ImgReg1IN_82,ImgReg1IN_81,ImgReg1IN_80})) ;
    triStateBuffer_16 loop3_5_TriState2L (.D ({OutputImg2[111],OutputImg2[110],
                      OutputImg2[109],OutputImg2[108],OutputImg2[107],
                      OutputImg2[106],OutputImg2[105],OutputImg2[104],
                      OutputImg2[103],OutputImg2[102],OutputImg2[101],
                      OutputImg2[100],OutputImg2[99],OutputImg2[98],
                      OutputImg2[97],OutputImg2[96]}), .EN (nx23674), .F ({
                      ImgReg2IN_95,ImgReg2IN_94,ImgReg2IN_93,ImgReg2IN_92,
                      ImgReg2IN_91,ImgReg2IN_90,ImgReg2IN_89,ImgReg2IN_88,
                      ImgReg2IN_87,ImgReg2IN_86,ImgReg2IN_85,ImgReg2IN_84,
                      ImgReg2IN_83,ImgReg2IN_82,ImgReg2IN_81,ImgReg2IN_80})) ;
    triStateBuffer_16 loop3_5_TriState3L (.D ({OutputImg3[111],OutputImg3[110],
                      OutputImg3[109],OutputImg3[108],OutputImg3[107],
                      OutputImg3[106],OutputImg3[105],OutputImg3[104],
                      OutputImg3[103],OutputImg3[102],OutputImg3[101],
                      OutputImg3[100],OutputImg3[99],OutputImg3[98],
                      OutputImg3[97],OutputImg3[96]}), .EN (nx23674), .F ({
                      ImgReg3IN_95,ImgReg3IN_94,ImgReg3IN_93,ImgReg3IN_92,
                      ImgReg3IN_91,ImgReg3IN_90,ImgReg3IN_89,ImgReg3IN_88,
                      ImgReg3IN_87,ImgReg3IN_86,ImgReg3IN_85,ImgReg3IN_84,
                      ImgReg3IN_83,ImgReg3IN_82,ImgReg3IN_81,ImgReg3IN_80})) ;
    triStateBuffer_16 loop3_5_TriState4L (.D ({OutputImg4[111],OutputImg4[110],
                      OutputImg4[109],OutputImg4[108],OutputImg4[107],
                      OutputImg4[106],OutputImg4[105],OutputImg4[104],
                      OutputImg4[103],OutputImg4[102],OutputImg4[101],
                      OutputImg4[100],OutputImg4[99],OutputImg4[98],
                      OutputImg4[97],OutputImg4[96]}), .EN (nx23674), .F ({
                      ImgReg4IN_95,ImgReg4IN_94,ImgReg4IN_93,ImgReg4IN_92,
                      ImgReg4IN_91,ImgReg4IN_90,ImgReg4IN_89,ImgReg4IN_88,
                      ImgReg4IN_87,ImgReg4IN_86,ImgReg4IN_85,ImgReg4IN_84,
                      ImgReg4IN_83,ImgReg4IN_82,ImgReg4IN_81,ImgReg4IN_80})) ;
    triStateBuffer_16 loop3_5_TriState5L (.D ({OutputImg5[111],OutputImg5[110],
                      OutputImg5[109],OutputImg5[108],OutputImg5[107],
                      OutputImg5[106],OutputImg5[105],OutputImg5[104],
                      OutputImg5[103],OutputImg5[102],OutputImg5[101],
                      OutputImg5[100],OutputImg5[99],OutputImg5[98],
                      OutputImg5[97],OutputImg5[96]}), .EN (nx23676), .F ({
                      ImgReg5IN_95,ImgReg5IN_94,ImgReg5IN_93,ImgReg5IN_92,
                      ImgReg5IN_91,ImgReg5IN_90,ImgReg5IN_89,ImgReg5IN_88,
                      ImgReg5IN_87,ImgReg5IN_86,ImgReg5IN_85,ImgReg5IN_84,
                      ImgReg5IN_83,ImgReg5IN_82,ImgReg5IN_81,ImgReg5IN_80})) ;
    triStateBuffer_16 loop3_5_TriState0N (.D ({DATA[95],DATA[94],DATA[93],
                      DATA[92],DATA[91],DATA[90],DATA[89],DATA[88],DATA[87],
                      DATA[86],DATA[85],DATA[84],DATA[83],DATA[82],DATA[81],
                      DATA[80]}), .EN (nx23654), .F ({ImgReg0IN_95,ImgReg0IN_94,
                      ImgReg0IN_93,ImgReg0IN_92,ImgReg0IN_91,ImgReg0IN_90,
                      ImgReg0IN_89,ImgReg0IN_88,ImgReg0IN_87,ImgReg0IN_86,
                      ImgReg0IN_85,ImgReg0IN_84,ImgReg0IN_83,ImgReg0IN_82,
                      ImgReg0IN_81,ImgReg0IN_80})) ;
    triStateBuffer_16 loop3_5_TriState1N (.D ({DATA[95],DATA[94],DATA[93],
                      DATA[92],DATA[91],DATA[90],DATA[89],DATA[88],DATA[87],
                      DATA[86],DATA[85],DATA[84],DATA[83],DATA[82],DATA[81],
                      DATA[80]}), .EN (nx23642), .F ({ImgReg1IN_95,ImgReg1IN_94,
                      ImgReg1IN_93,ImgReg1IN_92,ImgReg1IN_91,ImgReg1IN_90,
                      ImgReg1IN_89,ImgReg1IN_88,ImgReg1IN_87,ImgReg1IN_86,
                      ImgReg1IN_85,ImgReg1IN_84,ImgReg1IN_83,ImgReg1IN_82,
                      ImgReg1IN_81,ImgReg1IN_80})) ;
    triStateBuffer_16 loop3_5_TriState2N (.D ({DATA[95],DATA[94],DATA[93],
                      DATA[92],DATA[91],DATA[90],DATA[89],DATA[88],DATA[87],
                      DATA[86],DATA[85],DATA[84],DATA[83],DATA[82],DATA[81],
                      DATA[80]}), .EN (nx23630), .F ({ImgReg2IN_95,ImgReg2IN_94,
                      ImgReg2IN_93,ImgReg2IN_92,ImgReg2IN_91,ImgReg2IN_90,
                      ImgReg2IN_89,ImgReg2IN_88,ImgReg2IN_87,ImgReg2IN_86,
                      ImgReg2IN_85,ImgReg2IN_84,ImgReg2IN_83,ImgReg2IN_82,
                      ImgReg2IN_81,ImgReg2IN_80})) ;
    triStateBuffer_16 loop3_5_TriState3N (.D ({DATA[95],DATA[94],DATA[93],
                      DATA[92],DATA[91],DATA[90],DATA[89],DATA[88],DATA[87],
                      DATA[86],DATA[85],DATA[84],DATA[83],DATA[82],DATA[81],
                      DATA[80]}), .EN (nx23618), .F ({ImgReg3IN_95,ImgReg3IN_94,
                      ImgReg3IN_93,ImgReg3IN_92,ImgReg3IN_91,ImgReg3IN_90,
                      ImgReg3IN_89,ImgReg3IN_88,ImgReg3IN_87,ImgReg3IN_86,
                      ImgReg3IN_85,ImgReg3IN_84,ImgReg3IN_83,ImgReg3IN_82,
                      ImgReg3IN_81,ImgReg3IN_80})) ;
    triStateBuffer_16 loop3_5_TriState4N (.D ({DATA[95],DATA[94],DATA[93],
                      DATA[92],DATA[91],DATA[90],DATA[89],DATA[88],DATA[87],
                      DATA[86],DATA[85],DATA[84],DATA[83],DATA[82],DATA[81],
                      DATA[80]}), .EN (nx23606), .F ({ImgReg4IN_95,ImgReg4IN_94,
                      ImgReg4IN_93,ImgReg4IN_92,ImgReg4IN_91,ImgReg4IN_90,
                      ImgReg4IN_89,ImgReg4IN_88,ImgReg4IN_87,ImgReg4IN_86,
                      ImgReg4IN_85,ImgReg4IN_84,ImgReg4IN_83,ImgReg4IN_82,
                      ImgReg4IN_81,ImgReg4IN_80})) ;
    triStateBuffer_16 loop3_5_TriState5N (.D ({DATA[95],DATA[94],DATA[93],
                      DATA[92],DATA[91],DATA[90],DATA[89],DATA[88],DATA[87],
                      DATA[86],DATA[85],DATA[84],DATA[83],DATA[82],DATA[81],
                      DATA[80]}), .EN (nx23594), .F ({ImgReg5IN_95,ImgReg5IN_94,
                      ImgReg5IN_93,ImgReg5IN_92,ImgReg5IN_91,ImgReg5IN_90,
                      ImgReg5IN_89,ImgReg5IN_88,ImgReg5IN_87,ImgReg5IN_86,
                      ImgReg5IN_85,ImgReg5IN_84,ImgReg5IN_83,ImgReg5IN_82,
                      ImgReg5IN_81,ImgReg5IN_80})) ;
    triStateBuffer_16 loop3_5_TriState0U (.D ({OutputImg1[95],OutputImg1[94],
                      OutputImg1[93],OutputImg1[92],OutputImg1[91],
                      OutputImg1[90],OutputImg1[89],OutputImg1[88],
                      OutputImg1[87],OutputImg1[86],OutputImg1[85],
                      OutputImg1[84],OutputImg1[83],OutputImg1[82],
                      OutputImg1[81],OutputImg1[80]}), .EN (nx23792), .F ({
                      ImgReg0IN_95,ImgReg0IN_94,ImgReg0IN_93,ImgReg0IN_92,
                      ImgReg0IN_91,ImgReg0IN_90,ImgReg0IN_89,ImgReg0IN_88,
                      ImgReg0IN_87,ImgReg0IN_86,ImgReg0IN_85,ImgReg0IN_84,
                      ImgReg0IN_83,ImgReg0IN_82,ImgReg0IN_81,ImgReg0IN_80})) ;
    triStateBuffer_16 loop3_5_TriState1U (.D ({OutputImg2[95],OutputImg2[94],
                      OutputImg2[93],OutputImg2[92],OutputImg2[91],
                      OutputImg2[90],OutputImg2[89],OutputImg2[88],
                      OutputImg2[87],OutputImg2[86],OutputImg2[85],
                      OutputImg2[84],OutputImg2[83],OutputImg2[82],
                      OutputImg2[81],OutputImg2[80]}), .EN (nx23792), .F ({
                      ImgReg1IN_95,ImgReg1IN_94,ImgReg1IN_93,ImgReg1IN_92,
                      ImgReg1IN_91,ImgReg1IN_90,ImgReg1IN_89,ImgReg1IN_88,
                      ImgReg1IN_87,ImgReg1IN_86,ImgReg1IN_85,ImgReg1IN_84,
                      ImgReg1IN_83,ImgReg1IN_82,ImgReg1IN_81,ImgReg1IN_80})) ;
    triStateBuffer_16 loop3_5_TriState2U (.D ({OutputImg3[95],OutputImg3[94],
                      OutputImg3[93],OutputImg3[92],OutputImg3[91],
                      OutputImg3[90],OutputImg3[89],OutputImg3[88],
                      OutputImg3[87],OutputImg3[86],OutputImg3[85],
                      OutputImg3[84],OutputImg3[83],OutputImg3[82],
                      OutputImg3[81],OutputImg3[80]}), .EN (nx23792), .F ({
                      ImgReg2IN_95,ImgReg2IN_94,ImgReg2IN_93,ImgReg2IN_92,
                      ImgReg2IN_91,ImgReg2IN_90,ImgReg2IN_89,ImgReg2IN_88,
                      ImgReg2IN_87,ImgReg2IN_86,ImgReg2IN_85,ImgReg2IN_84,
                      ImgReg2IN_83,ImgReg2IN_82,ImgReg2IN_81,ImgReg2IN_80})) ;
    triStateBuffer_16 loop3_5_TriState3U (.D ({OutputImg4[95],OutputImg4[94],
                      OutputImg4[93],OutputImg4[92],OutputImg4[91],
                      OutputImg4[90],OutputImg4[89],OutputImg4[88],
                      OutputImg4[87],OutputImg4[86],OutputImg4[85],
                      OutputImg4[84],OutputImg4[83],OutputImg4[82],
                      OutputImg4[81],OutputImg4[80]}), .EN (nx23794), .F ({
                      ImgReg3IN_95,ImgReg3IN_94,ImgReg3IN_93,ImgReg3IN_92,
                      ImgReg3IN_91,ImgReg3IN_90,ImgReg3IN_89,ImgReg3IN_88,
                      ImgReg3IN_87,ImgReg3IN_86,ImgReg3IN_85,ImgReg3IN_84,
                      ImgReg3IN_83,ImgReg3IN_82,ImgReg3IN_81,ImgReg3IN_80})) ;
    triStateBuffer_16 loop3_5_TriState4U (.D ({OutputImg5[95],OutputImg5[94],
                      OutputImg5[93],OutputImg5[92],OutputImg5[91],
                      OutputImg5[90],OutputImg5[89],OutputImg5[88],
                      OutputImg5[87],OutputImg5[86],OutputImg5[85],
                      OutputImg5[84],OutputImg5[83],OutputImg5[82],
                      OutputImg5[81],OutputImg5[80]}), .EN (nx23794), .F ({
                      ImgReg4IN_95,ImgReg4IN_94,ImgReg4IN_93,ImgReg4IN_92,
                      ImgReg4IN_91,ImgReg4IN_90,ImgReg4IN_89,ImgReg4IN_88,
                      ImgReg4IN_87,ImgReg4IN_86,ImgReg4IN_85,ImgReg4IN_84,
                      ImgReg4IN_83,ImgReg4IN_82,ImgReg4IN_81,ImgReg4IN_80})) ;
    nBitRegister_16 loop3_5_reg1 (.D ({ImgReg0IN_95,ImgReg0IN_94,ImgReg0IN_93,
                    ImgReg0IN_92,ImgReg0IN_91,ImgReg0IN_90,ImgReg0IN_89,
                    ImgReg0IN_88,ImgReg0IN_87,ImgReg0IN_86,ImgReg0IN_85,
                    ImgReg0IN_84,ImgReg0IN_83,ImgReg0IN_82,ImgReg0IN_81,
                    ImgReg0IN_80}), .CLK (nx23858), .RST (RST), .EN (nx23718), .Q (
                    {OutputImg0[95],OutputImg0[94],OutputImg0[93],OutputImg0[92]
                    ,OutputImg0[91],OutputImg0[90],OutputImg0[89],OutputImg0[88]
                    ,OutputImg0[87],OutputImg0[86],OutputImg0[85],OutputImg0[84]
                    ,OutputImg0[83],OutputImg0[82],OutputImg0[81],OutputImg0[80]
                    })) ;
    nBitRegister_16 loop3_5_reg2 (.D ({ImgReg1IN_95,ImgReg1IN_94,ImgReg1IN_93,
                    ImgReg1IN_92,ImgReg1IN_91,ImgReg1IN_90,ImgReg1IN_89,
                    ImgReg1IN_88,ImgReg1IN_87,ImgReg1IN_86,ImgReg1IN_85,
                    ImgReg1IN_84,ImgReg1IN_83,ImgReg1IN_82,ImgReg1IN_81,
                    ImgReg1IN_80}), .CLK (nx23860), .RST (RST), .EN (nx23728), .Q (
                    {OutputImg1[95],OutputImg1[94],OutputImg1[93],OutputImg1[92]
                    ,OutputImg1[91],OutputImg1[90],OutputImg1[89],OutputImg1[88]
                    ,OutputImg1[87],OutputImg1[86],OutputImg1[85],OutputImg1[84]
                    ,OutputImg1[83],OutputImg1[82],OutputImg1[81],OutputImg1[80]
                    })) ;
    nBitRegister_16 loop3_5_reg3 (.D ({ImgReg2IN_95,ImgReg2IN_94,ImgReg2IN_93,
                    ImgReg2IN_92,ImgReg2IN_91,ImgReg2IN_90,ImgReg2IN_89,
                    ImgReg2IN_88,ImgReg2IN_87,ImgReg2IN_86,ImgReg2IN_85,
                    ImgReg2IN_84,ImgReg2IN_83,ImgReg2IN_82,ImgReg2IN_81,
                    ImgReg2IN_80}), .CLK (nx23860), .RST (RST), .EN (nx23738), .Q (
                    {OutputImg2[95],OutputImg2[94],OutputImg2[93],OutputImg2[92]
                    ,OutputImg2[91],OutputImg2[90],OutputImg2[89],OutputImg2[88]
                    ,OutputImg2[87],OutputImg2[86],OutputImg2[85],OutputImg2[84]
                    ,OutputImg2[83],OutputImg2[82],OutputImg2[81],OutputImg2[80]
                    })) ;
    nBitRegister_16 loop3_5_reg4 (.D ({ImgReg3IN_95,ImgReg3IN_94,ImgReg3IN_93,
                    ImgReg3IN_92,ImgReg3IN_91,ImgReg3IN_90,ImgReg3IN_89,
                    ImgReg3IN_88,ImgReg3IN_87,ImgReg3IN_86,ImgReg3IN_85,
                    ImgReg3IN_84,ImgReg3IN_83,ImgReg3IN_82,ImgReg3IN_81,
                    ImgReg3IN_80}), .CLK (nx23862), .RST (RST), .EN (nx23748), .Q (
                    {OutputImg3[95],OutputImg3[94],OutputImg3[93],OutputImg3[92]
                    ,OutputImg3[91],OutputImg3[90],OutputImg3[89],OutputImg3[88]
                    ,OutputImg3[87],OutputImg3[86],OutputImg3[85],OutputImg3[84]
                    ,OutputImg3[83],OutputImg3[82],OutputImg3[81],OutputImg3[80]
                    })) ;
    nBitRegister_16 loop3_5_reg5 (.D ({ImgReg4IN_95,ImgReg4IN_94,ImgReg4IN_93,
                    ImgReg4IN_92,ImgReg4IN_91,ImgReg4IN_90,ImgReg4IN_89,
                    ImgReg4IN_88,ImgReg4IN_87,ImgReg4IN_86,ImgReg4IN_85,
                    ImgReg4IN_84,ImgReg4IN_83,ImgReg4IN_82,ImgReg4IN_81,
                    ImgReg4IN_80}), .CLK (nx23862), .RST (RST), .EN (nx23758), .Q (
                    {OutputImg4[95],OutputImg4[94],OutputImg4[93],OutputImg4[92]
                    ,OutputImg4[91],OutputImg4[90],OutputImg4[89],OutputImg4[88]
                    ,OutputImg4[87],OutputImg4[86],OutputImg4[85],OutputImg4[84]
                    ,OutputImg4[83],OutputImg4[82],OutputImg4[81],OutputImg4[80]
                    })) ;
    nBitRegister_16 loop3_5_reg6 (.D ({ImgReg5IN_95,ImgReg5IN_94,ImgReg5IN_93,
                    ImgReg5IN_92,ImgReg5IN_91,ImgReg5IN_90,ImgReg5IN_89,
                    ImgReg5IN_88,ImgReg5IN_87,ImgReg5IN_86,ImgReg5IN_85,
                    ImgReg5IN_84,ImgReg5IN_83,ImgReg5IN_82,ImgReg5IN_81,
                    ImgReg5IN_80}), .CLK (nx23864), .RST (RST), .EN (nx23768), .Q (
                    {OutputImg5[95],OutputImg5[94],OutputImg5[93],OutputImg5[92]
                    ,OutputImg5[91],OutputImg5[90],OutputImg5[89],OutputImg5[88]
                    ,OutputImg5[87],OutputImg5[86],OutputImg5[85],OutputImg5[84]
                    ,OutputImg5[83],OutputImg5[82],OutputImg5[81],OutputImg5[80]
                    })) ;
    triStateBuffer_16 loop3_6_TriState0L (.D ({OutputImg0[127],OutputImg0[126],
                      OutputImg0[125],OutputImg0[124],OutputImg0[123],
                      OutputImg0[122],OutputImg0[121],OutputImg0[120],
                      OutputImg0[119],OutputImg0[118],OutputImg0[117],
                      OutputImg0[116],OutputImg0[115],OutputImg0[114],
                      OutputImg0[113],OutputImg0[112]}), .EN (nx23676), .F ({
                      ImgReg0IN_111,ImgReg0IN_110,ImgReg0IN_109,ImgReg0IN_108,
                      ImgReg0IN_107,ImgReg0IN_106,ImgReg0IN_105,ImgReg0IN_104,
                      ImgReg0IN_103,ImgReg0IN_102,ImgReg0IN_101,ImgReg0IN_100,
                      ImgReg0IN_99,ImgReg0IN_98,ImgReg0IN_97,ImgReg0IN_96})) ;
    triStateBuffer_16 loop3_6_TriState1L (.D ({OutputImg1[127],OutputImg1[126],
                      OutputImg1[125],OutputImg1[124],OutputImg1[123],
                      OutputImg1[122],OutputImg1[121],OutputImg1[120],
                      OutputImg1[119],OutputImg1[118],OutputImg1[117],
                      OutputImg1[116],OutputImg1[115],OutputImg1[114],
                      OutputImg1[113],OutputImg1[112]}), .EN (nx23676), .F ({
                      ImgReg1IN_111,ImgReg1IN_110,ImgReg1IN_109,ImgReg1IN_108,
                      ImgReg1IN_107,ImgReg1IN_106,ImgReg1IN_105,ImgReg1IN_104,
                      ImgReg1IN_103,ImgReg1IN_102,ImgReg1IN_101,ImgReg1IN_100,
                      ImgReg1IN_99,ImgReg1IN_98,ImgReg1IN_97,ImgReg1IN_96})) ;
    triStateBuffer_16 loop3_6_TriState2L (.D ({OutputImg2[127],OutputImg2[126],
                      OutputImg2[125],OutputImg2[124],OutputImg2[123],
                      OutputImg2[122],OutputImg2[121],OutputImg2[120],
                      OutputImg2[119],OutputImg2[118],OutputImg2[117],
                      OutputImg2[116],OutputImg2[115],OutputImg2[114],
                      OutputImg2[113],OutputImg2[112]}), .EN (nx23676), .F ({
                      ImgReg2IN_111,ImgReg2IN_110,ImgReg2IN_109,ImgReg2IN_108,
                      ImgReg2IN_107,ImgReg2IN_106,ImgReg2IN_105,ImgReg2IN_104,
                      ImgReg2IN_103,ImgReg2IN_102,ImgReg2IN_101,ImgReg2IN_100,
                      ImgReg2IN_99,ImgReg2IN_98,ImgReg2IN_97,ImgReg2IN_96})) ;
    triStateBuffer_16 loop3_6_TriState3L (.D ({OutputImg3[127],OutputImg3[126],
                      OutputImg3[125],OutputImg3[124],OutputImg3[123],
                      OutputImg3[122],OutputImg3[121],OutputImg3[120],
                      OutputImg3[119],OutputImg3[118],OutputImg3[117],
                      OutputImg3[116],OutputImg3[115],OutputImg3[114],
                      OutputImg3[113],OutputImg3[112]}), .EN (nx23676), .F ({
                      ImgReg3IN_111,ImgReg3IN_110,ImgReg3IN_109,ImgReg3IN_108,
                      ImgReg3IN_107,ImgReg3IN_106,ImgReg3IN_105,ImgReg3IN_104,
                      ImgReg3IN_103,ImgReg3IN_102,ImgReg3IN_101,ImgReg3IN_100,
                      ImgReg3IN_99,ImgReg3IN_98,ImgReg3IN_97,ImgReg3IN_96})) ;
    triStateBuffer_16 loop3_6_TriState4L (.D ({OutputImg4[127],OutputImg4[126],
                      OutputImg4[125],OutputImg4[124],OutputImg4[123],
                      OutputImg4[122],OutputImg4[121],OutputImg4[120],
                      OutputImg4[119],OutputImg4[118],OutputImg4[117],
                      OutputImg4[116],OutputImg4[115],OutputImg4[114],
                      OutputImg4[113],OutputImg4[112]}), .EN (nx23676), .F ({
                      ImgReg4IN_111,ImgReg4IN_110,ImgReg4IN_109,ImgReg4IN_108,
                      ImgReg4IN_107,ImgReg4IN_106,ImgReg4IN_105,ImgReg4IN_104,
                      ImgReg4IN_103,ImgReg4IN_102,ImgReg4IN_101,ImgReg4IN_100,
                      ImgReg4IN_99,ImgReg4IN_98,ImgReg4IN_97,ImgReg4IN_96})) ;
    triStateBuffer_16 loop3_6_TriState5L (.D ({OutputImg5[127],OutputImg5[126],
                      OutputImg5[125],OutputImg5[124],OutputImg5[123],
                      OutputImg5[122],OutputImg5[121],OutputImg5[120],
                      OutputImg5[119],OutputImg5[118],OutputImg5[117],
                      OutputImg5[116],OutputImg5[115],OutputImg5[114],
                      OutputImg5[113],OutputImg5[112]}), .EN (nx23676), .F ({
                      ImgReg5IN_111,ImgReg5IN_110,ImgReg5IN_109,ImgReg5IN_108,
                      ImgReg5IN_107,ImgReg5IN_106,ImgReg5IN_105,ImgReg5IN_104,
                      ImgReg5IN_103,ImgReg5IN_102,ImgReg5IN_101,ImgReg5IN_100,
                      ImgReg5IN_99,ImgReg5IN_98,ImgReg5IN_97,ImgReg5IN_96})) ;
    triStateBuffer_16 loop3_6_TriState0N (.D ({DATA[111],DATA[110],DATA[109],
                      DATA[108],DATA[107],DATA[106],DATA[105],DATA[104],
                      DATA[103],DATA[102],DATA[101],DATA[100],DATA[99],DATA[98],
                      DATA[97],DATA[96]}), .EN (nx23654), .F ({ImgReg0IN_111,
                      ImgReg0IN_110,ImgReg0IN_109,ImgReg0IN_108,ImgReg0IN_107,
                      ImgReg0IN_106,ImgReg0IN_105,ImgReg0IN_104,ImgReg0IN_103,
                      ImgReg0IN_102,ImgReg0IN_101,ImgReg0IN_100,ImgReg0IN_99,
                      ImgReg0IN_98,ImgReg0IN_97,ImgReg0IN_96})) ;
    triStateBuffer_16 loop3_6_TriState1N (.D ({DATA[111],DATA[110],DATA[109],
                      DATA[108],DATA[107],DATA[106],DATA[105],DATA[104],
                      DATA[103],DATA[102],DATA[101],DATA[100],DATA[99],DATA[98],
                      DATA[97],DATA[96]}), .EN (nx23642), .F ({ImgReg1IN_111,
                      ImgReg1IN_110,ImgReg1IN_109,ImgReg1IN_108,ImgReg1IN_107,
                      ImgReg1IN_106,ImgReg1IN_105,ImgReg1IN_104,ImgReg1IN_103,
                      ImgReg1IN_102,ImgReg1IN_101,ImgReg1IN_100,ImgReg1IN_99,
                      ImgReg1IN_98,ImgReg1IN_97,ImgReg1IN_96})) ;
    triStateBuffer_16 loop3_6_TriState2N (.D ({DATA[111],DATA[110],DATA[109],
                      DATA[108],DATA[107],DATA[106],DATA[105],DATA[104],
                      DATA[103],DATA[102],DATA[101],DATA[100],DATA[99],DATA[98],
                      DATA[97],DATA[96]}), .EN (nx23630), .F ({ImgReg2IN_111,
                      ImgReg2IN_110,ImgReg2IN_109,ImgReg2IN_108,ImgReg2IN_107,
                      ImgReg2IN_106,ImgReg2IN_105,ImgReg2IN_104,ImgReg2IN_103,
                      ImgReg2IN_102,ImgReg2IN_101,ImgReg2IN_100,ImgReg2IN_99,
                      ImgReg2IN_98,ImgReg2IN_97,ImgReg2IN_96})) ;
    triStateBuffer_16 loop3_6_TriState3N (.D ({DATA[111],DATA[110],DATA[109],
                      DATA[108],DATA[107],DATA[106],DATA[105],DATA[104],
                      DATA[103],DATA[102],DATA[101],DATA[100],DATA[99],DATA[98],
                      DATA[97],DATA[96]}), .EN (nx23618), .F ({ImgReg3IN_111,
                      ImgReg3IN_110,ImgReg3IN_109,ImgReg3IN_108,ImgReg3IN_107,
                      ImgReg3IN_106,ImgReg3IN_105,ImgReg3IN_104,ImgReg3IN_103,
                      ImgReg3IN_102,ImgReg3IN_101,ImgReg3IN_100,ImgReg3IN_99,
                      ImgReg3IN_98,ImgReg3IN_97,ImgReg3IN_96})) ;
    triStateBuffer_16 loop3_6_TriState4N (.D ({DATA[111],DATA[110],DATA[109],
                      DATA[108],DATA[107],DATA[106],DATA[105],DATA[104],
                      DATA[103],DATA[102],DATA[101],DATA[100],DATA[99],DATA[98],
                      DATA[97],DATA[96]}), .EN (nx23606), .F ({ImgReg4IN_111,
                      ImgReg4IN_110,ImgReg4IN_109,ImgReg4IN_108,ImgReg4IN_107,
                      ImgReg4IN_106,ImgReg4IN_105,ImgReg4IN_104,ImgReg4IN_103,
                      ImgReg4IN_102,ImgReg4IN_101,ImgReg4IN_100,ImgReg4IN_99,
                      ImgReg4IN_98,ImgReg4IN_97,ImgReg4IN_96})) ;
    triStateBuffer_16 loop3_6_TriState5N (.D ({DATA[111],DATA[110],DATA[109],
                      DATA[108],DATA[107],DATA[106],DATA[105],DATA[104],
                      DATA[103],DATA[102],DATA[101],DATA[100],DATA[99],DATA[98],
                      DATA[97],DATA[96]}), .EN (nx23594), .F ({ImgReg5IN_111,
                      ImgReg5IN_110,ImgReg5IN_109,ImgReg5IN_108,ImgReg5IN_107,
                      ImgReg5IN_106,ImgReg5IN_105,ImgReg5IN_104,ImgReg5IN_103,
                      ImgReg5IN_102,ImgReg5IN_101,ImgReg5IN_100,ImgReg5IN_99,
                      ImgReg5IN_98,ImgReg5IN_97,ImgReg5IN_96})) ;
    triStateBuffer_16 loop3_6_TriState0U (.D ({OutputImg1[111],OutputImg1[110],
                      OutputImg1[109],OutputImg1[108],OutputImg1[107],
                      OutputImg1[106],OutputImg1[105],OutputImg1[104],
                      OutputImg1[103],OutputImg1[102],OutputImg1[101],
                      OutputImg1[100],OutputImg1[99],OutputImg1[98],
                      OutputImg1[97],OutputImg1[96]}), .EN (nx23794), .F ({
                      ImgReg0IN_111,ImgReg0IN_110,ImgReg0IN_109,ImgReg0IN_108,
                      ImgReg0IN_107,ImgReg0IN_106,ImgReg0IN_105,ImgReg0IN_104,
                      ImgReg0IN_103,ImgReg0IN_102,ImgReg0IN_101,ImgReg0IN_100,
                      ImgReg0IN_99,ImgReg0IN_98,ImgReg0IN_97,ImgReg0IN_96})) ;
    triStateBuffer_16 loop3_6_TriState1U (.D ({OutputImg2[111],OutputImg2[110],
                      OutputImg2[109],OutputImg2[108],OutputImg2[107],
                      OutputImg2[106],OutputImg2[105],OutputImg2[104],
                      OutputImg2[103],OutputImg2[102],OutputImg2[101],
                      OutputImg2[100],OutputImg2[99],OutputImg2[98],
                      OutputImg2[97],OutputImg2[96]}), .EN (nx23794), .F ({
                      ImgReg1IN_111,ImgReg1IN_110,ImgReg1IN_109,ImgReg1IN_108,
                      ImgReg1IN_107,ImgReg1IN_106,ImgReg1IN_105,ImgReg1IN_104,
                      ImgReg1IN_103,ImgReg1IN_102,ImgReg1IN_101,ImgReg1IN_100,
                      ImgReg1IN_99,ImgReg1IN_98,ImgReg1IN_97,ImgReg1IN_96})) ;
    triStateBuffer_16 loop3_6_TriState2U (.D ({OutputImg3[111],OutputImg3[110],
                      OutputImg3[109],OutputImg3[108],OutputImg3[107],
                      OutputImg3[106],OutputImg3[105],OutputImg3[104],
                      OutputImg3[103],OutputImg3[102],OutputImg3[101],
                      OutputImg3[100],OutputImg3[99],OutputImg3[98],
                      OutputImg3[97],OutputImg3[96]}), .EN (nx23794), .F ({
                      ImgReg2IN_111,ImgReg2IN_110,ImgReg2IN_109,ImgReg2IN_108,
                      ImgReg2IN_107,ImgReg2IN_106,ImgReg2IN_105,ImgReg2IN_104,
                      ImgReg2IN_103,ImgReg2IN_102,ImgReg2IN_101,ImgReg2IN_100,
                      ImgReg2IN_99,ImgReg2IN_98,ImgReg2IN_97,ImgReg2IN_96})) ;
    triStateBuffer_16 loop3_6_TriState3U (.D ({OutputImg4[111],OutputImg4[110],
                      OutputImg4[109],OutputImg4[108],OutputImg4[107],
                      OutputImg4[106],OutputImg4[105],OutputImg4[104],
                      OutputImg4[103],OutputImg4[102],OutputImg4[101],
                      OutputImg4[100],OutputImg4[99],OutputImg4[98],
                      OutputImg4[97],OutputImg4[96]}), .EN (nx23794), .F ({
                      ImgReg3IN_111,ImgReg3IN_110,ImgReg3IN_109,ImgReg3IN_108,
                      ImgReg3IN_107,ImgReg3IN_106,ImgReg3IN_105,ImgReg3IN_104,
                      ImgReg3IN_103,ImgReg3IN_102,ImgReg3IN_101,ImgReg3IN_100,
                      ImgReg3IN_99,ImgReg3IN_98,ImgReg3IN_97,ImgReg3IN_96})) ;
    triStateBuffer_16 loop3_6_TriState4U (.D ({OutputImg5[111],OutputImg5[110],
                      OutputImg5[109],OutputImg5[108],OutputImg5[107],
                      OutputImg5[106],OutputImg5[105],OutputImg5[104],
                      OutputImg5[103],OutputImg5[102],OutputImg5[101],
                      OutputImg5[100],OutputImg5[99],OutputImg5[98],
                      OutputImg5[97],OutputImg5[96]}), .EN (nx23794), .F ({
                      ImgReg4IN_111,ImgReg4IN_110,ImgReg4IN_109,ImgReg4IN_108,
                      ImgReg4IN_107,ImgReg4IN_106,ImgReg4IN_105,ImgReg4IN_104,
                      ImgReg4IN_103,ImgReg4IN_102,ImgReg4IN_101,ImgReg4IN_100,
                      ImgReg4IN_99,ImgReg4IN_98,ImgReg4IN_97,ImgReg4IN_96})) ;
    nBitRegister_16 loop3_6_reg1 (.D ({ImgReg0IN_111,ImgReg0IN_110,ImgReg0IN_109
                    ,ImgReg0IN_108,ImgReg0IN_107,ImgReg0IN_106,ImgReg0IN_105,
                    ImgReg0IN_104,ImgReg0IN_103,ImgReg0IN_102,ImgReg0IN_101,
                    ImgReg0IN_100,ImgReg0IN_99,ImgReg0IN_98,ImgReg0IN_97,
                    ImgReg0IN_96}), .CLK (nx23864), .RST (RST), .EN (nx23718), .Q (
                    {OutputImg0[111],OutputImg0[110],OutputImg0[109],
                    OutputImg0[108],OutputImg0[107],OutputImg0[106],
                    OutputImg0[105],OutputImg0[104],OutputImg0[103],
                    OutputImg0[102],OutputImg0[101],OutputImg0[100],
                    OutputImg0[99],OutputImg0[98],OutputImg0[97],OutputImg0[96]}
                    )) ;
    nBitRegister_16 loop3_6_reg2 (.D ({ImgReg1IN_111,ImgReg1IN_110,ImgReg1IN_109
                    ,ImgReg1IN_108,ImgReg1IN_107,ImgReg1IN_106,ImgReg1IN_105,
                    ImgReg1IN_104,ImgReg1IN_103,ImgReg1IN_102,ImgReg1IN_101,
                    ImgReg1IN_100,ImgReg1IN_99,ImgReg1IN_98,ImgReg1IN_97,
                    ImgReg1IN_96}), .CLK (nx23866), .RST (RST), .EN (nx23728), .Q (
                    {OutputImg1[111],OutputImg1[110],OutputImg1[109],
                    OutputImg1[108],OutputImg1[107],OutputImg1[106],
                    OutputImg1[105],OutputImg1[104],OutputImg1[103],
                    OutputImg1[102],OutputImg1[101],OutputImg1[100],
                    OutputImg1[99],OutputImg1[98],OutputImg1[97],OutputImg1[96]}
                    )) ;
    nBitRegister_16 loop3_6_reg3 (.D ({ImgReg2IN_111,ImgReg2IN_110,ImgReg2IN_109
                    ,ImgReg2IN_108,ImgReg2IN_107,ImgReg2IN_106,ImgReg2IN_105,
                    ImgReg2IN_104,ImgReg2IN_103,ImgReg2IN_102,ImgReg2IN_101,
                    ImgReg2IN_100,ImgReg2IN_99,ImgReg2IN_98,ImgReg2IN_97,
                    ImgReg2IN_96}), .CLK (nx23866), .RST (RST), .EN (nx23738), .Q (
                    {OutputImg2[111],OutputImg2[110],OutputImg2[109],
                    OutputImg2[108],OutputImg2[107],OutputImg2[106],
                    OutputImg2[105],OutputImg2[104],OutputImg2[103],
                    OutputImg2[102],OutputImg2[101],OutputImg2[100],
                    OutputImg2[99],OutputImg2[98],OutputImg2[97],OutputImg2[96]}
                    )) ;
    nBitRegister_16 loop3_6_reg4 (.D ({ImgReg3IN_111,ImgReg3IN_110,ImgReg3IN_109
                    ,ImgReg3IN_108,ImgReg3IN_107,ImgReg3IN_106,ImgReg3IN_105,
                    ImgReg3IN_104,ImgReg3IN_103,ImgReg3IN_102,ImgReg3IN_101,
                    ImgReg3IN_100,ImgReg3IN_99,ImgReg3IN_98,ImgReg3IN_97,
                    ImgReg3IN_96}), .CLK (nx23868), .RST (RST), .EN (nx23748), .Q (
                    {OutputImg3[111],OutputImg3[110],OutputImg3[109],
                    OutputImg3[108],OutputImg3[107],OutputImg3[106],
                    OutputImg3[105],OutputImg3[104],OutputImg3[103],
                    OutputImg3[102],OutputImg3[101],OutputImg3[100],
                    OutputImg3[99],OutputImg3[98],OutputImg3[97],OutputImg3[96]}
                    )) ;
    nBitRegister_16 loop3_6_reg5 (.D ({ImgReg4IN_111,ImgReg4IN_110,ImgReg4IN_109
                    ,ImgReg4IN_108,ImgReg4IN_107,ImgReg4IN_106,ImgReg4IN_105,
                    ImgReg4IN_104,ImgReg4IN_103,ImgReg4IN_102,ImgReg4IN_101,
                    ImgReg4IN_100,ImgReg4IN_99,ImgReg4IN_98,ImgReg4IN_97,
                    ImgReg4IN_96}), .CLK (nx23868), .RST (RST), .EN (nx23758), .Q (
                    {OutputImg4[111],OutputImg4[110],OutputImg4[109],
                    OutputImg4[108],OutputImg4[107],OutputImg4[106],
                    OutputImg4[105],OutputImg4[104],OutputImg4[103],
                    OutputImg4[102],OutputImg4[101],OutputImg4[100],
                    OutputImg4[99],OutputImg4[98],OutputImg4[97],OutputImg4[96]}
                    )) ;
    nBitRegister_16 loop3_6_reg6 (.D ({ImgReg5IN_111,ImgReg5IN_110,ImgReg5IN_109
                    ,ImgReg5IN_108,ImgReg5IN_107,ImgReg5IN_106,ImgReg5IN_105,
                    ImgReg5IN_104,ImgReg5IN_103,ImgReg5IN_102,ImgReg5IN_101,
                    ImgReg5IN_100,ImgReg5IN_99,ImgReg5IN_98,ImgReg5IN_97,
                    ImgReg5IN_96}), .CLK (nx23870), .RST (RST), .EN (nx23768), .Q (
                    {OutputImg5[111],OutputImg5[110],OutputImg5[109],
                    OutputImg5[108],OutputImg5[107],OutputImg5[106],
                    OutputImg5[105],OutputImg5[104],OutputImg5[103],
                    OutputImg5[102],OutputImg5[101],OutputImg5[100],
                    OutputImg5[99],OutputImg5[98],OutputImg5[97],OutputImg5[96]}
                    )) ;
    triStateBuffer_16 loop3_7_TriState0L (.D ({OutputImg0[143],OutputImg0[142],
                      OutputImg0[141],OutputImg0[140],OutputImg0[139],
                      OutputImg0[138],OutputImg0[137],OutputImg0[136],
                      OutputImg0[135],OutputImg0[134],OutputImg0[133],
                      OutputImg0[132],OutputImg0[131],OutputImg0[130],
                      OutputImg0[129],OutputImg0[128]}), .EN (nx23678), .F ({
                      ImgReg0IN_127,ImgReg0IN_126,ImgReg0IN_125,ImgReg0IN_124,
                      ImgReg0IN_123,ImgReg0IN_122,ImgReg0IN_121,ImgReg0IN_120,
                      ImgReg0IN_119,ImgReg0IN_118,ImgReg0IN_117,ImgReg0IN_116,
                      ImgReg0IN_115,ImgReg0IN_114,ImgReg0IN_113,ImgReg0IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState1L (.D ({OutputImg1[143],OutputImg1[142],
                      OutputImg1[141],OutputImg1[140],OutputImg1[139],
                      OutputImg1[138],OutputImg1[137],OutputImg1[136],
                      OutputImg1[135],OutputImg1[134],OutputImg1[133],
                      OutputImg1[132],OutputImg1[131],OutputImg1[130],
                      OutputImg1[129],OutputImg1[128]}), .EN (nx23678), .F ({
                      ImgReg1IN_127,ImgReg1IN_126,ImgReg1IN_125,ImgReg1IN_124,
                      ImgReg1IN_123,ImgReg1IN_122,ImgReg1IN_121,ImgReg1IN_120,
                      ImgReg1IN_119,ImgReg1IN_118,ImgReg1IN_117,ImgReg1IN_116,
                      ImgReg1IN_115,ImgReg1IN_114,ImgReg1IN_113,ImgReg1IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState2L (.D ({OutputImg2[143],OutputImg2[142],
                      OutputImg2[141],OutputImg2[140],OutputImg2[139],
                      OutputImg2[138],OutputImg2[137],OutputImg2[136],
                      OutputImg2[135],OutputImg2[134],OutputImg2[133],
                      OutputImg2[132],OutputImg2[131],OutputImg2[130],
                      OutputImg2[129],OutputImg2[128]}), .EN (nx23678), .F ({
                      ImgReg2IN_127,ImgReg2IN_126,ImgReg2IN_125,ImgReg2IN_124,
                      ImgReg2IN_123,ImgReg2IN_122,ImgReg2IN_121,ImgReg2IN_120,
                      ImgReg2IN_119,ImgReg2IN_118,ImgReg2IN_117,ImgReg2IN_116,
                      ImgReg2IN_115,ImgReg2IN_114,ImgReg2IN_113,ImgReg2IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState3L (.D ({OutputImg3[143],OutputImg3[142],
                      OutputImg3[141],OutputImg3[140],OutputImg3[139],
                      OutputImg3[138],OutputImg3[137],OutputImg3[136],
                      OutputImg3[135],OutputImg3[134],OutputImg3[133],
                      OutputImg3[132],OutputImg3[131],OutputImg3[130],
                      OutputImg3[129],OutputImg3[128]}), .EN (nx23678), .F ({
                      ImgReg3IN_127,ImgReg3IN_126,ImgReg3IN_125,ImgReg3IN_124,
                      ImgReg3IN_123,ImgReg3IN_122,ImgReg3IN_121,ImgReg3IN_120,
                      ImgReg3IN_119,ImgReg3IN_118,ImgReg3IN_117,ImgReg3IN_116,
                      ImgReg3IN_115,ImgReg3IN_114,ImgReg3IN_113,ImgReg3IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState4L (.D ({OutputImg4[143],OutputImg4[142],
                      OutputImg4[141],OutputImg4[140],OutputImg4[139],
                      OutputImg4[138],OutputImg4[137],OutputImg4[136],
                      OutputImg4[135],OutputImg4[134],OutputImg4[133],
                      OutputImg4[132],OutputImg4[131],OutputImg4[130],
                      OutputImg4[129],OutputImg4[128]}), .EN (nx23678), .F ({
                      ImgReg4IN_127,ImgReg4IN_126,ImgReg4IN_125,ImgReg4IN_124,
                      ImgReg4IN_123,ImgReg4IN_122,ImgReg4IN_121,ImgReg4IN_120,
                      ImgReg4IN_119,ImgReg4IN_118,ImgReg4IN_117,ImgReg4IN_116,
                      ImgReg4IN_115,ImgReg4IN_114,ImgReg4IN_113,ImgReg4IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState5L (.D ({OutputImg5[143],OutputImg5[142],
                      OutputImg5[141],OutputImg5[140],OutputImg5[139],
                      OutputImg5[138],OutputImg5[137],OutputImg5[136],
                      OutputImg5[135],OutputImg5[134],OutputImg5[133],
                      OutputImg5[132],OutputImg5[131],OutputImg5[130],
                      OutputImg5[129],OutputImg5[128]}), .EN (nx23678), .F ({
                      ImgReg5IN_127,ImgReg5IN_126,ImgReg5IN_125,ImgReg5IN_124,
                      ImgReg5IN_123,ImgReg5IN_122,ImgReg5IN_121,ImgReg5IN_120,
                      ImgReg5IN_119,ImgReg5IN_118,ImgReg5IN_117,ImgReg5IN_116,
                      ImgReg5IN_115,ImgReg5IN_114,ImgReg5IN_113,ImgReg5IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState0N (.D ({DATA[127],DATA[126],DATA[125],
                      DATA[124],DATA[123],DATA[122],DATA[121],DATA[120],
                      DATA[119],DATA[118],DATA[117],DATA[116],DATA[115],
                      DATA[114],DATA[113],DATA[112]}), .EN (nx23656), .F ({
                      ImgReg0IN_127,ImgReg0IN_126,ImgReg0IN_125,ImgReg0IN_124,
                      ImgReg0IN_123,ImgReg0IN_122,ImgReg0IN_121,ImgReg0IN_120,
                      ImgReg0IN_119,ImgReg0IN_118,ImgReg0IN_117,ImgReg0IN_116,
                      ImgReg0IN_115,ImgReg0IN_114,ImgReg0IN_113,ImgReg0IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState1N (.D ({DATA[127],DATA[126],DATA[125],
                      DATA[124],DATA[123],DATA[122],DATA[121],DATA[120],
                      DATA[119],DATA[118],DATA[117],DATA[116],DATA[115],
                      DATA[114],DATA[113],DATA[112]}), .EN (nx23644), .F ({
                      ImgReg1IN_127,ImgReg1IN_126,ImgReg1IN_125,ImgReg1IN_124,
                      ImgReg1IN_123,ImgReg1IN_122,ImgReg1IN_121,ImgReg1IN_120,
                      ImgReg1IN_119,ImgReg1IN_118,ImgReg1IN_117,ImgReg1IN_116,
                      ImgReg1IN_115,ImgReg1IN_114,ImgReg1IN_113,ImgReg1IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState2N (.D ({DATA[127],DATA[126],DATA[125],
                      DATA[124],DATA[123],DATA[122],DATA[121],DATA[120],
                      DATA[119],DATA[118],DATA[117],DATA[116],DATA[115],
                      DATA[114],DATA[113],DATA[112]}), .EN (nx23632), .F ({
                      ImgReg2IN_127,ImgReg2IN_126,ImgReg2IN_125,ImgReg2IN_124,
                      ImgReg2IN_123,ImgReg2IN_122,ImgReg2IN_121,ImgReg2IN_120,
                      ImgReg2IN_119,ImgReg2IN_118,ImgReg2IN_117,ImgReg2IN_116,
                      ImgReg2IN_115,ImgReg2IN_114,ImgReg2IN_113,ImgReg2IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState3N (.D ({DATA[127],DATA[126],DATA[125],
                      DATA[124],DATA[123],DATA[122],DATA[121],DATA[120],
                      DATA[119],DATA[118],DATA[117],DATA[116],DATA[115],
                      DATA[114],DATA[113],DATA[112]}), .EN (nx23620), .F ({
                      ImgReg3IN_127,ImgReg3IN_126,ImgReg3IN_125,ImgReg3IN_124,
                      ImgReg3IN_123,ImgReg3IN_122,ImgReg3IN_121,ImgReg3IN_120,
                      ImgReg3IN_119,ImgReg3IN_118,ImgReg3IN_117,ImgReg3IN_116,
                      ImgReg3IN_115,ImgReg3IN_114,ImgReg3IN_113,ImgReg3IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState4N (.D ({DATA[127],DATA[126],DATA[125],
                      DATA[124],DATA[123],DATA[122],DATA[121],DATA[120],
                      DATA[119],DATA[118],DATA[117],DATA[116],DATA[115],
                      DATA[114],DATA[113],DATA[112]}), .EN (nx23608), .F ({
                      ImgReg4IN_127,ImgReg4IN_126,ImgReg4IN_125,ImgReg4IN_124,
                      ImgReg4IN_123,ImgReg4IN_122,ImgReg4IN_121,ImgReg4IN_120,
                      ImgReg4IN_119,ImgReg4IN_118,ImgReg4IN_117,ImgReg4IN_116,
                      ImgReg4IN_115,ImgReg4IN_114,ImgReg4IN_113,ImgReg4IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState5N (.D ({DATA[127],DATA[126],DATA[125],
                      DATA[124],DATA[123],DATA[122],DATA[121],DATA[120],
                      DATA[119],DATA[118],DATA[117],DATA[116],DATA[115],
                      DATA[114],DATA[113],DATA[112]}), .EN (nx23596), .F ({
                      ImgReg5IN_127,ImgReg5IN_126,ImgReg5IN_125,ImgReg5IN_124,
                      ImgReg5IN_123,ImgReg5IN_122,ImgReg5IN_121,ImgReg5IN_120,
                      ImgReg5IN_119,ImgReg5IN_118,ImgReg5IN_117,ImgReg5IN_116,
                      ImgReg5IN_115,ImgReg5IN_114,ImgReg5IN_113,ImgReg5IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState0U (.D ({OutputImg1[127],OutputImg1[126],
                      OutputImg1[125],OutputImg1[124],OutputImg1[123],
                      OutputImg1[122],OutputImg1[121],OutputImg1[120],
                      OutputImg1[119],OutputImg1[118],OutputImg1[117],
                      OutputImg1[116],OutputImg1[115],OutputImg1[114],
                      OutputImg1[113],OutputImg1[112]}), .EN (nx23796), .F ({
                      ImgReg0IN_127,ImgReg0IN_126,ImgReg0IN_125,ImgReg0IN_124,
                      ImgReg0IN_123,ImgReg0IN_122,ImgReg0IN_121,ImgReg0IN_120,
                      ImgReg0IN_119,ImgReg0IN_118,ImgReg0IN_117,ImgReg0IN_116,
                      ImgReg0IN_115,ImgReg0IN_114,ImgReg0IN_113,ImgReg0IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState1U (.D ({OutputImg2[127],OutputImg2[126],
                      OutputImg2[125],OutputImg2[124],OutputImg2[123],
                      OutputImg2[122],OutputImg2[121],OutputImg2[120],
                      OutputImg2[119],OutputImg2[118],OutputImg2[117],
                      OutputImg2[116],OutputImg2[115],OutputImg2[114],
                      OutputImg2[113],OutputImg2[112]}), .EN (nx23796), .F ({
                      ImgReg1IN_127,ImgReg1IN_126,ImgReg1IN_125,ImgReg1IN_124,
                      ImgReg1IN_123,ImgReg1IN_122,ImgReg1IN_121,ImgReg1IN_120,
                      ImgReg1IN_119,ImgReg1IN_118,ImgReg1IN_117,ImgReg1IN_116,
                      ImgReg1IN_115,ImgReg1IN_114,ImgReg1IN_113,ImgReg1IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState2U (.D ({OutputImg3[127],OutputImg3[126],
                      OutputImg3[125],OutputImg3[124],OutputImg3[123],
                      OutputImg3[122],OutputImg3[121],OutputImg3[120],
                      OutputImg3[119],OutputImg3[118],OutputImg3[117],
                      OutputImg3[116],OutputImg3[115],OutputImg3[114],
                      OutputImg3[113],OutputImg3[112]}), .EN (nx23796), .F ({
                      ImgReg2IN_127,ImgReg2IN_126,ImgReg2IN_125,ImgReg2IN_124,
                      ImgReg2IN_123,ImgReg2IN_122,ImgReg2IN_121,ImgReg2IN_120,
                      ImgReg2IN_119,ImgReg2IN_118,ImgReg2IN_117,ImgReg2IN_116,
                      ImgReg2IN_115,ImgReg2IN_114,ImgReg2IN_113,ImgReg2IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState3U (.D ({OutputImg4[127],OutputImg4[126],
                      OutputImg4[125],OutputImg4[124],OutputImg4[123],
                      OutputImg4[122],OutputImg4[121],OutputImg4[120],
                      OutputImg4[119],OutputImg4[118],OutputImg4[117],
                      OutputImg4[116],OutputImg4[115],OutputImg4[114],
                      OutputImg4[113],OutputImg4[112]}), .EN (nx23796), .F ({
                      ImgReg3IN_127,ImgReg3IN_126,ImgReg3IN_125,ImgReg3IN_124,
                      ImgReg3IN_123,ImgReg3IN_122,ImgReg3IN_121,ImgReg3IN_120,
                      ImgReg3IN_119,ImgReg3IN_118,ImgReg3IN_117,ImgReg3IN_116,
                      ImgReg3IN_115,ImgReg3IN_114,ImgReg3IN_113,ImgReg3IN_112})
                      ) ;
    triStateBuffer_16 loop3_7_TriState4U (.D ({OutputImg5[127],OutputImg5[126],
                      OutputImg5[125],OutputImg5[124],OutputImg5[123],
                      OutputImg5[122],OutputImg5[121],OutputImg5[120],
                      OutputImg5[119],OutputImg5[118],OutputImg5[117],
                      OutputImg5[116],OutputImg5[115],OutputImg5[114],
                      OutputImg5[113],OutputImg5[112]}), .EN (nx23796), .F ({
                      ImgReg4IN_127,ImgReg4IN_126,ImgReg4IN_125,ImgReg4IN_124,
                      ImgReg4IN_123,ImgReg4IN_122,ImgReg4IN_121,ImgReg4IN_120,
                      ImgReg4IN_119,ImgReg4IN_118,ImgReg4IN_117,ImgReg4IN_116,
                      ImgReg4IN_115,ImgReg4IN_114,ImgReg4IN_113,ImgReg4IN_112})
                      ) ;
    nBitRegister_16 loop3_7_reg1 (.D ({ImgReg0IN_127,ImgReg0IN_126,ImgReg0IN_125
                    ,ImgReg0IN_124,ImgReg0IN_123,ImgReg0IN_122,ImgReg0IN_121,
                    ImgReg0IN_120,ImgReg0IN_119,ImgReg0IN_118,ImgReg0IN_117,
                    ImgReg0IN_116,ImgReg0IN_115,ImgReg0IN_114,ImgReg0IN_113,
                    ImgReg0IN_112}), .CLK (nx23870), .RST (RST), .EN (nx23720), 
                    .Q ({OutputImg0[127],OutputImg0[126],OutputImg0[125],
                    OutputImg0[124],OutputImg0[123],OutputImg0[122],
                    OutputImg0[121],OutputImg0[120],OutputImg0[119],
                    OutputImg0[118],OutputImg0[117],OutputImg0[116],
                    OutputImg0[115],OutputImg0[114],OutputImg0[113],
                    OutputImg0[112]})) ;
    nBitRegister_16 loop3_7_reg2 (.D ({ImgReg1IN_127,ImgReg1IN_126,ImgReg1IN_125
                    ,ImgReg1IN_124,ImgReg1IN_123,ImgReg1IN_122,ImgReg1IN_121,
                    ImgReg1IN_120,ImgReg1IN_119,ImgReg1IN_118,ImgReg1IN_117,
                    ImgReg1IN_116,ImgReg1IN_115,ImgReg1IN_114,ImgReg1IN_113,
                    ImgReg1IN_112}), .CLK (nx23872), .RST (RST), .EN (nx23730), 
                    .Q ({OutputImg1[127],OutputImg1[126],OutputImg1[125],
                    OutputImg1[124],OutputImg1[123],OutputImg1[122],
                    OutputImg1[121],OutputImg1[120],OutputImg1[119],
                    OutputImg1[118],OutputImg1[117],OutputImg1[116],
                    OutputImg1[115],OutputImg1[114],OutputImg1[113],
                    OutputImg1[112]})) ;
    nBitRegister_16 loop3_7_reg3 (.D ({ImgReg2IN_127,ImgReg2IN_126,ImgReg2IN_125
                    ,ImgReg2IN_124,ImgReg2IN_123,ImgReg2IN_122,ImgReg2IN_121,
                    ImgReg2IN_120,ImgReg2IN_119,ImgReg2IN_118,ImgReg2IN_117,
                    ImgReg2IN_116,ImgReg2IN_115,ImgReg2IN_114,ImgReg2IN_113,
                    ImgReg2IN_112}), .CLK (nx23872), .RST (RST), .EN (nx23740), 
                    .Q ({OutputImg2[127],OutputImg2[126],OutputImg2[125],
                    OutputImg2[124],OutputImg2[123],OutputImg2[122],
                    OutputImg2[121],OutputImg2[120],OutputImg2[119],
                    OutputImg2[118],OutputImg2[117],OutputImg2[116],
                    OutputImg2[115],OutputImg2[114],OutputImg2[113],
                    OutputImg2[112]})) ;
    nBitRegister_16 loop3_7_reg4 (.D ({ImgReg3IN_127,ImgReg3IN_126,ImgReg3IN_125
                    ,ImgReg3IN_124,ImgReg3IN_123,ImgReg3IN_122,ImgReg3IN_121,
                    ImgReg3IN_120,ImgReg3IN_119,ImgReg3IN_118,ImgReg3IN_117,
                    ImgReg3IN_116,ImgReg3IN_115,ImgReg3IN_114,ImgReg3IN_113,
                    ImgReg3IN_112}), .CLK (nx23874), .RST (RST), .EN (nx23750), 
                    .Q ({OutputImg3[127],OutputImg3[126],OutputImg3[125],
                    OutputImg3[124],OutputImg3[123],OutputImg3[122],
                    OutputImg3[121],OutputImg3[120],OutputImg3[119],
                    OutputImg3[118],OutputImg3[117],OutputImg3[116],
                    OutputImg3[115],OutputImg3[114],OutputImg3[113],
                    OutputImg3[112]})) ;
    nBitRegister_16 loop3_7_reg5 (.D ({ImgReg4IN_127,ImgReg4IN_126,ImgReg4IN_125
                    ,ImgReg4IN_124,ImgReg4IN_123,ImgReg4IN_122,ImgReg4IN_121,
                    ImgReg4IN_120,ImgReg4IN_119,ImgReg4IN_118,ImgReg4IN_117,
                    ImgReg4IN_116,ImgReg4IN_115,ImgReg4IN_114,ImgReg4IN_113,
                    ImgReg4IN_112}), .CLK (nx23874), .RST (RST), .EN (nx23760), 
                    .Q ({OutputImg4[127],OutputImg4[126],OutputImg4[125],
                    OutputImg4[124],OutputImg4[123],OutputImg4[122],
                    OutputImg4[121],OutputImg4[120],OutputImg4[119],
                    OutputImg4[118],OutputImg4[117],OutputImg4[116],
                    OutputImg4[115],OutputImg4[114],OutputImg4[113],
                    OutputImg4[112]})) ;
    nBitRegister_16 loop3_7_reg6 (.D ({ImgReg5IN_127,ImgReg5IN_126,ImgReg5IN_125
                    ,ImgReg5IN_124,ImgReg5IN_123,ImgReg5IN_122,ImgReg5IN_121,
                    ImgReg5IN_120,ImgReg5IN_119,ImgReg5IN_118,ImgReg5IN_117,
                    ImgReg5IN_116,ImgReg5IN_115,ImgReg5IN_114,ImgReg5IN_113,
                    ImgReg5IN_112}), .CLK (nx23876), .RST (RST), .EN (nx23770), 
                    .Q ({OutputImg5[127],OutputImg5[126],OutputImg5[125],
                    OutputImg5[124],OutputImg5[123],OutputImg5[122],
                    OutputImg5[121],OutputImg5[120],OutputImg5[119],
                    OutputImg5[118],OutputImg5[117],OutputImg5[116],
                    OutputImg5[115],OutputImg5[114],OutputImg5[113],
                    OutputImg5[112]})) ;
    triStateBuffer_16 loop3_8_TriState0L (.D ({OutputImg0[159],OutputImg0[158],
                      OutputImg0[157],OutputImg0[156],OutputImg0[155],
                      OutputImg0[154],OutputImg0[153],OutputImg0[152],
                      OutputImg0[151],OutputImg0[150],OutputImg0[149],
                      OutputImg0[148],OutputImg0[147],OutputImg0[146],
                      OutputImg0[145],OutputImg0[144]}), .EN (nx23678), .F ({
                      ImgReg0IN_143,ImgReg0IN_142,ImgReg0IN_141,ImgReg0IN_140,
                      ImgReg0IN_139,ImgReg0IN_138,ImgReg0IN_137,ImgReg0IN_136,
                      ImgReg0IN_135,ImgReg0IN_134,ImgReg0IN_133,ImgReg0IN_132,
                      ImgReg0IN_131,ImgReg0IN_130,ImgReg0IN_129,ImgReg0IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState1L (.D ({OutputImg1[159],OutputImg1[158],
                      OutputImg1[157],OutputImg1[156],OutputImg1[155],
                      OutputImg1[154],OutputImg1[153],OutputImg1[152],
                      OutputImg1[151],OutputImg1[150],OutputImg1[149],
                      OutputImg1[148],OutputImg1[147],OutputImg1[146],
                      OutputImg1[145],OutputImg1[144]}), .EN (nx23680), .F ({
                      ImgReg1IN_143,ImgReg1IN_142,ImgReg1IN_141,ImgReg1IN_140,
                      ImgReg1IN_139,ImgReg1IN_138,ImgReg1IN_137,ImgReg1IN_136,
                      ImgReg1IN_135,ImgReg1IN_134,ImgReg1IN_133,ImgReg1IN_132,
                      ImgReg1IN_131,ImgReg1IN_130,ImgReg1IN_129,ImgReg1IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState2L (.D ({OutputImg2[159],OutputImg2[158],
                      OutputImg2[157],OutputImg2[156],OutputImg2[155],
                      OutputImg2[154],OutputImg2[153],OutputImg2[152],
                      OutputImg2[151],OutputImg2[150],OutputImg2[149],
                      OutputImg2[148],OutputImg2[147],OutputImg2[146],
                      OutputImg2[145],OutputImg2[144]}), .EN (nx23680), .F ({
                      ImgReg2IN_143,ImgReg2IN_142,ImgReg2IN_141,ImgReg2IN_140,
                      ImgReg2IN_139,ImgReg2IN_138,ImgReg2IN_137,ImgReg2IN_136,
                      ImgReg2IN_135,ImgReg2IN_134,ImgReg2IN_133,ImgReg2IN_132,
                      ImgReg2IN_131,ImgReg2IN_130,ImgReg2IN_129,ImgReg2IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState3L (.D ({OutputImg3[159],OutputImg3[158],
                      OutputImg3[157],OutputImg3[156],OutputImg3[155],
                      OutputImg3[154],OutputImg3[153],OutputImg3[152],
                      OutputImg3[151],OutputImg3[150],OutputImg3[149],
                      OutputImg3[148],OutputImg3[147],OutputImg3[146],
                      OutputImg3[145],OutputImg3[144]}), .EN (nx23680), .F ({
                      ImgReg3IN_143,ImgReg3IN_142,ImgReg3IN_141,ImgReg3IN_140,
                      ImgReg3IN_139,ImgReg3IN_138,ImgReg3IN_137,ImgReg3IN_136,
                      ImgReg3IN_135,ImgReg3IN_134,ImgReg3IN_133,ImgReg3IN_132,
                      ImgReg3IN_131,ImgReg3IN_130,ImgReg3IN_129,ImgReg3IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState4L (.D ({OutputImg4[159],OutputImg4[158],
                      OutputImg4[157],OutputImg4[156],OutputImg4[155],
                      OutputImg4[154],OutputImg4[153],OutputImg4[152],
                      OutputImg4[151],OutputImg4[150],OutputImg4[149],
                      OutputImg4[148],OutputImg4[147],OutputImg4[146],
                      OutputImg4[145],OutputImg4[144]}), .EN (nx23680), .F ({
                      ImgReg4IN_143,ImgReg4IN_142,ImgReg4IN_141,ImgReg4IN_140,
                      ImgReg4IN_139,ImgReg4IN_138,ImgReg4IN_137,ImgReg4IN_136,
                      ImgReg4IN_135,ImgReg4IN_134,ImgReg4IN_133,ImgReg4IN_132,
                      ImgReg4IN_131,ImgReg4IN_130,ImgReg4IN_129,ImgReg4IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState5L (.D ({OutputImg5[159],OutputImg5[158],
                      OutputImg5[157],OutputImg5[156],OutputImg5[155],
                      OutputImg5[154],OutputImg5[153],OutputImg5[152],
                      OutputImg5[151],OutputImg5[150],OutputImg5[149],
                      OutputImg5[148],OutputImg5[147],OutputImg5[146],
                      OutputImg5[145],OutputImg5[144]}), .EN (nx23680), .F ({
                      ImgReg5IN_143,ImgReg5IN_142,ImgReg5IN_141,ImgReg5IN_140,
                      ImgReg5IN_139,ImgReg5IN_138,ImgReg5IN_137,ImgReg5IN_136,
                      ImgReg5IN_135,ImgReg5IN_134,ImgReg5IN_133,ImgReg5IN_132,
                      ImgReg5IN_131,ImgReg5IN_130,ImgReg5IN_129,ImgReg5IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState0N (.D ({DATA[143],DATA[142],DATA[141],
                      DATA[140],DATA[139],DATA[138],DATA[137],DATA[136],
                      DATA[135],DATA[134],DATA[133],DATA[132],DATA[131],
                      DATA[130],DATA[129],DATA[128]}), .EN (nx23656), .F ({
                      ImgReg0IN_143,ImgReg0IN_142,ImgReg0IN_141,ImgReg0IN_140,
                      ImgReg0IN_139,ImgReg0IN_138,ImgReg0IN_137,ImgReg0IN_136,
                      ImgReg0IN_135,ImgReg0IN_134,ImgReg0IN_133,ImgReg0IN_132,
                      ImgReg0IN_131,ImgReg0IN_130,ImgReg0IN_129,ImgReg0IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState1N (.D ({DATA[143],DATA[142],DATA[141],
                      DATA[140],DATA[139],DATA[138],DATA[137],DATA[136],
                      DATA[135],DATA[134],DATA[133],DATA[132],DATA[131],
                      DATA[130],DATA[129],DATA[128]}), .EN (nx23644), .F ({
                      ImgReg1IN_143,ImgReg1IN_142,ImgReg1IN_141,ImgReg1IN_140,
                      ImgReg1IN_139,ImgReg1IN_138,ImgReg1IN_137,ImgReg1IN_136,
                      ImgReg1IN_135,ImgReg1IN_134,ImgReg1IN_133,ImgReg1IN_132,
                      ImgReg1IN_131,ImgReg1IN_130,ImgReg1IN_129,ImgReg1IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState2N (.D ({DATA[143],DATA[142],DATA[141],
                      DATA[140],DATA[139],DATA[138],DATA[137],DATA[136],
                      DATA[135],DATA[134],DATA[133],DATA[132],DATA[131],
                      DATA[130],DATA[129],DATA[128]}), .EN (nx23632), .F ({
                      ImgReg2IN_143,ImgReg2IN_142,ImgReg2IN_141,ImgReg2IN_140,
                      ImgReg2IN_139,ImgReg2IN_138,ImgReg2IN_137,ImgReg2IN_136,
                      ImgReg2IN_135,ImgReg2IN_134,ImgReg2IN_133,ImgReg2IN_132,
                      ImgReg2IN_131,ImgReg2IN_130,ImgReg2IN_129,ImgReg2IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState3N (.D ({DATA[143],DATA[142],DATA[141],
                      DATA[140],DATA[139],DATA[138],DATA[137],DATA[136],
                      DATA[135],DATA[134],DATA[133],DATA[132],DATA[131],
                      DATA[130],DATA[129],DATA[128]}), .EN (nx23620), .F ({
                      ImgReg3IN_143,ImgReg3IN_142,ImgReg3IN_141,ImgReg3IN_140,
                      ImgReg3IN_139,ImgReg3IN_138,ImgReg3IN_137,ImgReg3IN_136,
                      ImgReg3IN_135,ImgReg3IN_134,ImgReg3IN_133,ImgReg3IN_132,
                      ImgReg3IN_131,ImgReg3IN_130,ImgReg3IN_129,ImgReg3IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState4N (.D ({DATA[143],DATA[142],DATA[141],
                      DATA[140],DATA[139],DATA[138],DATA[137],DATA[136],
                      DATA[135],DATA[134],DATA[133],DATA[132],DATA[131],
                      DATA[130],DATA[129],DATA[128]}), .EN (nx23608), .F ({
                      ImgReg4IN_143,ImgReg4IN_142,ImgReg4IN_141,ImgReg4IN_140,
                      ImgReg4IN_139,ImgReg4IN_138,ImgReg4IN_137,ImgReg4IN_136,
                      ImgReg4IN_135,ImgReg4IN_134,ImgReg4IN_133,ImgReg4IN_132,
                      ImgReg4IN_131,ImgReg4IN_130,ImgReg4IN_129,ImgReg4IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState5N (.D ({DATA[143],DATA[142],DATA[141],
                      DATA[140],DATA[139],DATA[138],DATA[137],DATA[136],
                      DATA[135],DATA[134],DATA[133],DATA[132],DATA[131],
                      DATA[130],DATA[129],DATA[128]}), .EN (nx23596), .F ({
                      ImgReg5IN_143,ImgReg5IN_142,ImgReg5IN_141,ImgReg5IN_140,
                      ImgReg5IN_139,ImgReg5IN_138,ImgReg5IN_137,ImgReg5IN_136,
                      ImgReg5IN_135,ImgReg5IN_134,ImgReg5IN_133,ImgReg5IN_132,
                      ImgReg5IN_131,ImgReg5IN_130,ImgReg5IN_129,ImgReg5IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState0U (.D ({OutputImg1[143],OutputImg1[142],
                      OutputImg1[141],OutputImg1[140],OutputImg1[139],
                      OutputImg1[138],OutputImg1[137],OutputImg1[136],
                      OutputImg1[135],OutputImg1[134],OutputImg1[133],
                      OutputImg1[132],OutputImg1[131],OutputImg1[130],
                      OutputImg1[129],OutputImg1[128]}), .EN (nx23796), .F ({
                      ImgReg0IN_143,ImgReg0IN_142,ImgReg0IN_141,ImgReg0IN_140,
                      ImgReg0IN_139,ImgReg0IN_138,ImgReg0IN_137,ImgReg0IN_136,
                      ImgReg0IN_135,ImgReg0IN_134,ImgReg0IN_133,ImgReg0IN_132,
                      ImgReg0IN_131,ImgReg0IN_130,ImgReg0IN_129,ImgReg0IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState1U (.D ({OutputImg2[143],OutputImg2[142],
                      OutputImg2[141],OutputImg2[140],OutputImg2[139],
                      OutputImg2[138],OutputImg2[137],OutputImg2[136],
                      OutputImg2[135],OutputImg2[134],OutputImg2[133],
                      OutputImg2[132],OutputImg2[131],OutputImg2[130],
                      OutputImg2[129],OutputImg2[128]}), .EN (nx23796), .F ({
                      ImgReg1IN_143,ImgReg1IN_142,ImgReg1IN_141,ImgReg1IN_140,
                      ImgReg1IN_139,ImgReg1IN_138,ImgReg1IN_137,ImgReg1IN_136,
                      ImgReg1IN_135,ImgReg1IN_134,ImgReg1IN_133,ImgReg1IN_132,
                      ImgReg1IN_131,ImgReg1IN_130,ImgReg1IN_129,ImgReg1IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState2U (.D ({OutputImg3[143],OutputImg3[142],
                      OutputImg3[141],OutputImg3[140],OutputImg3[139],
                      OutputImg3[138],OutputImg3[137],OutputImg3[136],
                      OutputImg3[135],OutputImg3[134],OutputImg3[133],
                      OutputImg3[132],OutputImg3[131],OutputImg3[130],
                      OutputImg3[129],OutputImg3[128]}), .EN (nx23798), .F ({
                      ImgReg2IN_143,ImgReg2IN_142,ImgReg2IN_141,ImgReg2IN_140,
                      ImgReg2IN_139,ImgReg2IN_138,ImgReg2IN_137,ImgReg2IN_136,
                      ImgReg2IN_135,ImgReg2IN_134,ImgReg2IN_133,ImgReg2IN_132,
                      ImgReg2IN_131,ImgReg2IN_130,ImgReg2IN_129,ImgReg2IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState3U (.D ({OutputImg4[143],OutputImg4[142],
                      OutputImg4[141],OutputImg4[140],OutputImg4[139],
                      OutputImg4[138],OutputImg4[137],OutputImg4[136],
                      OutputImg4[135],OutputImg4[134],OutputImg4[133],
                      OutputImg4[132],OutputImg4[131],OutputImg4[130],
                      OutputImg4[129],OutputImg4[128]}), .EN (nx23798), .F ({
                      ImgReg3IN_143,ImgReg3IN_142,ImgReg3IN_141,ImgReg3IN_140,
                      ImgReg3IN_139,ImgReg3IN_138,ImgReg3IN_137,ImgReg3IN_136,
                      ImgReg3IN_135,ImgReg3IN_134,ImgReg3IN_133,ImgReg3IN_132,
                      ImgReg3IN_131,ImgReg3IN_130,ImgReg3IN_129,ImgReg3IN_128})
                      ) ;
    triStateBuffer_16 loop3_8_TriState4U (.D ({OutputImg5[143],OutputImg5[142],
                      OutputImg5[141],OutputImg5[140],OutputImg5[139],
                      OutputImg5[138],OutputImg5[137],OutputImg5[136],
                      OutputImg5[135],OutputImg5[134],OutputImg5[133],
                      OutputImg5[132],OutputImg5[131],OutputImg5[130],
                      OutputImg5[129],OutputImg5[128]}), .EN (nx23798), .F ({
                      ImgReg4IN_143,ImgReg4IN_142,ImgReg4IN_141,ImgReg4IN_140,
                      ImgReg4IN_139,ImgReg4IN_138,ImgReg4IN_137,ImgReg4IN_136,
                      ImgReg4IN_135,ImgReg4IN_134,ImgReg4IN_133,ImgReg4IN_132,
                      ImgReg4IN_131,ImgReg4IN_130,ImgReg4IN_129,ImgReg4IN_128})
                      ) ;
    nBitRegister_16 loop3_8_reg1 (.D ({ImgReg0IN_143,ImgReg0IN_142,ImgReg0IN_141
                    ,ImgReg0IN_140,ImgReg0IN_139,ImgReg0IN_138,ImgReg0IN_137,
                    ImgReg0IN_136,ImgReg0IN_135,ImgReg0IN_134,ImgReg0IN_133,
                    ImgReg0IN_132,ImgReg0IN_131,ImgReg0IN_130,ImgReg0IN_129,
                    ImgReg0IN_128}), .CLK (nx23876), .RST (RST), .EN (nx23720), 
                    .Q ({OutputImg0[143],OutputImg0[142],OutputImg0[141],
                    OutputImg0[140],OutputImg0[139],OutputImg0[138],
                    OutputImg0[137],OutputImg0[136],OutputImg0[135],
                    OutputImg0[134],OutputImg0[133],OutputImg0[132],
                    OutputImg0[131],OutputImg0[130],OutputImg0[129],
                    OutputImg0[128]})) ;
    nBitRegister_16 loop3_8_reg2 (.D ({ImgReg1IN_143,ImgReg1IN_142,ImgReg1IN_141
                    ,ImgReg1IN_140,ImgReg1IN_139,ImgReg1IN_138,ImgReg1IN_137,
                    ImgReg1IN_136,ImgReg1IN_135,ImgReg1IN_134,ImgReg1IN_133,
                    ImgReg1IN_132,ImgReg1IN_131,ImgReg1IN_130,ImgReg1IN_129,
                    ImgReg1IN_128}), .CLK (nx23878), .RST (RST), .EN (nx23730), 
                    .Q ({OutputImg1[143],OutputImg1[142],OutputImg1[141],
                    OutputImg1[140],OutputImg1[139],OutputImg1[138],
                    OutputImg1[137],OutputImg1[136],OutputImg1[135],
                    OutputImg1[134],OutputImg1[133],OutputImg1[132],
                    OutputImg1[131],OutputImg1[130],OutputImg1[129],
                    OutputImg1[128]})) ;
    nBitRegister_16 loop3_8_reg3 (.D ({ImgReg2IN_143,ImgReg2IN_142,ImgReg2IN_141
                    ,ImgReg2IN_140,ImgReg2IN_139,ImgReg2IN_138,ImgReg2IN_137,
                    ImgReg2IN_136,ImgReg2IN_135,ImgReg2IN_134,ImgReg2IN_133,
                    ImgReg2IN_132,ImgReg2IN_131,ImgReg2IN_130,ImgReg2IN_129,
                    ImgReg2IN_128}), .CLK (nx23878), .RST (RST), .EN (nx23740), 
                    .Q ({OutputImg2[143],OutputImg2[142],OutputImg2[141],
                    OutputImg2[140],OutputImg2[139],OutputImg2[138],
                    OutputImg2[137],OutputImg2[136],OutputImg2[135],
                    OutputImg2[134],OutputImg2[133],OutputImg2[132],
                    OutputImg2[131],OutputImg2[130],OutputImg2[129],
                    OutputImg2[128]})) ;
    nBitRegister_16 loop3_8_reg4 (.D ({ImgReg3IN_143,ImgReg3IN_142,ImgReg3IN_141
                    ,ImgReg3IN_140,ImgReg3IN_139,ImgReg3IN_138,ImgReg3IN_137,
                    ImgReg3IN_136,ImgReg3IN_135,ImgReg3IN_134,ImgReg3IN_133,
                    ImgReg3IN_132,ImgReg3IN_131,ImgReg3IN_130,ImgReg3IN_129,
                    ImgReg3IN_128}), .CLK (nx23880), .RST (RST), .EN (nx23750), 
                    .Q ({OutputImg3[143],OutputImg3[142],OutputImg3[141],
                    OutputImg3[140],OutputImg3[139],OutputImg3[138],
                    OutputImg3[137],OutputImg3[136],OutputImg3[135],
                    OutputImg3[134],OutputImg3[133],OutputImg3[132],
                    OutputImg3[131],OutputImg3[130],OutputImg3[129],
                    OutputImg3[128]})) ;
    nBitRegister_16 loop3_8_reg5 (.D ({ImgReg4IN_143,ImgReg4IN_142,ImgReg4IN_141
                    ,ImgReg4IN_140,ImgReg4IN_139,ImgReg4IN_138,ImgReg4IN_137,
                    ImgReg4IN_136,ImgReg4IN_135,ImgReg4IN_134,ImgReg4IN_133,
                    ImgReg4IN_132,ImgReg4IN_131,ImgReg4IN_130,ImgReg4IN_129,
                    ImgReg4IN_128}), .CLK (nx23880), .RST (RST), .EN (nx23760), 
                    .Q ({OutputImg4[143],OutputImg4[142],OutputImg4[141],
                    OutputImg4[140],OutputImg4[139],OutputImg4[138],
                    OutputImg4[137],OutputImg4[136],OutputImg4[135],
                    OutputImg4[134],OutputImg4[133],OutputImg4[132],
                    OutputImg4[131],OutputImg4[130],OutputImg4[129],
                    OutputImg4[128]})) ;
    nBitRegister_16 loop3_8_reg6 (.D ({ImgReg5IN_143,ImgReg5IN_142,ImgReg5IN_141
                    ,ImgReg5IN_140,ImgReg5IN_139,ImgReg5IN_138,ImgReg5IN_137,
                    ImgReg5IN_136,ImgReg5IN_135,ImgReg5IN_134,ImgReg5IN_133,
                    ImgReg5IN_132,ImgReg5IN_131,ImgReg5IN_130,ImgReg5IN_129,
                    ImgReg5IN_128}), .CLK (nx23882), .RST (RST), .EN (nx23770), 
                    .Q ({OutputImg5[143],OutputImg5[142],OutputImg5[141],
                    OutputImg5[140],OutputImg5[139],OutputImg5[138],
                    OutputImg5[137],OutputImg5[136],OutputImg5[135],
                    OutputImg5[134],OutputImg5[133],OutputImg5[132],
                    OutputImg5[131],OutputImg5[130],OutputImg5[129],
                    OutputImg5[128]})) ;
    triStateBuffer_16 loop3_9_TriState0L (.D ({OutputImg0[175],OutputImg0[174],
                      OutputImg0[173],OutputImg0[172],OutputImg0[171],
                      OutputImg0[170],OutputImg0[169],OutputImg0[168],
                      OutputImg0[167],OutputImg0[166],OutputImg0[165],
                      OutputImg0[164],OutputImg0[163],OutputImg0[162],
                      OutputImg0[161],OutputImg0[160]}), .EN (nx23680), .F ({
                      ImgReg0IN_159,ImgReg0IN_158,ImgReg0IN_157,ImgReg0IN_156,
                      ImgReg0IN_155,ImgReg0IN_154,ImgReg0IN_153,ImgReg0IN_152,
                      ImgReg0IN_151,ImgReg0IN_150,ImgReg0IN_149,ImgReg0IN_148,
                      ImgReg0IN_147,ImgReg0IN_146,ImgReg0IN_145,ImgReg0IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState1L (.D ({OutputImg1[175],OutputImg1[174],
                      OutputImg1[173],OutputImg1[172],OutputImg1[171],
                      OutputImg1[170],OutputImg1[169],OutputImg1[168],
                      OutputImg1[167],OutputImg1[166],OutputImg1[165],
                      OutputImg1[164],OutputImg1[163],OutputImg1[162],
                      OutputImg1[161],OutputImg1[160]}), .EN (nx23680), .F ({
                      ImgReg1IN_159,ImgReg1IN_158,ImgReg1IN_157,ImgReg1IN_156,
                      ImgReg1IN_155,ImgReg1IN_154,ImgReg1IN_153,ImgReg1IN_152,
                      ImgReg1IN_151,ImgReg1IN_150,ImgReg1IN_149,ImgReg1IN_148,
                      ImgReg1IN_147,ImgReg1IN_146,ImgReg1IN_145,ImgReg1IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState2L (.D ({OutputImg2[175],OutputImg2[174],
                      OutputImg2[173],OutputImg2[172],OutputImg2[171],
                      OutputImg2[170],OutputImg2[169],OutputImg2[168],
                      OutputImg2[167],OutputImg2[166],OutputImg2[165],
                      OutputImg2[164],OutputImg2[163],OutputImg2[162],
                      OutputImg2[161],OutputImg2[160]}), .EN (nx23682), .F ({
                      ImgReg2IN_159,ImgReg2IN_158,ImgReg2IN_157,ImgReg2IN_156,
                      ImgReg2IN_155,ImgReg2IN_154,ImgReg2IN_153,ImgReg2IN_152,
                      ImgReg2IN_151,ImgReg2IN_150,ImgReg2IN_149,ImgReg2IN_148,
                      ImgReg2IN_147,ImgReg2IN_146,ImgReg2IN_145,ImgReg2IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState3L (.D ({OutputImg3[175],OutputImg3[174],
                      OutputImg3[173],OutputImg3[172],OutputImg3[171],
                      OutputImg3[170],OutputImg3[169],OutputImg3[168],
                      OutputImg3[167],OutputImg3[166],OutputImg3[165],
                      OutputImg3[164],OutputImg3[163],OutputImg3[162],
                      OutputImg3[161],OutputImg3[160]}), .EN (nx23682), .F ({
                      ImgReg3IN_159,ImgReg3IN_158,ImgReg3IN_157,ImgReg3IN_156,
                      ImgReg3IN_155,ImgReg3IN_154,ImgReg3IN_153,ImgReg3IN_152,
                      ImgReg3IN_151,ImgReg3IN_150,ImgReg3IN_149,ImgReg3IN_148,
                      ImgReg3IN_147,ImgReg3IN_146,ImgReg3IN_145,ImgReg3IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState4L (.D ({OutputImg4[175],OutputImg4[174],
                      OutputImg4[173],OutputImg4[172],OutputImg4[171],
                      OutputImg4[170],OutputImg4[169],OutputImg4[168],
                      OutputImg4[167],OutputImg4[166],OutputImg4[165],
                      OutputImg4[164],OutputImg4[163],OutputImg4[162],
                      OutputImg4[161],OutputImg4[160]}), .EN (nx23682), .F ({
                      ImgReg4IN_159,ImgReg4IN_158,ImgReg4IN_157,ImgReg4IN_156,
                      ImgReg4IN_155,ImgReg4IN_154,ImgReg4IN_153,ImgReg4IN_152,
                      ImgReg4IN_151,ImgReg4IN_150,ImgReg4IN_149,ImgReg4IN_148,
                      ImgReg4IN_147,ImgReg4IN_146,ImgReg4IN_145,ImgReg4IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState5L (.D ({OutputImg5[175],OutputImg5[174],
                      OutputImg5[173],OutputImg5[172],OutputImg5[171],
                      OutputImg5[170],OutputImg5[169],OutputImg5[168],
                      OutputImg5[167],OutputImg5[166],OutputImg5[165],
                      OutputImg5[164],OutputImg5[163],OutputImg5[162],
                      OutputImg5[161],OutputImg5[160]}), .EN (nx23682), .F ({
                      ImgReg5IN_159,ImgReg5IN_158,ImgReg5IN_157,ImgReg5IN_156,
                      ImgReg5IN_155,ImgReg5IN_154,ImgReg5IN_153,ImgReg5IN_152,
                      ImgReg5IN_151,ImgReg5IN_150,ImgReg5IN_149,ImgReg5IN_148,
                      ImgReg5IN_147,ImgReg5IN_146,ImgReg5IN_145,ImgReg5IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState0N (.D ({DATA[159],DATA[158],DATA[157],
                      DATA[156],DATA[155],DATA[154],DATA[153],DATA[152],
                      DATA[151],DATA[150],DATA[149],DATA[148],DATA[147],
                      DATA[146],DATA[145],DATA[144]}), .EN (nx23656), .F ({
                      ImgReg0IN_159,ImgReg0IN_158,ImgReg0IN_157,ImgReg0IN_156,
                      ImgReg0IN_155,ImgReg0IN_154,ImgReg0IN_153,ImgReg0IN_152,
                      ImgReg0IN_151,ImgReg0IN_150,ImgReg0IN_149,ImgReg0IN_148,
                      ImgReg0IN_147,ImgReg0IN_146,ImgReg0IN_145,ImgReg0IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState1N (.D ({DATA[159],DATA[158],DATA[157],
                      DATA[156],DATA[155],DATA[154],DATA[153],DATA[152],
                      DATA[151],DATA[150],DATA[149],DATA[148],DATA[147],
                      DATA[146],DATA[145],DATA[144]}), .EN (nx23644), .F ({
                      ImgReg1IN_159,ImgReg1IN_158,ImgReg1IN_157,ImgReg1IN_156,
                      ImgReg1IN_155,ImgReg1IN_154,ImgReg1IN_153,ImgReg1IN_152,
                      ImgReg1IN_151,ImgReg1IN_150,ImgReg1IN_149,ImgReg1IN_148,
                      ImgReg1IN_147,ImgReg1IN_146,ImgReg1IN_145,ImgReg1IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState2N (.D ({DATA[159],DATA[158],DATA[157],
                      DATA[156],DATA[155],DATA[154],DATA[153],DATA[152],
                      DATA[151],DATA[150],DATA[149],DATA[148],DATA[147],
                      DATA[146],DATA[145],DATA[144]}), .EN (nx23632), .F ({
                      ImgReg2IN_159,ImgReg2IN_158,ImgReg2IN_157,ImgReg2IN_156,
                      ImgReg2IN_155,ImgReg2IN_154,ImgReg2IN_153,ImgReg2IN_152,
                      ImgReg2IN_151,ImgReg2IN_150,ImgReg2IN_149,ImgReg2IN_148,
                      ImgReg2IN_147,ImgReg2IN_146,ImgReg2IN_145,ImgReg2IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState3N (.D ({DATA[159],DATA[158],DATA[157],
                      DATA[156],DATA[155],DATA[154],DATA[153],DATA[152],
                      DATA[151],DATA[150],DATA[149],DATA[148],DATA[147],
                      DATA[146],DATA[145],DATA[144]}), .EN (nx23620), .F ({
                      ImgReg3IN_159,ImgReg3IN_158,ImgReg3IN_157,ImgReg3IN_156,
                      ImgReg3IN_155,ImgReg3IN_154,ImgReg3IN_153,ImgReg3IN_152,
                      ImgReg3IN_151,ImgReg3IN_150,ImgReg3IN_149,ImgReg3IN_148,
                      ImgReg3IN_147,ImgReg3IN_146,ImgReg3IN_145,ImgReg3IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState4N (.D ({DATA[159],DATA[158],DATA[157],
                      DATA[156],DATA[155],DATA[154],DATA[153],DATA[152],
                      DATA[151],DATA[150],DATA[149],DATA[148],DATA[147],
                      DATA[146],DATA[145],DATA[144]}), .EN (nx23608), .F ({
                      ImgReg4IN_159,ImgReg4IN_158,ImgReg4IN_157,ImgReg4IN_156,
                      ImgReg4IN_155,ImgReg4IN_154,ImgReg4IN_153,ImgReg4IN_152,
                      ImgReg4IN_151,ImgReg4IN_150,ImgReg4IN_149,ImgReg4IN_148,
                      ImgReg4IN_147,ImgReg4IN_146,ImgReg4IN_145,ImgReg4IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState5N (.D ({DATA[159],DATA[158],DATA[157],
                      DATA[156],DATA[155],DATA[154],DATA[153],DATA[152],
                      DATA[151],DATA[150],DATA[149],DATA[148],DATA[147],
                      DATA[146],DATA[145],DATA[144]}), .EN (nx23596), .F ({
                      ImgReg5IN_159,ImgReg5IN_158,ImgReg5IN_157,ImgReg5IN_156,
                      ImgReg5IN_155,ImgReg5IN_154,ImgReg5IN_153,ImgReg5IN_152,
                      ImgReg5IN_151,ImgReg5IN_150,ImgReg5IN_149,ImgReg5IN_148,
                      ImgReg5IN_147,ImgReg5IN_146,ImgReg5IN_145,ImgReg5IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState0U (.D ({OutputImg1[159],OutputImg1[158],
                      OutputImg1[157],OutputImg1[156],OutputImg1[155],
                      OutputImg1[154],OutputImg1[153],OutputImg1[152],
                      OutputImg1[151],OutputImg1[150],OutputImg1[149],
                      OutputImg1[148],OutputImg1[147],OutputImg1[146],
                      OutputImg1[145],OutputImg1[144]}), .EN (nx23798), .F ({
                      ImgReg0IN_159,ImgReg0IN_158,ImgReg0IN_157,ImgReg0IN_156,
                      ImgReg0IN_155,ImgReg0IN_154,ImgReg0IN_153,ImgReg0IN_152,
                      ImgReg0IN_151,ImgReg0IN_150,ImgReg0IN_149,ImgReg0IN_148,
                      ImgReg0IN_147,ImgReg0IN_146,ImgReg0IN_145,ImgReg0IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState1U (.D ({OutputImg2[159],OutputImg2[158],
                      OutputImg2[157],OutputImg2[156],OutputImg2[155],
                      OutputImg2[154],OutputImg2[153],OutputImg2[152],
                      OutputImg2[151],OutputImg2[150],OutputImg2[149],
                      OutputImg2[148],OutputImg2[147],OutputImg2[146],
                      OutputImg2[145],OutputImg2[144]}), .EN (nx23798), .F ({
                      ImgReg1IN_159,ImgReg1IN_158,ImgReg1IN_157,ImgReg1IN_156,
                      ImgReg1IN_155,ImgReg1IN_154,ImgReg1IN_153,ImgReg1IN_152,
                      ImgReg1IN_151,ImgReg1IN_150,ImgReg1IN_149,ImgReg1IN_148,
                      ImgReg1IN_147,ImgReg1IN_146,ImgReg1IN_145,ImgReg1IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState2U (.D ({OutputImg3[159],OutputImg3[158],
                      OutputImg3[157],OutputImg3[156],OutputImg3[155],
                      OutputImg3[154],OutputImg3[153],OutputImg3[152],
                      OutputImg3[151],OutputImg3[150],OutputImg3[149],
                      OutputImg3[148],OutputImg3[147],OutputImg3[146],
                      OutputImg3[145],OutputImg3[144]}), .EN (nx23798), .F ({
                      ImgReg2IN_159,ImgReg2IN_158,ImgReg2IN_157,ImgReg2IN_156,
                      ImgReg2IN_155,ImgReg2IN_154,ImgReg2IN_153,ImgReg2IN_152,
                      ImgReg2IN_151,ImgReg2IN_150,ImgReg2IN_149,ImgReg2IN_148,
                      ImgReg2IN_147,ImgReg2IN_146,ImgReg2IN_145,ImgReg2IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState3U (.D ({OutputImg4[159],OutputImg4[158],
                      OutputImg4[157],OutputImg4[156],OutputImg4[155],
                      OutputImg4[154],OutputImg4[153],OutputImg4[152],
                      OutputImg4[151],OutputImg4[150],OutputImg4[149],
                      OutputImg4[148],OutputImg4[147],OutputImg4[146],
                      OutputImg4[145],OutputImg4[144]}), .EN (nx23798), .F ({
                      ImgReg3IN_159,ImgReg3IN_158,ImgReg3IN_157,ImgReg3IN_156,
                      ImgReg3IN_155,ImgReg3IN_154,ImgReg3IN_153,ImgReg3IN_152,
                      ImgReg3IN_151,ImgReg3IN_150,ImgReg3IN_149,ImgReg3IN_148,
                      ImgReg3IN_147,ImgReg3IN_146,ImgReg3IN_145,ImgReg3IN_144})
                      ) ;
    triStateBuffer_16 loop3_9_TriState4U (.D ({OutputImg5[159],OutputImg5[158],
                      OutputImg5[157],OutputImg5[156],OutputImg5[155],
                      OutputImg5[154],OutputImg5[153],OutputImg5[152],
                      OutputImg5[151],OutputImg5[150],OutputImg5[149],
                      OutputImg5[148],OutputImg5[147],OutputImg5[146],
                      OutputImg5[145],OutputImg5[144]}), .EN (nx23800), .F ({
                      ImgReg4IN_159,ImgReg4IN_158,ImgReg4IN_157,ImgReg4IN_156,
                      ImgReg4IN_155,ImgReg4IN_154,ImgReg4IN_153,ImgReg4IN_152,
                      ImgReg4IN_151,ImgReg4IN_150,ImgReg4IN_149,ImgReg4IN_148,
                      ImgReg4IN_147,ImgReg4IN_146,ImgReg4IN_145,ImgReg4IN_144})
                      ) ;
    nBitRegister_16 loop3_9_reg1 (.D ({ImgReg0IN_159,ImgReg0IN_158,ImgReg0IN_157
                    ,ImgReg0IN_156,ImgReg0IN_155,ImgReg0IN_154,ImgReg0IN_153,
                    ImgReg0IN_152,ImgReg0IN_151,ImgReg0IN_150,ImgReg0IN_149,
                    ImgReg0IN_148,ImgReg0IN_147,ImgReg0IN_146,ImgReg0IN_145,
                    ImgReg0IN_144}), .CLK (nx23882), .RST (RST), .EN (nx23720), 
                    .Q ({OutputImg0[159],OutputImg0[158],OutputImg0[157],
                    OutputImg0[156],OutputImg0[155],OutputImg0[154],
                    OutputImg0[153],OutputImg0[152],OutputImg0[151],
                    OutputImg0[150],OutputImg0[149],OutputImg0[148],
                    OutputImg0[147],OutputImg0[146],OutputImg0[145],
                    OutputImg0[144]})) ;
    nBitRegister_16 loop3_9_reg2 (.D ({ImgReg1IN_159,ImgReg1IN_158,ImgReg1IN_157
                    ,ImgReg1IN_156,ImgReg1IN_155,ImgReg1IN_154,ImgReg1IN_153,
                    ImgReg1IN_152,ImgReg1IN_151,ImgReg1IN_150,ImgReg1IN_149,
                    ImgReg1IN_148,ImgReg1IN_147,ImgReg1IN_146,ImgReg1IN_145,
                    ImgReg1IN_144}), .CLK (nx23884), .RST (RST), .EN (nx23730), 
                    .Q ({OutputImg1[159],OutputImg1[158],OutputImg1[157],
                    OutputImg1[156],OutputImg1[155],OutputImg1[154],
                    OutputImg1[153],OutputImg1[152],OutputImg1[151],
                    OutputImg1[150],OutputImg1[149],OutputImg1[148],
                    OutputImg1[147],OutputImg1[146],OutputImg1[145],
                    OutputImg1[144]})) ;
    nBitRegister_16 loop3_9_reg3 (.D ({ImgReg2IN_159,ImgReg2IN_158,ImgReg2IN_157
                    ,ImgReg2IN_156,ImgReg2IN_155,ImgReg2IN_154,ImgReg2IN_153,
                    ImgReg2IN_152,ImgReg2IN_151,ImgReg2IN_150,ImgReg2IN_149,
                    ImgReg2IN_148,ImgReg2IN_147,ImgReg2IN_146,ImgReg2IN_145,
                    ImgReg2IN_144}), .CLK (nx23884), .RST (RST), .EN (nx23740), 
                    .Q ({OutputImg2[159],OutputImg2[158],OutputImg2[157],
                    OutputImg2[156],OutputImg2[155],OutputImg2[154],
                    OutputImg2[153],OutputImg2[152],OutputImg2[151],
                    OutputImg2[150],OutputImg2[149],OutputImg2[148],
                    OutputImg2[147],OutputImg2[146],OutputImg2[145],
                    OutputImg2[144]})) ;
    nBitRegister_16 loop3_9_reg4 (.D ({ImgReg3IN_159,ImgReg3IN_158,ImgReg3IN_157
                    ,ImgReg3IN_156,ImgReg3IN_155,ImgReg3IN_154,ImgReg3IN_153,
                    ImgReg3IN_152,ImgReg3IN_151,ImgReg3IN_150,ImgReg3IN_149,
                    ImgReg3IN_148,ImgReg3IN_147,ImgReg3IN_146,ImgReg3IN_145,
                    ImgReg3IN_144}), .CLK (nx23886), .RST (RST), .EN (nx23750), 
                    .Q ({OutputImg3[159],OutputImg3[158],OutputImg3[157],
                    OutputImg3[156],OutputImg3[155],OutputImg3[154],
                    OutputImg3[153],OutputImg3[152],OutputImg3[151],
                    OutputImg3[150],OutputImg3[149],OutputImg3[148],
                    OutputImg3[147],OutputImg3[146],OutputImg3[145],
                    OutputImg3[144]})) ;
    nBitRegister_16 loop3_9_reg5 (.D ({ImgReg4IN_159,ImgReg4IN_158,ImgReg4IN_157
                    ,ImgReg4IN_156,ImgReg4IN_155,ImgReg4IN_154,ImgReg4IN_153,
                    ImgReg4IN_152,ImgReg4IN_151,ImgReg4IN_150,ImgReg4IN_149,
                    ImgReg4IN_148,ImgReg4IN_147,ImgReg4IN_146,ImgReg4IN_145,
                    ImgReg4IN_144}), .CLK (nx23886), .RST (RST), .EN (nx23760), 
                    .Q ({OutputImg4[159],OutputImg4[158],OutputImg4[157],
                    OutputImg4[156],OutputImg4[155],OutputImg4[154],
                    OutputImg4[153],OutputImg4[152],OutputImg4[151],
                    OutputImg4[150],OutputImg4[149],OutputImg4[148],
                    OutputImg4[147],OutputImg4[146],OutputImg4[145],
                    OutputImg4[144]})) ;
    nBitRegister_16 loop3_9_reg6 (.D ({ImgReg5IN_159,ImgReg5IN_158,ImgReg5IN_157
                    ,ImgReg5IN_156,ImgReg5IN_155,ImgReg5IN_154,ImgReg5IN_153,
                    ImgReg5IN_152,ImgReg5IN_151,ImgReg5IN_150,ImgReg5IN_149,
                    ImgReg5IN_148,ImgReg5IN_147,ImgReg5IN_146,ImgReg5IN_145,
                    ImgReg5IN_144}), .CLK (nx23888), .RST (RST), .EN (nx23770), 
                    .Q ({OutputImg5[159],OutputImg5[158],OutputImg5[157],
                    OutputImg5[156],OutputImg5[155],OutputImg5[154],
                    OutputImg5[153],OutputImg5[152],OutputImg5[151],
                    OutputImg5[150],OutputImg5[149],OutputImg5[148],
                    OutputImg5[147],OutputImg5[146],OutputImg5[145],
                    OutputImg5[144]})) ;
    triStateBuffer_16 loop3_10_TriState0L (.D ({OutputImg0[191],OutputImg0[190],
                      OutputImg0[189],OutputImg0[188],OutputImg0[187],
                      OutputImg0[186],OutputImg0[185],OutputImg0[184],
                      OutputImg0[183],OutputImg0[182],OutputImg0[181],
                      OutputImg0[180],OutputImg0[179],OutputImg0[178],
                      OutputImg0[177],OutputImg0[176]}), .EN (nx23682), .F ({
                      ImgReg0IN_175,ImgReg0IN_174,ImgReg0IN_173,ImgReg0IN_172,
                      ImgReg0IN_171,ImgReg0IN_170,ImgReg0IN_169,ImgReg0IN_168,
                      ImgReg0IN_167,ImgReg0IN_166,ImgReg0IN_165,ImgReg0IN_164,
                      ImgReg0IN_163,ImgReg0IN_162,ImgReg0IN_161,ImgReg0IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState1L (.D ({OutputImg1[191],OutputImg1[190],
                      OutputImg1[189],OutputImg1[188],OutputImg1[187],
                      OutputImg1[186],OutputImg1[185],OutputImg1[184],
                      OutputImg1[183],OutputImg1[182],OutputImg1[181],
                      OutputImg1[180],OutputImg1[179],OutputImg1[178],
                      OutputImg1[177],OutputImg1[176]}), .EN (nx23682), .F ({
                      ImgReg1IN_175,ImgReg1IN_174,ImgReg1IN_173,ImgReg1IN_172,
                      ImgReg1IN_171,ImgReg1IN_170,ImgReg1IN_169,ImgReg1IN_168,
                      ImgReg1IN_167,ImgReg1IN_166,ImgReg1IN_165,ImgReg1IN_164,
                      ImgReg1IN_163,ImgReg1IN_162,ImgReg1IN_161,ImgReg1IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState2L (.D ({OutputImg2[191],OutputImg2[190],
                      OutputImg2[189],OutputImg2[188],OutputImg2[187],
                      OutputImg2[186],OutputImg2[185],OutputImg2[184],
                      OutputImg2[183],OutputImg2[182],OutputImg2[181],
                      OutputImg2[180],OutputImg2[179],OutputImg2[178],
                      OutputImg2[177],OutputImg2[176]}), .EN (nx23682), .F ({
                      ImgReg2IN_175,ImgReg2IN_174,ImgReg2IN_173,ImgReg2IN_172,
                      ImgReg2IN_171,ImgReg2IN_170,ImgReg2IN_169,ImgReg2IN_168,
                      ImgReg2IN_167,ImgReg2IN_166,ImgReg2IN_165,ImgReg2IN_164,
                      ImgReg2IN_163,ImgReg2IN_162,ImgReg2IN_161,ImgReg2IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState3L (.D ({OutputImg3[191],OutputImg3[190],
                      OutputImg3[189],OutputImg3[188],OutputImg3[187],
                      OutputImg3[186],OutputImg3[185],OutputImg3[184],
                      OutputImg3[183],OutputImg3[182],OutputImg3[181],
                      OutputImg3[180],OutputImg3[179],OutputImg3[178],
                      OutputImg3[177],OutputImg3[176]}), .EN (nx23684), .F ({
                      ImgReg3IN_175,ImgReg3IN_174,ImgReg3IN_173,ImgReg3IN_172,
                      ImgReg3IN_171,ImgReg3IN_170,ImgReg3IN_169,ImgReg3IN_168,
                      ImgReg3IN_167,ImgReg3IN_166,ImgReg3IN_165,ImgReg3IN_164,
                      ImgReg3IN_163,ImgReg3IN_162,ImgReg3IN_161,ImgReg3IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState4L (.D ({OutputImg4[191],OutputImg4[190],
                      OutputImg4[189],OutputImg4[188],OutputImg4[187],
                      OutputImg4[186],OutputImg4[185],OutputImg4[184],
                      OutputImg4[183],OutputImg4[182],OutputImg4[181],
                      OutputImg4[180],OutputImg4[179],OutputImg4[178],
                      OutputImg4[177],OutputImg4[176]}), .EN (nx23684), .F ({
                      ImgReg4IN_175,ImgReg4IN_174,ImgReg4IN_173,ImgReg4IN_172,
                      ImgReg4IN_171,ImgReg4IN_170,ImgReg4IN_169,ImgReg4IN_168,
                      ImgReg4IN_167,ImgReg4IN_166,ImgReg4IN_165,ImgReg4IN_164,
                      ImgReg4IN_163,ImgReg4IN_162,ImgReg4IN_161,ImgReg4IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState5L (.D ({OutputImg5[191],OutputImg5[190],
                      OutputImg5[189],OutputImg5[188],OutputImg5[187],
                      OutputImg5[186],OutputImg5[185],OutputImg5[184],
                      OutputImg5[183],OutputImg5[182],OutputImg5[181],
                      OutputImg5[180],OutputImg5[179],OutputImg5[178],
                      OutputImg5[177],OutputImg5[176]}), .EN (nx23684), .F ({
                      ImgReg5IN_175,ImgReg5IN_174,ImgReg5IN_173,ImgReg5IN_172,
                      ImgReg5IN_171,ImgReg5IN_170,ImgReg5IN_169,ImgReg5IN_168,
                      ImgReg5IN_167,ImgReg5IN_166,ImgReg5IN_165,ImgReg5IN_164,
                      ImgReg5IN_163,ImgReg5IN_162,ImgReg5IN_161,ImgReg5IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState0N (.D ({DATA[175],DATA[174],DATA[173],
                      DATA[172],DATA[171],DATA[170],DATA[169],DATA[168],
                      DATA[167],DATA[166],DATA[165],DATA[164],DATA[163],
                      DATA[162],DATA[161],DATA[160]}), .EN (nx23656), .F ({
                      ImgReg0IN_175,ImgReg0IN_174,ImgReg0IN_173,ImgReg0IN_172,
                      ImgReg0IN_171,ImgReg0IN_170,ImgReg0IN_169,ImgReg0IN_168,
                      ImgReg0IN_167,ImgReg0IN_166,ImgReg0IN_165,ImgReg0IN_164,
                      ImgReg0IN_163,ImgReg0IN_162,ImgReg0IN_161,ImgReg0IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState1N (.D ({DATA[175],DATA[174],DATA[173],
                      DATA[172],DATA[171],DATA[170],DATA[169],DATA[168],
                      DATA[167],DATA[166],DATA[165],DATA[164],DATA[163],
                      DATA[162],DATA[161],DATA[160]}), .EN (nx23644), .F ({
                      ImgReg1IN_175,ImgReg1IN_174,ImgReg1IN_173,ImgReg1IN_172,
                      ImgReg1IN_171,ImgReg1IN_170,ImgReg1IN_169,ImgReg1IN_168,
                      ImgReg1IN_167,ImgReg1IN_166,ImgReg1IN_165,ImgReg1IN_164,
                      ImgReg1IN_163,ImgReg1IN_162,ImgReg1IN_161,ImgReg1IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState2N (.D ({DATA[175],DATA[174],DATA[173],
                      DATA[172],DATA[171],DATA[170],DATA[169],DATA[168],
                      DATA[167],DATA[166],DATA[165],DATA[164],DATA[163],
                      DATA[162],DATA[161],DATA[160]}), .EN (nx23632), .F ({
                      ImgReg2IN_175,ImgReg2IN_174,ImgReg2IN_173,ImgReg2IN_172,
                      ImgReg2IN_171,ImgReg2IN_170,ImgReg2IN_169,ImgReg2IN_168,
                      ImgReg2IN_167,ImgReg2IN_166,ImgReg2IN_165,ImgReg2IN_164,
                      ImgReg2IN_163,ImgReg2IN_162,ImgReg2IN_161,ImgReg2IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState3N (.D ({DATA[175],DATA[174],DATA[173],
                      DATA[172],DATA[171],DATA[170],DATA[169],DATA[168],
                      DATA[167],DATA[166],DATA[165],DATA[164],DATA[163],
                      DATA[162],DATA[161],DATA[160]}), .EN (nx23620), .F ({
                      ImgReg3IN_175,ImgReg3IN_174,ImgReg3IN_173,ImgReg3IN_172,
                      ImgReg3IN_171,ImgReg3IN_170,ImgReg3IN_169,ImgReg3IN_168,
                      ImgReg3IN_167,ImgReg3IN_166,ImgReg3IN_165,ImgReg3IN_164,
                      ImgReg3IN_163,ImgReg3IN_162,ImgReg3IN_161,ImgReg3IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState4N (.D ({DATA[175],DATA[174],DATA[173],
                      DATA[172],DATA[171],DATA[170],DATA[169],DATA[168],
                      DATA[167],DATA[166],DATA[165],DATA[164],DATA[163],
                      DATA[162],DATA[161],DATA[160]}), .EN (nx23608), .F ({
                      ImgReg4IN_175,ImgReg4IN_174,ImgReg4IN_173,ImgReg4IN_172,
                      ImgReg4IN_171,ImgReg4IN_170,ImgReg4IN_169,ImgReg4IN_168,
                      ImgReg4IN_167,ImgReg4IN_166,ImgReg4IN_165,ImgReg4IN_164,
                      ImgReg4IN_163,ImgReg4IN_162,ImgReg4IN_161,ImgReg4IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState5N (.D ({DATA[175],DATA[174],DATA[173],
                      DATA[172],DATA[171],DATA[170],DATA[169],DATA[168],
                      DATA[167],DATA[166],DATA[165],DATA[164],DATA[163],
                      DATA[162],DATA[161],DATA[160]}), .EN (nx23596), .F ({
                      ImgReg5IN_175,ImgReg5IN_174,ImgReg5IN_173,ImgReg5IN_172,
                      ImgReg5IN_171,ImgReg5IN_170,ImgReg5IN_169,ImgReg5IN_168,
                      ImgReg5IN_167,ImgReg5IN_166,ImgReg5IN_165,ImgReg5IN_164,
                      ImgReg5IN_163,ImgReg5IN_162,ImgReg5IN_161,ImgReg5IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState0U (.D ({OutputImg1[175],OutputImg1[174],
                      OutputImg1[173],OutputImg1[172],OutputImg1[171],
                      OutputImg1[170],OutputImg1[169],OutputImg1[168],
                      OutputImg1[167],OutputImg1[166],OutputImg1[165],
                      OutputImg1[164],OutputImg1[163],OutputImg1[162],
                      OutputImg1[161],OutputImg1[160]}), .EN (nx23800), .F ({
                      ImgReg0IN_175,ImgReg0IN_174,ImgReg0IN_173,ImgReg0IN_172,
                      ImgReg0IN_171,ImgReg0IN_170,ImgReg0IN_169,ImgReg0IN_168,
                      ImgReg0IN_167,ImgReg0IN_166,ImgReg0IN_165,ImgReg0IN_164,
                      ImgReg0IN_163,ImgReg0IN_162,ImgReg0IN_161,ImgReg0IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState1U (.D ({OutputImg2[175],OutputImg2[174],
                      OutputImg2[173],OutputImg2[172],OutputImg2[171],
                      OutputImg2[170],OutputImg2[169],OutputImg2[168],
                      OutputImg2[167],OutputImg2[166],OutputImg2[165],
                      OutputImg2[164],OutputImg2[163],OutputImg2[162],
                      OutputImg2[161],OutputImg2[160]}), .EN (nx23800), .F ({
                      ImgReg1IN_175,ImgReg1IN_174,ImgReg1IN_173,ImgReg1IN_172,
                      ImgReg1IN_171,ImgReg1IN_170,ImgReg1IN_169,ImgReg1IN_168,
                      ImgReg1IN_167,ImgReg1IN_166,ImgReg1IN_165,ImgReg1IN_164,
                      ImgReg1IN_163,ImgReg1IN_162,ImgReg1IN_161,ImgReg1IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState2U (.D ({OutputImg3[175],OutputImg3[174],
                      OutputImg3[173],OutputImg3[172],OutputImg3[171],
                      OutputImg3[170],OutputImg3[169],OutputImg3[168],
                      OutputImg3[167],OutputImg3[166],OutputImg3[165],
                      OutputImg3[164],OutputImg3[163],OutputImg3[162],
                      OutputImg3[161],OutputImg3[160]}), .EN (nx23800), .F ({
                      ImgReg2IN_175,ImgReg2IN_174,ImgReg2IN_173,ImgReg2IN_172,
                      ImgReg2IN_171,ImgReg2IN_170,ImgReg2IN_169,ImgReg2IN_168,
                      ImgReg2IN_167,ImgReg2IN_166,ImgReg2IN_165,ImgReg2IN_164,
                      ImgReg2IN_163,ImgReg2IN_162,ImgReg2IN_161,ImgReg2IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState3U (.D ({OutputImg4[175],OutputImg4[174],
                      OutputImg4[173],OutputImg4[172],OutputImg4[171],
                      OutputImg4[170],OutputImg4[169],OutputImg4[168],
                      OutputImg4[167],OutputImg4[166],OutputImg4[165],
                      OutputImg4[164],OutputImg4[163],OutputImg4[162],
                      OutputImg4[161],OutputImg4[160]}), .EN (nx23800), .F ({
                      ImgReg3IN_175,ImgReg3IN_174,ImgReg3IN_173,ImgReg3IN_172,
                      ImgReg3IN_171,ImgReg3IN_170,ImgReg3IN_169,ImgReg3IN_168,
                      ImgReg3IN_167,ImgReg3IN_166,ImgReg3IN_165,ImgReg3IN_164,
                      ImgReg3IN_163,ImgReg3IN_162,ImgReg3IN_161,ImgReg3IN_160})
                      ) ;
    triStateBuffer_16 loop3_10_TriState4U (.D ({OutputImg5[175],OutputImg5[174],
                      OutputImg5[173],OutputImg5[172],OutputImg5[171],
                      OutputImg5[170],OutputImg5[169],OutputImg5[168],
                      OutputImg5[167],OutputImg5[166],OutputImg5[165],
                      OutputImg5[164],OutputImg5[163],OutputImg5[162],
                      OutputImg5[161],OutputImg5[160]}), .EN (nx23800), .F ({
                      ImgReg4IN_175,ImgReg4IN_174,ImgReg4IN_173,ImgReg4IN_172,
                      ImgReg4IN_171,ImgReg4IN_170,ImgReg4IN_169,ImgReg4IN_168,
                      ImgReg4IN_167,ImgReg4IN_166,ImgReg4IN_165,ImgReg4IN_164,
                      ImgReg4IN_163,ImgReg4IN_162,ImgReg4IN_161,ImgReg4IN_160})
                      ) ;
    nBitRegister_16 loop3_10_reg1 (.D ({ImgReg0IN_175,ImgReg0IN_174,
                    ImgReg0IN_173,ImgReg0IN_172,ImgReg0IN_171,ImgReg0IN_170,
                    ImgReg0IN_169,ImgReg0IN_168,ImgReg0IN_167,ImgReg0IN_166,
                    ImgReg0IN_165,ImgReg0IN_164,ImgReg0IN_163,ImgReg0IN_162,
                    ImgReg0IN_161,ImgReg0IN_160}), .CLK (nx23888), .RST (RST), .EN (
                    nx23720), .Q ({OutputImg0[175],OutputImg0[174],
                    OutputImg0[173],OutputImg0[172],OutputImg0[171],
                    OutputImg0[170],OutputImg0[169],OutputImg0[168],
                    OutputImg0[167],OutputImg0[166],OutputImg0[165],
                    OutputImg0[164],OutputImg0[163],OutputImg0[162],
                    OutputImg0[161],OutputImg0[160]})) ;
    nBitRegister_16 loop3_10_reg2 (.D ({ImgReg1IN_175,ImgReg1IN_174,
                    ImgReg1IN_173,ImgReg1IN_172,ImgReg1IN_171,ImgReg1IN_170,
                    ImgReg1IN_169,ImgReg1IN_168,ImgReg1IN_167,ImgReg1IN_166,
                    ImgReg1IN_165,ImgReg1IN_164,ImgReg1IN_163,ImgReg1IN_162,
                    ImgReg1IN_161,ImgReg1IN_160}), .CLK (nx23890), .RST (RST), .EN (
                    nx23730), .Q ({OutputImg1[175],OutputImg1[174],
                    OutputImg1[173],OutputImg1[172],OutputImg1[171],
                    OutputImg1[170],OutputImg1[169],OutputImg1[168],
                    OutputImg1[167],OutputImg1[166],OutputImg1[165],
                    OutputImg1[164],OutputImg1[163],OutputImg1[162],
                    OutputImg1[161],OutputImg1[160]})) ;
    nBitRegister_16 loop3_10_reg3 (.D ({ImgReg2IN_175,ImgReg2IN_174,
                    ImgReg2IN_173,ImgReg2IN_172,ImgReg2IN_171,ImgReg2IN_170,
                    ImgReg2IN_169,ImgReg2IN_168,ImgReg2IN_167,ImgReg2IN_166,
                    ImgReg2IN_165,ImgReg2IN_164,ImgReg2IN_163,ImgReg2IN_162,
                    ImgReg2IN_161,ImgReg2IN_160}), .CLK (nx23890), .RST (RST), .EN (
                    nx23740), .Q ({OutputImg2[175],OutputImg2[174],
                    OutputImg2[173],OutputImg2[172],OutputImg2[171],
                    OutputImg2[170],OutputImg2[169],OutputImg2[168],
                    OutputImg2[167],OutputImg2[166],OutputImg2[165],
                    OutputImg2[164],OutputImg2[163],OutputImg2[162],
                    OutputImg2[161],OutputImg2[160]})) ;
    nBitRegister_16 loop3_10_reg4 (.D ({ImgReg3IN_175,ImgReg3IN_174,
                    ImgReg3IN_173,ImgReg3IN_172,ImgReg3IN_171,ImgReg3IN_170,
                    ImgReg3IN_169,ImgReg3IN_168,ImgReg3IN_167,ImgReg3IN_166,
                    ImgReg3IN_165,ImgReg3IN_164,ImgReg3IN_163,ImgReg3IN_162,
                    ImgReg3IN_161,ImgReg3IN_160}), .CLK (nx23892), .RST (RST), .EN (
                    nx23750), .Q ({OutputImg3[175],OutputImg3[174],
                    OutputImg3[173],OutputImg3[172],OutputImg3[171],
                    OutputImg3[170],OutputImg3[169],OutputImg3[168],
                    OutputImg3[167],OutputImg3[166],OutputImg3[165],
                    OutputImg3[164],OutputImg3[163],OutputImg3[162],
                    OutputImg3[161],OutputImg3[160]})) ;
    nBitRegister_16 loop3_10_reg5 (.D ({ImgReg4IN_175,ImgReg4IN_174,
                    ImgReg4IN_173,ImgReg4IN_172,ImgReg4IN_171,ImgReg4IN_170,
                    ImgReg4IN_169,ImgReg4IN_168,ImgReg4IN_167,ImgReg4IN_166,
                    ImgReg4IN_165,ImgReg4IN_164,ImgReg4IN_163,ImgReg4IN_162,
                    ImgReg4IN_161,ImgReg4IN_160}), .CLK (nx23892), .RST (RST), .EN (
                    nx23760), .Q ({OutputImg4[175],OutputImg4[174],
                    OutputImg4[173],OutputImg4[172],OutputImg4[171],
                    OutputImg4[170],OutputImg4[169],OutputImg4[168],
                    OutputImg4[167],OutputImg4[166],OutputImg4[165],
                    OutputImg4[164],OutputImg4[163],OutputImg4[162],
                    OutputImg4[161],OutputImg4[160]})) ;
    nBitRegister_16 loop3_10_reg6 (.D ({ImgReg5IN_175,ImgReg5IN_174,
                    ImgReg5IN_173,ImgReg5IN_172,ImgReg5IN_171,ImgReg5IN_170,
                    ImgReg5IN_169,ImgReg5IN_168,ImgReg5IN_167,ImgReg5IN_166,
                    ImgReg5IN_165,ImgReg5IN_164,ImgReg5IN_163,ImgReg5IN_162,
                    ImgReg5IN_161,ImgReg5IN_160}), .CLK (nx23894), .RST (RST), .EN (
                    nx23770), .Q ({OutputImg5[175],OutputImg5[174],
                    OutputImg5[173],OutputImg5[172],OutputImg5[171],
                    OutputImg5[170],OutputImg5[169],OutputImg5[168],
                    OutputImg5[167],OutputImg5[166],OutputImg5[165],
                    OutputImg5[164],OutputImg5[163],OutputImg5[162],
                    OutputImg5[161],OutputImg5[160]})) ;
    triStateBuffer_16 loop3_11_TriState0L (.D ({OutputImg0[207],OutputImg0[206],
                      OutputImg0[205],OutputImg0[204],OutputImg0[203],
                      OutputImg0[202],OutputImg0[201],OutputImg0[200],
                      OutputImg0[199],OutputImg0[198],OutputImg0[197],
                      OutputImg0[196],OutputImg0[195],OutputImg0[194],
                      OutputImg0[193],OutputImg0[192]}), .EN (nx23684), .F ({
                      ImgReg0IN_191,ImgReg0IN_190,ImgReg0IN_189,ImgReg0IN_188,
                      ImgReg0IN_187,ImgReg0IN_186,ImgReg0IN_185,ImgReg0IN_184,
                      ImgReg0IN_183,ImgReg0IN_182,ImgReg0IN_181,ImgReg0IN_180,
                      ImgReg0IN_179,ImgReg0IN_178,ImgReg0IN_177,ImgReg0IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState1L (.D ({OutputImg1[207],OutputImg1[206],
                      OutputImg1[205],OutputImg1[204],OutputImg1[203],
                      OutputImg1[202],OutputImg1[201],OutputImg1[200],
                      OutputImg1[199],OutputImg1[198],OutputImg1[197],
                      OutputImg1[196],OutputImg1[195],OutputImg1[194],
                      OutputImg1[193],OutputImg1[192]}), .EN (nx23684), .F ({
                      ImgReg1IN_191,ImgReg1IN_190,ImgReg1IN_189,ImgReg1IN_188,
                      ImgReg1IN_187,ImgReg1IN_186,ImgReg1IN_185,ImgReg1IN_184,
                      ImgReg1IN_183,ImgReg1IN_182,ImgReg1IN_181,ImgReg1IN_180,
                      ImgReg1IN_179,ImgReg1IN_178,ImgReg1IN_177,ImgReg1IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState2L (.D ({OutputImg2[207],OutputImg2[206],
                      OutputImg2[205],OutputImg2[204],OutputImg2[203],
                      OutputImg2[202],OutputImg2[201],OutputImg2[200],
                      OutputImg2[199],OutputImg2[198],OutputImg2[197],
                      OutputImg2[196],OutputImg2[195],OutputImg2[194],
                      OutputImg2[193],OutputImg2[192]}), .EN (nx23684), .F ({
                      ImgReg2IN_191,ImgReg2IN_190,ImgReg2IN_189,ImgReg2IN_188,
                      ImgReg2IN_187,ImgReg2IN_186,ImgReg2IN_185,ImgReg2IN_184,
                      ImgReg2IN_183,ImgReg2IN_182,ImgReg2IN_181,ImgReg2IN_180,
                      ImgReg2IN_179,ImgReg2IN_178,ImgReg2IN_177,ImgReg2IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState3L (.D ({OutputImg3[207],OutputImg3[206],
                      OutputImg3[205],OutputImg3[204],OutputImg3[203],
                      OutputImg3[202],OutputImg3[201],OutputImg3[200],
                      OutputImg3[199],OutputImg3[198],OutputImg3[197],
                      OutputImg3[196],OutputImg3[195],OutputImg3[194],
                      OutputImg3[193],OutputImg3[192]}), .EN (nx23684), .F ({
                      ImgReg3IN_191,ImgReg3IN_190,ImgReg3IN_189,ImgReg3IN_188,
                      ImgReg3IN_187,ImgReg3IN_186,ImgReg3IN_185,ImgReg3IN_184,
                      ImgReg3IN_183,ImgReg3IN_182,ImgReg3IN_181,ImgReg3IN_180,
                      ImgReg3IN_179,ImgReg3IN_178,ImgReg3IN_177,ImgReg3IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState4L (.D ({OutputImg4[207],OutputImg4[206],
                      OutputImg4[205],OutputImg4[204],OutputImg4[203],
                      OutputImg4[202],OutputImg4[201],OutputImg4[200],
                      OutputImg4[199],OutputImg4[198],OutputImg4[197],
                      OutputImg4[196],OutputImg4[195],OutputImg4[194],
                      OutputImg4[193],OutputImg4[192]}), .EN (nx23686), .F ({
                      ImgReg4IN_191,ImgReg4IN_190,ImgReg4IN_189,ImgReg4IN_188,
                      ImgReg4IN_187,ImgReg4IN_186,ImgReg4IN_185,ImgReg4IN_184,
                      ImgReg4IN_183,ImgReg4IN_182,ImgReg4IN_181,ImgReg4IN_180,
                      ImgReg4IN_179,ImgReg4IN_178,ImgReg4IN_177,ImgReg4IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState5L (.D ({OutputImg5[207],OutputImg5[206],
                      OutputImg5[205],OutputImg5[204],OutputImg5[203],
                      OutputImg5[202],OutputImg5[201],OutputImg5[200],
                      OutputImg5[199],OutputImg5[198],OutputImg5[197],
                      OutputImg5[196],OutputImg5[195],OutputImg5[194],
                      OutputImg5[193],OutputImg5[192]}), .EN (nx23686), .F ({
                      ImgReg5IN_191,ImgReg5IN_190,ImgReg5IN_189,ImgReg5IN_188,
                      ImgReg5IN_187,ImgReg5IN_186,ImgReg5IN_185,ImgReg5IN_184,
                      ImgReg5IN_183,ImgReg5IN_182,ImgReg5IN_181,ImgReg5IN_180,
                      ImgReg5IN_179,ImgReg5IN_178,ImgReg5IN_177,ImgReg5IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState0N (.D ({DATA[191],DATA[190],DATA[189],
                      DATA[188],DATA[187],DATA[186],DATA[185],DATA[184],
                      DATA[183],DATA[182],DATA[181],DATA[180],DATA[179],
                      DATA[178],DATA[177],DATA[176]}), .EN (nx23656), .F ({
                      ImgReg0IN_191,ImgReg0IN_190,ImgReg0IN_189,ImgReg0IN_188,
                      ImgReg0IN_187,ImgReg0IN_186,ImgReg0IN_185,ImgReg0IN_184,
                      ImgReg0IN_183,ImgReg0IN_182,ImgReg0IN_181,ImgReg0IN_180,
                      ImgReg0IN_179,ImgReg0IN_178,ImgReg0IN_177,ImgReg0IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState1N (.D ({DATA[191],DATA[190],DATA[189],
                      DATA[188],DATA[187],DATA[186],DATA[185],DATA[184],
                      DATA[183],DATA[182],DATA[181],DATA[180],DATA[179],
                      DATA[178],DATA[177],DATA[176]}), .EN (nx23644), .F ({
                      ImgReg1IN_191,ImgReg1IN_190,ImgReg1IN_189,ImgReg1IN_188,
                      ImgReg1IN_187,ImgReg1IN_186,ImgReg1IN_185,ImgReg1IN_184,
                      ImgReg1IN_183,ImgReg1IN_182,ImgReg1IN_181,ImgReg1IN_180,
                      ImgReg1IN_179,ImgReg1IN_178,ImgReg1IN_177,ImgReg1IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState2N (.D ({DATA[191],DATA[190],DATA[189],
                      DATA[188],DATA[187],DATA[186],DATA[185],DATA[184],
                      DATA[183],DATA[182],DATA[181],DATA[180],DATA[179],
                      DATA[178],DATA[177],DATA[176]}), .EN (nx23632), .F ({
                      ImgReg2IN_191,ImgReg2IN_190,ImgReg2IN_189,ImgReg2IN_188,
                      ImgReg2IN_187,ImgReg2IN_186,ImgReg2IN_185,ImgReg2IN_184,
                      ImgReg2IN_183,ImgReg2IN_182,ImgReg2IN_181,ImgReg2IN_180,
                      ImgReg2IN_179,ImgReg2IN_178,ImgReg2IN_177,ImgReg2IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState3N (.D ({DATA[191],DATA[190],DATA[189],
                      DATA[188],DATA[187],DATA[186],DATA[185],DATA[184],
                      DATA[183],DATA[182],DATA[181],DATA[180],DATA[179],
                      DATA[178],DATA[177],DATA[176]}), .EN (nx23620), .F ({
                      ImgReg3IN_191,ImgReg3IN_190,ImgReg3IN_189,ImgReg3IN_188,
                      ImgReg3IN_187,ImgReg3IN_186,ImgReg3IN_185,ImgReg3IN_184,
                      ImgReg3IN_183,ImgReg3IN_182,ImgReg3IN_181,ImgReg3IN_180,
                      ImgReg3IN_179,ImgReg3IN_178,ImgReg3IN_177,ImgReg3IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState4N (.D ({DATA[191],DATA[190],DATA[189],
                      DATA[188],DATA[187],DATA[186],DATA[185],DATA[184],
                      DATA[183],DATA[182],DATA[181],DATA[180],DATA[179],
                      DATA[178],DATA[177],DATA[176]}), .EN (nx23608), .F ({
                      ImgReg4IN_191,ImgReg4IN_190,ImgReg4IN_189,ImgReg4IN_188,
                      ImgReg4IN_187,ImgReg4IN_186,ImgReg4IN_185,ImgReg4IN_184,
                      ImgReg4IN_183,ImgReg4IN_182,ImgReg4IN_181,ImgReg4IN_180,
                      ImgReg4IN_179,ImgReg4IN_178,ImgReg4IN_177,ImgReg4IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState5N (.D ({DATA[191],DATA[190],DATA[189],
                      DATA[188],DATA[187],DATA[186],DATA[185],DATA[184],
                      DATA[183],DATA[182],DATA[181],DATA[180],DATA[179],
                      DATA[178],DATA[177],DATA[176]}), .EN (nx23596), .F ({
                      ImgReg5IN_191,ImgReg5IN_190,ImgReg5IN_189,ImgReg5IN_188,
                      ImgReg5IN_187,ImgReg5IN_186,ImgReg5IN_185,ImgReg5IN_184,
                      ImgReg5IN_183,ImgReg5IN_182,ImgReg5IN_181,ImgReg5IN_180,
                      ImgReg5IN_179,ImgReg5IN_178,ImgReg5IN_177,ImgReg5IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState0U (.D ({OutputImg1[191],OutputImg1[190],
                      OutputImg1[189],OutputImg1[188],OutputImg1[187],
                      OutputImg1[186],OutputImg1[185],OutputImg1[184],
                      OutputImg1[183],OutputImg1[182],OutputImg1[181],
                      OutputImg1[180],OutputImg1[179],OutputImg1[178],
                      OutputImg1[177],OutputImg1[176]}), .EN (nx23800), .F ({
                      ImgReg0IN_191,ImgReg0IN_190,ImgReg0IN_189,ImgReg0IN_188,
                      ImgReg0IN_187,ImgReg0IN_186,ImgReg0IN_185,ImgReg0IN_184,
                      ImgReg0IN_183,ImgReg0IN_182,ImgReg0IN_181,ImgReg0IN_180,
                      ImgReg0IN_179,ImgReg0IN_178,ImgReg0IN_177,ImgReg0IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState1U (.D ({OutputImg2[191],OutputImg2[190],
                      OutputImg2[189],OutputImg2[188],OutputImg2[187],
                      OutputImg2[186],OutputImg2[185],OutputImg2[184],
                      OutputImg2[183],OutputImg2[182],OutputImg2[181],
                      OutputImg2[180],OutputImg2[179],OutputImg2[178],
                      OutputImg2[177],OutputImg2[176]}), .EN (nx23802), .F ({
                      ImgReg1IN_191,ImgReg1IN_190,ImgReg1IN_189,ImgReg1IN_188,
                      ImgReg1IN_187,ImgReg1IN_186,ImgReg1IN_185,ImgReg1IN_184,
                      ImgReg1IN_183,ImgReg1IN_182,ImgReg1IN_181,ImgReg1IN_180,
                      ImgReg1IN_179,ImgReg1IN_178,ImgReg1IN_177,ImgReg1IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState2U (.D ({OutputImg3[191],OutputImg3[190],
                      OutputImg3[189],OutputImg3[188],OutputImg3[187],
                      OutputImg3[186],OutputImg3[185],OutputImg3[184],
                      OutputImg3[183],OutputImg3[182],OutputImg3[181],
                      OutputImg3[180],OutputImg3[179],OutputImg3[178],
                      OutputImg3[177],OutputImg3[176]}), .EN (nx23802), .F ({
                      ImgReg2IN_191,ImgReg2IN_190,ImgReg2IN_189,ImgReg2IN_188,
                      ImgReg2IN_187,ImgReg2IN_186,ImgReg2IN_185,ImgReg2IN_184,
                      ImgReg2IN_183,ImgReg2IN_182,ImgReg2IN_181,ImgReg2IN_180,
                      ImgReg2IN_179,ImgReg2IN_178,ImgReg2IN_177,ImgReg2IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState3U (.D ({OutputImg4[191],OutputImg4[190],
                      OutputImg4[189],OutputImg4[188],OutputImg4[187],
                      OutputImg4[186],OutputImg4[185],OutputImg4[184],
                      OutputImg4[183],OutputImg4[182],OutputImg4[181],
                      OutputImg4[180],OutputImg4[179],OutputImg4[178],
                      OutputImg4[177],OutputImg4[176]}), .EN (nx23802), .F ({
                      ImgReg3IN_191,ImgReg3IN_190,ImgReg3IN_189,ImgReg3IN_188,
                      ImgReg3IN_187,ImgReg3IN_186,ImgReg3IN_185,ImgReg3IN_184,
                      ImgReg3IN_183,ImgReg3IN_182,ImgReg3IN_181,ImgReg3IN_180,
                      ImgReg3IN_179,ImgReg3IN_178,ImgReg3IN_177,ImgReg3IN_176})
                      ) ;
    triStateBuffer_16 loop3_11_TriState4U (.D ({OutputImg5[191],OutputImg5[190],
                      OutputImg5[189],OutputImg5[188],OutputImg5[187],
                      OutputImg5[186],OutputImg5[185],OutputImg5[184],
                      OutputImg5[183],OutputImg5[182],OutputImg5[181],
                      OutputImg5[180],OutputImg5[179],OutputImg5[178],
                      OutputImg5[177],OutputImg5[176]}), .EN (nx23802), .F ({
                      ImgReg4IN_191,ImgReg4IN_190,ImgReg4IN_189,ImgReg4IN_188,
                      ImgReg4IN_187,ImgReg4IN_186,ImgReg4IN_185,ImgReg4IN_184,
                      ImgReg4IN_183,ImgReg4IN_182,ImgReg4IN_181,ImgReg4IN_180,
                      ImgReg4IN_179,ImgReg4IN_178,ImgReg4IN_177,ImgReg4IN_176})
                      ) ;
    nBitRegister_16 loop3_11_reg1 (.D ({ImgReg0IN_191,ImgReg0IN_190,
                    ImgReg0IN_189,ImgReg0IN_188,ImgReg0IN_187,ImgReg0IN_186,
                    ImgReg0IN_185,ImgReg0IN_184,ImgReg0IN_183,ImgReg0IN_182,
                    ImgReg0IN_181,ImgReg0IN_180,ImgReg0IN_179,ImgReg0IN_178,
                    ImgReg0IN_177,ImgReg0IN_176}), .CLK (nx23894), .RST (RST), .EN (
                    nx23720), .Q ({OutputImg0[191],OutputImg0[190],
                    OutputImg0[189],OutputImg0[188],OutputImg0[187],
                    OutputImg0[186],OutputImg0[185],OutputImg0[184],
                    OutputImg0[183],OutputImg0[182],OutputImg0[181],
                    OutputImg0[180],OutputImg0[179],OutputImg0[178],
                    OutputImg0[177],OutputImg0[176]})) ;
    nBitRegister_16 loop3_11_reg2 (.D ({ImgReg1IN_191,ImgReg1IN_190,
                    ImgReg1IN_189,ImgReg1IN_188,ImgReg1IN_187,ImgReg1IN_186,
                    ImgReg1IN_185,ImgReg1IN_184,ImgReg1IN_183,ImgReg1IN_182,
                    ImgReg1IN_181,ImgReg1IN_180,ImgReg1IN_179,ImgReg1IN_178,
                    ImgReg1IN_177,ImgReg1IN_176}), .CLK (nx23896), .RST (RST), .EN (
                    nx23730), .Q ({OutputImg1[191],OutputImg1[190],
                    OutputImg1[189],OutputImg1[188],OutputImg1[187],
                    OutputImg1[186],OutputImg1[185],OutputImg1[184],
                    OutputImg1[183],OutputImg1[182],OutputImg1[181],
                    OutputImg1[180],OutputImg1[179],OutputImg1[178],
                    OutputImg1[177],OutputImg1[176]})) ;
    nBitRegister_16 loop3_11_reg3 (.D ({ImgReg2IN_191,ImgReg2IN_190,
                    ImgReg2IN_189,ImgReg2IN_188,ImgReg2IN_187,ImgReg2IN_186,
                    ImgReg2IN_185,ImgReg2IN_184,ImgReg2IN_183,ImgReg2IN_182,
                    ImgReg2IN_181,ImgReg2IN_180,ImgReg2IN_179,ImgReg2IN_178,
                    ImgReg2IN_177,ImgReg2IN_176}), .CLK (nx23896), .RST (RST), .EN (
                    nx23740), .Q ({OutputImg2[191],OutputImg2[190],
                    OutputImg2[189],OutputImg2[188],OutputImg2[187],
                    OutputImg2[186],OutputImg2[185],OutputImg2[184],
                    OutputImg2[183],OutputImg2[182],OutputImg2[181],
                    OutputImg2[180],OutputImg2[179],OutputImg2[178],
                    OutputImg2[177],OutputImg2[176]})) ;
    nBitRegister_16 loop3_11_reg4 (.D ({ImgReg3IN_191,ImgReg3IN_190,
                    ImgReg3IN_189,ImgReg3IN_188,ImgReg3IN_187,ImgReg3IN_186,
                    ImgReg3IN_185,ImgReg3IN_184,ImgReg3IN_183,ImgReg3IN_182,
                    ImgReg3IN_181,ImgReg3IN_180,ImgReg3IN_179,ImgReg3IN_178,
                    ImgReg3IN_177,ImgReg3IN_176}), .CLK (nx23898), .RST (RST), .EN (
                    nx23750), .Q ({OutputImg3[191],OutputImg3[190],
                    OutputImg3[189],OutputImg3[188],OutputImg3[187],
                    OutputImg3[186],OutputImg3[185],OutputImg3[184],
                    OutputImg3[183],OutputImg3[182],OutputImg3[181],
                    OutputImg3[180],OutputImg3[179],OutputImg3[178],
                    OutputImg3[177],OutputImg3[176]})) ;
    nBitRegister_16 loop3_11_reg5 (.D ({ImgReg4IN_191,ImgReg4IN_190,
                    ImgReg4IN_189,ImgReg4IN_188,ImgReg4IN_187,ImgReg4IN_186,
                    ImgReg4IN_185,ImgReg4IN_184,ImgReg4IN_183,ImgReg4IN_182,
                    ImgReg4IN_181,ImgReg4IN_180,ImgReg4IN_179,ImgReg4IN_178,
                    ImgReg4IN_177,ImgReg4IN_176}), .CLK (nx23898), .RST (RST), .EN (
                    nx23760), .Q ({OutputImg4[191],OutputImg4[190],
                    OutputImg4[189],OutputImg4[188],OutputImg4[187],
                    OutputImg4[186],OutputImg4[185],OutputImg4[184],
                    OutputImg4[183],OutputImg4[182],OutputImg4[181],
                    OutputImg4[180],OutputImg4[179],OutputImg4[178],
                    OutputImg4[177],OutputImg4[176]})) ;
    nBitRegister_16 loop3_11_reg6 (.D ({ImgReg5IN_191,ImgReg5IN_190,
                    ImgReg5IN_189,ImgReg5IN_188,ImgReg5IN_187,ImgReg5IN_186,
                    ImgReg5IN_185,ImgReg5IN_184,ImgReg5IN_183,ImgReg5IN_182,
                    ImgReg5IN_181,ImgReg5IN_180,ImgReg5IN_179,ImgReg5IN_178,
                    ImgReg5IN_177,ImgReg5IN_176}), .CLK (nx23900), .RST (RST), .EN (
                    nx23770), .Q ({OutputImg5[191],OutputImg5[190],
                    OutputImg5[189],OutputImg5[188],OutputImg5[187],
                    OutputImg5[186],OutputImg5[185],OutputImg5[184],
                    OutputImg5[183],OutputImg5[182],OutputImg5[181],
                    OutputImg5[180],OutputImg5[179],OutputImg5[178],
                    OutputImg5[177],OutputImg5[176]})) ;
    triStateBuffer_16 loop3_12_TriState0L (.D ({OutputImg0[223],OutputImg0[222],
                      OutputImg0[221],OutputImg0[220],OutputImg0[219],
                      OutputImg0[218],OutputImg0[217],OutputImg0[216],
                      OutputImg0[215],OutputImg0[214],OutputImg0[213],
                      OutputImg0[212],OutputImg0[211],OutputImg0[210],
                      OutputImg0[209],OutputImg0[208]}), .EN (nx23686), .F ({
                      ImgReg0IN_207,ImgReg0IN_206,ImgReg0IN_205,ImgReg0IN_204,
                      ImgReg0IN_203,ImgReg0IN_202,ImgReg0IN_201,ImgReg0IN_200,
                      ImgReg0IN_199,ImgReg0IN_198,ImgReg0IN_197,ImgReg0IN_196,
                      ImgReg0IN_195,ImgReg0IN_194,ImgReg0IN_193,ImgReg0IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState1L (.D ({OutputImg1[223],OutputImg1[222],
                      OutputImg1[221],OutputImg1[220],OutputImg1[219],
                      OutputImg1[218],OutputImg1[217],OutputImg1[216],
                      OutputImg1[215],OutputImg1[214],OutputImg1[213],
                      OutputImg1[212],OutputImg1[211],OutputImg1[210],
                      OutputImg1[209],OutputImg1[208]}), .EN (nx23686), .F ({
                      ImgReg1IN_207,ImgReg1IN_206,ImgReg1IN_205,ImgReg1IN_204,
                      ImgReg1IN_203,ImgReg1IN_202,ImgReg1IN_201,ImgReg1IN_200,
                      ImgReg1IN_199,ImgReg1IN_198,ImgReg1IN_197,ImgReg1IN_196,
                      ImgReg1IN_195,ImgReg1IN_194,ImgReg1IN_193,ImgReg1IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState2L (.D ({OutputImg2[223],OutputImg2[222],
                      OutputImg2[221],OutputImg2[220],OutputImg2[219],
                      OutputImg2[218],OutputImg2[217],OutputImg2[216],
                      OutputImg2[215],OutputImg2[214],OutputImg2[213],
                      OutputImg2[212],OutputImg2[211],OutputImg2[210],
                      OutputImg2[209],OutputImg2[208]}), .EN (nx23686), .F ({
                      ImgReg2IN_207,ImgReg2IN_206,ImgReg2IN_205,ImgReg2IN_204,
                      ImgReg2IN_203,ImgReg2IN_202,ImgReg2IN_201,ImgReg2IN_200,
                      ImgReg2IN_199,ImgReg2IN_198,ImgReg2IN_197,ImgReg2IN_196,
                      ImgReg2IN_195,ImgReg2IN_194,ImgReg2IN_193,ImgReg2IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState3L (.D ({OutputImg3[223],OutputImg3[222],
                      OutputImg3[221],OutputImg3[220],OutputImg3[219],
                      OutputImg3[218],OutputImg3[217],OutputImg3[216],
                      OutputImg3[215],OutputImg3[214],OutputImg3[213],
                      OutputImg3[212],OutputImg3[211],OutputImg3[210],
                      OutputImg3[209],OutputImg3[208]}), .EN (nx23686), .F ({
                      ImgReg3IN_207,ImgReg3IN_206,ImgReg3IN_205,ImgReg3IN_204,
                      ImgReg3IN_203,ImgReg3IN_202,ImgReg3IN_201,ImgReg3IN_200,
                      ImgReg3IN_199,ImgReg3IN_198,ImgReg3IN_197,ImgReg3IN_196,
                      ImgReg3IN_195,ImgReg3IN_194,ImgReg3IN_193,ImgReg3IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState4L (.D ({OutputImg4[223],OutputImg4[222],
                      OutputImg4[221],OutputImg4[220],OutputImg4[219],
                      OutputImg4[218],OutputImg4[217],OutputImg4[216],
                      OutputImg4[215],OutputImg4[214],OutputImg4[213],
                      OutputImg4[212],OutputImg4[211],OutputImg4[210],
                      OutputImg4[209],OutputImg4[208]}), .EN (nx23686), .F ({
                      ImgReg4IN_207,ImgReg4IN_206,ImgReg4IN_205,ImgReg4IN_204,
                      ImgReg4IN_203,ImgReg4IN_202,ImgReg4IN_201,ImgReg4IN_200,
                      ImgReg4IN_199,ImgReg4IN_198,ImgReg4IN_197,ImgReg4IN_196,
                      ImgReg4IN_195,ImgReg4IN_194,ImgReg4IN_193,ImgReg4IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState5L (.D ({OutputImg5[223],OutputImg5[222],
                      OutputImg5[221],OutputImg5[220],OutputImg5[219],
                      OutputImg5[218],OutputImg5[217],OutputImg5[216],
                      OutputImg5[215],OutputImg5[214],OutputImg5[213],
                      OutputImg5[212],OutputImg5[211],OutputImg5[210],
                      OutputImg5[209],OutputImg5[208]}), .EN (nx23688), .F ({
                      ImgReg5IN_207,ImgReg5IN_206,ImgReg5IN_205,ImgReg5IN_204,
                      ImgReg5IN_203,ImgReg5IN_202,ImgReg5IN_201,ImgReg5IN_200,
                      ImgReg5IN_199,ImgReg5IN_198,ImgReg5IN_197,ImgReg5IN_196,
                      ImgReg5IN_195,ImgReg5IN_194,ImgReg5IN_193,ImgReg5IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState0N (.D ({DATA[207],DATA[206],DATA[205],
                      DATA[204],DATA[203],DATA[202],DATA[201],DATA[200],
                      DATA[199],DATA[198],DATA[197],DATA[196],DATA[195],
                      DATA[194],DATA[193],DATA[192]}), .EN (nx23656), .F ({
                      ImgReg0IN_207,ImgReg0IN_206,ImgReg0IN_205,ImgReg0IN_204,
                      ImgReg0IN_203,ImgReg0IN_202,ImgReg0IN_201,ImgReg0IN_200,
                      ImgReg0IN_199,ImgReg0IN_198,ImgReg0IN_197,ImgReg0IN_196,
                      ImgReg0IN_195,ImgReg0IN_194,ImgReg0IN_193,ImgReg0IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState1N (.D ({DATA[207],DATA[206],DATA[205],
                      DATA[204],DATA[203],DATA[202],DATA[201],DATA[200],
                      DATA[199],DATA[198],DATA[197],DATA[196],DATA[195],
                      DATA[194],DATA[193],DATA[192]}), .EN (nx23644), .F ({
                      ImgReg1IN_207,ImgReg1IN_206,ImgReg1IN_205,ImgReg1IN_204,
                      ImgReg1IN_203,ImgReg1IN_202,ImgReg1IN_201,ImgReg1IN_200,
                      ImgReg1IN_199,ImgReg1IN_198,ImgReg1IN_197,ImgReg1IN_196,
                      ImgReg1IN_195,ImgReg1IN_194,ImgReg1IN_193,ImgReg1IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState2N (.D ({DATA[207],DATA[206],DATA[205],
                      DATA[204],DATA[203],DATA[202],DATA[201],DATA[200],
                      DATA[199],DATA[198],DATA[197],DATA[196],DATA[195],
                      DATA[194],DATA[193],DATA[192]}), .EN (nx23632), .F ({
                      ImgReg2IN_207,ImgReg2IN_206,ImgReg2IN_205,ImgReg2IN_204,
                      ImgReg2IN_203,ImgReg2IN_202,ImgReg2IN_201,ImgReg2IN_200,
                      ImgReg2IN_199,ImgReg2IN_198,ImgReg2IN_197,ImgReg2IN_196,
                      ImgReg2IN_195,ImgReg2IN_194,ImgReg2IN_193,ImgReg2IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState3N (.D ({DATA[207],DATA[206],DATA[205],
                      DATA[204],DATA[203],DATA[202],DATA[201],DATA[200],
                      DATA[199],DATA[198],DATA[197],DATA[196],DATA[195],
                      DATA[194],DATA[193],DATA[192]}), .EN (nx23620), .F ({
                      ImgReg3IN_207,ImgReg3IN_206,ImgReg3IN_205,ImgReg3IN_204,
                      ImgReg3IN_203,ImgReg3IN_202,ImgReg3IN_201,ImgReg3IN_200,
                      ImgReg3IN_199,ImgReg3IN_198,ImgReg3IN_197,ImgReg3IN_196,
                      ImgReg3IN_195,ImgReg3IN_194,ImgReg3IN_193,ImgReg3IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState4N (.D ({DATA[207],DATA[206],DATA[205],
                      DATA[204],DATA[203],DATA[202],DATA[201],DATA[200],
                      DATA[199],DATA[198],DATA[197],DATA[196],DATA[195],
                      DATA[194],DATA[193],DATA[192]}), .EN (nx23608), .F ({
                      ImgReg4IN_207,ImgReg4IN_206,ImgReg4IN_205,ImgReg4IN_204,
                      ImgReg4IN_203,ImgReg4IN_202,ImgReg4IN_201,ImgReg4IN_200,
                      ImgReg4IN_199,ImgReg4IN_198,ImgReg4IN_197,ImgReg4IN_196,
                      ImgReg4IN_195,ImgReg4IN_194,ImgReg4IN_193,ImgReg4IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState5N (.D ({DATA[207],DATA[206],DATA[205],
                      DATA[204],DATA[203],DATA[202],DATA[201],DATA[200],
                      DATA[199],DATA[198],DATA[197],DATA[196],DATA[195],
                      DATA[194],DATA[193],DATA[192]}), .EN (nx23596), .F ({
                      ImgReg5IN_207,ImgReg5IN_206,ImgReg5IN_205,ImgReg5IN_204,
                      ImgReg5IN_203,ImgReg5IN_202,ImgReg5IN_201,ImgReg5IN_200,
                      ImgReg5IN_199,ImgReg5IN_198,ImgReg5IN_197,ImgReg5IN_196,
                      ImgReg5IN_195,ImgReg5IN_194,ImgReg5IN_193,ImgReg5IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState0U (.D ({OutputImg1[207],OutputImg1[206],
                      OutputImg1[205],OutputImg1[204],OutputImg1[203],
                      OutputImg1[202],OutputImg1[201],OutputImg1[200],
                      OutputImg1[199],OutputImg1[198],OutputImg1[197],
                      OutputImg1[196],OutputImg1[195],OutputImg1[194],
                      OutputImg1[193],OutputImg1[192]}), .EN (nx23802), .F ({
                      ImgReg0IN_207,ImgReg0IN_206,ImgReg0IN_205,ImgReg0IN_204,
                      ImgReg0IN_203,ImgReg0IN_202,ImgReg0IN_201,ImgReg0IN_200,
                      ImgReg0IN_199,ImgReg0IN_198,ImgReg0IN_197,ImgReg0IN_196,
                      ImgReg0IN_195,ImgReg0IN_194,ImgReg0IN_193,ImgReg0IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState1U (.D ({OutputImg2[207],OutputImg2[206],
                      OutputImg2[205],OutputImg2[204],OutputImg2[203],
                      OutputImg2[202],OutputImg2[201],OutputImg2[200],
                      OutputImg2[199],OutputImg2[198],OutputImg2[197],
                      OutputImg2[196],OutputImg2[195],OutputImg2[194],
                      OutputImg2[193],OutputImg2[192]}), .EN (nx23802), .F ({
                      ImgReg1IN_207,ImgReg1IN_206,ImgReg1IN_205,ImgReg1IN_204,
                      ImgReg1IN_203,ImgReg1IN_202,ImgReg1IN_201,ImgReg1IN_200,
                      ImgReg1IN_199,ImgReg1IN_198,ImgReg1IN_197,ImgReg1IN_196,
                      ImgReg1IN_195,ImgReg1IN_194,ImgReg1IN_193,ImgReg1IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState2U (.D ({OutputImg3[207],OutputImg3[206],
                      OutputImg3[205],OutputImg3[204],OutputImg3[203],
                      OutputImg3[202],OutputImg3[201],OutputImg3[200],
                      OutputImg3[199],OutputImg3[198],OutputImg3[197],
                      OutputImg3[196],OutputImg3[195],OutputImg3[194],
                      OutputImg3[193],OutputImg3[192]}), .EN (nx23802), .F ({
                      ImgReg2IN_207,ImgReg2IN_206,ImgReg2IN_205,ImgReg2IN_204,
                      ImgReg2IN_203,ImgReg2IN_202,ImgReg2IN_201,ImgReg2IN_200,
                      ImgReg2IN_199,ImgReg2IN_198,ImgReg2IN_197,ImgReg2IN_196,
                      ImgReg2IN_195,ImgReg2IN_194,ImgReg2IN_193,ImgReg2IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState3U (.D ({OutputImg4[207],OutputImg4[206],
                      OutputImg4[205],OutputImg4[204],OutputImg4[203],
                      OutputImg4[202],OutputImg4[201],OutputImg4[200],
                      OutputImg4[199],OutputImg4[198],OutputImg4[197],
                      OutputImg4[196],OutputImg4[195],OutputImg4[194],
                      OutputImg4[193],OutputImg4[192]}), .EN (nx23804), .F ({
                      ImgReg3IN_207,ImgReg3IN_206,ImgReg3IN_205,ImgReg3IN_204,
                      ImgReg3IN_203,ImgReg3IN_202,ImgReg3IN_201,ImgReg3IN_200,
                      ImgReg3IN_199,ImgReg3IN_198,ImgReg3IN_197,ImgReg3IN_196,
                      ImgReg3IN_195,ImgReg3IN_194,ImgReg3IN_193,ImgReg3IN_192})
                      ) ;
    triStateBuffer_16 loop3_12_TriState4U (.D ({OutputImg5[207],OutputImg5[206],
                      OutputImg5[205],OutputImg5[204],OutputImg5[203],
                      OutputImg5[202],OutputImg5[201],OutputImg5[200],
                      OutputImg5[199],OutputImg5[198],OutputImg5[197],
                      OutputImg5[196],OutputImg5[195],OutputImg5[194],
                      OutputImg5[193],OutputImg5[192]}), .EN (nx23804), .F ({
                      ImgReg4IN_207,ImgReg4IN_206,ImgReg4IN_205,ImgReg4IN_204,
                      ImgReg4IN_203,ImgReg4IN_202,ImgReg4IN_201,ImgReg4IN_200,
                      ImgReg4IN_199,ImgReg4IN_198,ImgReg4IN_197,ImgReg4IN_196,
                      ImgReg4IN_195,ImgReg4IN_194,ImgReg4IN_193,ImgReg4IN_192})
                      ) ;
    nBitRegister_16 loop3_12_reg1 (.D ({ImgReg0IN_207,ImgReg0IN_206,
                    ImgReg0IN_205,ImgReg0IN_204,ImgReg0IN_203,ImgReg0IN_202,
                    ImgReg0IN_201,ImgReg0IN_200,ImgReg0IN_199,ImgReg0IN_198,
                    ImgReg0IN_197,ImgReg0IN_196,ImgReg0IN_195,ImgReg0IN_194,
                    ImgReg0IN_193,ImgReg0IN_192}), .CLK (nx23900), .RST (RST), .EN (
                    nx23720), .Q ({OutputImg0[207],OutputImg0[206],
                    OutputImg0[205],OutputImg0[204],OutputImg0[203],
                    OutputImg0[202],OutputImg0[201],OutputImg0[200],
                    OutputImg0[199],OutputImg0[198],OutputImg0[197],
                    OutputImg0[196],OutputImg0[195],OutputImg0[194],
                    OutputImg0[193],OutputImg0[192]})) ;
    nBitRegister_16 loop3_12_reg2 (.D ({ImgReg1IN_207,ImgReg1IN_206,
                    ImgReg1IN_205,ImgReg1IN_204,ImgReg1IN_203,ImgReg1IN_202,
                    ImgReg1IN_201,ImgReg1IN_200,ImgReg1IN_199,ImgReg1IN_198,
                    ImgReg1IN_197,ImgReg1IN_196,ImgReg1IN_195,ImgReg1IN_194,
                    ImgReg1IN_193,ImgReg1IN_192}), .CLK (nx23902), .RST (RST), .EN (
                    nx23730), .Q ({OutputImg1[207],OutputImg1[206],
                    OutputImg1[205],OutputImg1[204],OutputImg1[203],
                    OutputImg1[202],OutputImg1[201],OutputImg1[200],
                    OutputImg1[199],OutputImg1[198],OutputImg1[197],
                    OutputImg1[196],OutputImg1[195],OutputImg1[194],
                    OutputImg1[193],OutputImg1[192]})) ;
    nBitRegister_16 loop3_12_reg3 (.D ({ImgReg2IN_207,ImgReg2IN_206,
                    ImgReg2IN_205,ImgReg2IN_204,ImgReg2IN_203,ImgReg2IN_202,
                    ImgReg2IN_201,ImgReg2IN_200,ImgReg2IN_199,ImgReg2IN_198,
                    ImgReg2IN_197,ImgReg2IN_196,ImgReg2IN_195,ImgReg2IN_194,
                    ImgReg2IN_193,ImgReg2IN_192}), .CLK (nx23902), .RST (RST), .EN (
                    nx23740), .Q ({OutputImg2[207],OutputImg2[206],
                    OutputImg2[205],OutputImg2[204],OutputImg2[203],
                    OutputImg2[202],OutputImg2[201],OutputImg2[200],
                    OutputImg2[199],OutputImg2[198],OutputImg2[197],
                    OutputImg2[196],OutputImg2[195],OutputImg2[194],
                    OutputImg2[193],OutputImg2[192]})) ;
    nBitRegister_16 loop3_12_reg4 (.D ({ImgReg3IN_207,ImgReg3IN_206,
                    ImgReg3IN_205,ImgReg3IN_204,ImgReg3IN_203,ImgReg3IN_202,
                    ImgReg3IN_201,ImgReg3IN_200,ImgReg3IN_199,ImgReg3IN_198,
                    ImgReg3IN_197,ImgReg3IN_196,ImgReg3IN_195,ImgReg3IN_194,
                    ImgReg3IN_193,ImgReg3IN_192}), .CLK (nx23904), .RST (RST), .EN (
                    nx23750), .Q ({OutputImg3[207],OutputImg3[206],
                    OutputImg3[205],OutputImg3[204],OutputImg3[203],
                    OutputImg3[202],OutputImg3[201],OutputImg3[200],
                    OutputImg3[199],OutputImg3[198],OutputImg3[197],
                    OutputImg3[196],OutputImg3[195],OutputImg3[194],
                    OutputImg3[193],OutputImg3[192]})) ;
    nBitRegister_16 loop3_12_reg5 (.D ({ImgReg4IN_207,ImgReg4IN_206,
                    ImgReg4IN_205,ImgReg4IN_204,ImgReg4IN_203,ImgReg4IN_202,
                    ImgReg4IN_201,ImgReg4IN_200,ImgReg4IN_199,ImgReg4IN_198,
                    ImgReg4IN_197,ImgReg4IN_196,ImgReg4IN_195,ImgReg4IN_194,
                    ImgReg4IN_193,ImgReg4IN_192}), .CLK (nx23904), .RST (RST), .EN (
                    nx23760), .Q ({OutputImg4[207],OutputImg4[206],
                    OutputImg4[205],OutputImg4[204],OutputImg4[203],
                    OutputImg4[202],OutputImg4[201],OutputImg4[200],
                    OutputImg4[199],OutputImg4[198],OutputImg4[197],
                    OutputImg4[196],OutputImg4[195],OutputImg4[194],
                    OutputImg4[193],OutputImg4[192]})) ;
    nBitRegister_16 loop3_12_reg6 (.D ({ImgReg5IN_207,ImgReg5IN_206,
                    ImgReg5IN_205,ImgReg5IN_204,ImgReg5IN_203,ImgReg5IN_202,
                    ImgReg5IN_201,ImgReg5IN_200,ImgReg5IN_199,ImgReg5IN_198,
                    ImgReg5IN_197,ImgReg5IN_196,ImgReg5IN_195,ImgReg5IN_194,
                    ImgReg5IN_193,ImgReg5IN_192}), .CLK (nx23906), .RST (RST), .EN (
                    nx23770), .Q ({OutputImg5[207],OutputImg5[206],
                    OutputImg5[205],OutputImg5[204],OutputImg5[203],
                    OutputImg5[202],OutputImg5[201],OutputImg5[200],
                    OutputImg5[199],OutputImg5[198],OutputImg5[197],
                    OutputImg5[196],OutputImg5[195],OutputImg5[194],
                    OutputImg5[193],OutputImg5[192]})) ;
    triStateBuffer_16 loop3_13_TriState0L (.D ({OutputImg0[239],OutputImg0[238],
                      OutputImg0[237],OutputImg0[236],OutputImg0[235],
                      OutputImg0[234],OutputImg0[233],OutputImg0[232],
                      OutputImg0[231],OutputImg0[230],OutputImg0[229],
                      OutputImg0[228],OutputImg0[227],OutputImg0[226],
                      OutputImg0[225],OutputImg0[224]}), .EN (nx23688), .F ({
                      ImgReg0IN_223,ImgReg0IN_222,ImgReg0IN_221,ImgReg0IN_220,
                      ImgReg0IN_219,ImgReg0IN_218,ImgReg0IN_217,ImgReg0IN_216,
                      ImgReg0IN_215,ImgReg0IN_214,ImgReg0IN_213,ImgReg0IN_212,
                      ImgReg0IN_211,ImgReg0IN_210,ImgReg0IN_209,ImgReg0IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState1L (.D ({OutputImg1[239],OutputImg1[238],
                      OutputImg1[237],OutputImg1[236],OutputImg1[235],
                      OutputImg1[234],OutputImg1[233],OutputImg1[232],
                      OutputImg1[231],OutputImg1[230],OutputImg1[229],
                      OutputImg1[228],OutputImg1[227],OutputImg1[226],
                      OutputImg1[225],OutputImg1[224]}), .EN (nx23688), .F ({
                      ImgReg1IN_223,ImgReg1IN_222,ImgReg1IN_221,ImgReg1IN_220,
                      ImgReg1IN_219,ImgReg1IN_218,ImgReg1IN_217,ImgReg1IN_216,
                      ImgReg1IN_215,ImgReg1IN_214,ImgReg1IN_213,ImgReg1IN_212,
                      ImgReg1IN_211,ImgReg1IN_210,ImgReg1IN_209,ImgReg1IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState2L (.D ({OutputImg2[239],OutputImg2[238],
                      OutputImg2[237],OutputImg2[236],OutputImg2[235],
                      OutputImg2[234],OutputImg2[233],OutputImg2[232],
                      OutputImg2[231],OutputImg2[230],OutputImg2[229],
                      OutputImg2[228],OutputImg2[227],OutputImg2[226],
                      OutputImg2[225],OutputImg2[224]}), .EN (nx23688), .F ({
                      ImgReg2IN_223,ImgReg2IN_222,ImgReg2IN_221,ImgReg2IN_220,
                      ImgReg2IN_219,ImgReg2IN_218,ImgReg2IN_217,ImgReg2IN_216,
                      ImgReg2IN_215,ImgReg2IN_214,ImgReg2IN_213,ImgReg2IN_212,
                      ImgReg2IN_211,ImgReg2IN_210,ImgReg2IN_209,ImgReg2IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState3L (.D ({OutputImg3[239],OutputImg3[238],
                      OutputImg3[237],OutputImg3[236],OutputImg3[235],
                      OutputImg3[234],OutputImg3[233],OutputImg3[232],
                      OutputImg3[231],OutputImg3[230],OutputImg3[229],
                      OutputImg3[228],OutputImg3[227],OutputImg3[226],
                      OutputImg3[225],OutputImg3[224]}), .EN (nx23688), .F ({
                      ImgReg3IN_223,ImgReg3IN_222,ImgReg3IN_221,ImgReg3IN_220,
                      ImgReg3IN_219,ImgReg3IN_218,ImgReg3IN_217,ImgReg3IN_216,
                      ImgReg3IN_215,ImgReg3IN_214,ImgReg3IN_213,ImgReg3IN_212,
                      ImgReg3IN_211,ImgReg3IN_210,ImgReg3IN_209,ImgReg3IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState4L (.D ({OutputImg4[239],OutputImg4[238],
                      OutputImg4[237],OutputImg4[236],OutputImg4[235],
                      OutputImg4[234],OutputImg4[233],OutputImg4[232],
                      OutputImg4[231],OutputImg4[230],OutputImg4[229],
                      OutputImg4[228],OutputImg4[227],OutputImg4[226],
                      OutputImg4[225],OutputImg4[224]}), .EN (nx23688), .F ({
                      ImgReg4IN_223,ImgReg4IN_222,ImgReg4IN_221,ImgReg4IN_220,
                      ImgReg4IN_219,ImgReg4IN_218,ImgReg4IN_217,ImgReg4IN_216,
                      ImgReg4IN_215,ImgReg4IN_214,ImgReg4IN_213,ImgReg4IN_212,
                      ImgReg4IN_211,ImgReg4IN_210,ImgReg4IN_209,ImgReg4IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState5L (.D ({OutputImg5[239],OutputImg5[238],
                      OutputImg5[237],OutputImg5[236],OutputImg5[235],
                      OutputImg5[234],OutputImg5[233],OutputImg5[232],
                      OutputImg5[231],OutputImg5[230],OutputImg5[229],
                      OutputImg5[228],OutputImg5[227],OutputImg5[226],
                      OutputImg5[225],OutputImg5[224]}), .EN (nx23688), .F ({
                      ImgReg5IN_223,ImgReg5IN_222,ImgReg5IN_221,ImgReg5IN_220,
                      ImgReg5IN_219,ImgReg5IN_218,ImgReg5IN_217,ImgReg5IN_216,
                      ImgReg5IN_215,ImgReg5IN_214,ImgReg5IN_213,ImgReg5IN_212,
                      ImgReg5IN_211,ImgReg5IN_210,ImgReg5IN_209,ImgReg5IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState0N (.D ({DATA[223],DATA[222],DATA[221],
                      DATA[220],DATA[219],DATA[218],DATA[217],DATA[216],
                      DATA[215],DATA[214],DATA[213],DATA[212],DATA[211],
                      DATA[210],DATA[209],DATA[208]}), .EN (nx23656), .F ({
                      ImgReg0IN_223,ImgReg0IN_222,ImgReg0IN_221,ImgReg0IN_220,
                      ImgReg0IN_219,ImgReg0IN_218,ImgReg0IN_217,ImgReg0IN_216,
                      ImgReg0IN_215,ImgReg0IN_214,ImgReg0IN_213,ImgReg0IN_212,
                      ImgReg0IN_211,ImgReg0IN_210,ImgReg0IN_209,ImgReg0IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState1N (.D ({DATA[223],DATA[222],DATA[221],
                      DATA[220],DATA[219],DATA[218],DATA[217],DATA[216],
                      DATA[215],DATA[214],DATA[213],DATA[212],DATA[211],
                      DATA[210],DATA[209],DATA[208]}), .EN (nx23644), .F ({
                      ImgReg1IN_223,ImgReg1IN_222,ImgReg1IN_221,ImgReg1IN_220,
                      ImgReg1IN_219,ImgReg1IN_218,ImgReg1IN_217,ImgReg1IN_216,
                      ImgReg1IN_215,ImgReg1IN_214,ImgReg1IN_213,ImgReg1IN_212,
                      ImgReg1IN_211,ImgReg1IN_210,ImgReg1IN_209,ImgReg1IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState2N (.D ({DATA[223],DATA[222],DATA[221],
                      DATA[220],DATA[219],DATA[218],DATA[217],DATA[216],
                      DATA[215],DATA[214],DATA[213],DATA[212],DATA[211],
                      DATA[210],DATA[209],DATA[208]}), .EN (nx23632), .F ({
                      ImgReg2IN_223,ImgReg2IN_222,ImgReg2IN_221,ImgReg2IN_220,
                      ImgReg2IN_219,ImgReg2IN_218,ImgReg2IN_217,ImgReg2IN_216,
                      ImgReg2IN_215,ImgReg2IN_214,ImgReg2IN_213,ImgReg2IN_212,
                      ImgReg2IN_211,ImgReg2IN_210,ImgReg2IN_209,ImgReg2IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState3N (.D ({DATA[223],DATA[222],DATA[221],
                      DATA[220],DATA[219],DATA[218],DATA[217],DATA[216],
                      DATA[215],DATA[214],DATA[213],DATA[212],DATA[211],
                      DATA[210],DATA[209],DATA[208]}), .EN (nx23620), .F ({
                      ImgReg3IN_223,ImgReg3IN_222,ImgReg3IN_221,ImgReg3IN_220,
                      ImgReg3IN_219,ImgReg3IN_218,ImgReg3IN_217,ImgReg3IN_216,
                      ImgReg3IN_215,ImgReg3IN_214,ImgReg3IN_213,ImgReg3IN_212,
                      ImgReg3IN_211,ImgReg3IN_210,ImgReg3IN_209,ImgReg3IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState4N (.D ({DATA[223],DATA[222],DATA[221],
                      DATA[220],DATA[219],DATA[218],DATA[217],DATA[216],
                      DATA[215],DATA[214],DATA[213],DATA[212],DATA[211],
                      DATA[210],DATA[209],DATA[208]}), .EN (nx23608), .F ({
                      ImgReg4IN_223,ImgReg4IN_222,ImgReg4IN_221,ImgReg4IN_220,
                      ImgReg4IN_219,ImgReg4IN_218,ImgReg4IN_217,ImgReg4IN_216,
                      ImgReg4IN_215,ImgReg4IN_214,ImgReg4IN_213,ImgReg4IN_212,
                      ImgReg4IN_211,ImgReg4IN_210,ImgReg4IN_209,ImgReg4IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState5N (.D ({DATA[223],DATA[222],DATA[221],
                      DATA[220],DATA[219],DATA[218],DATA[217],DATA[216],
                      DATA[215],DATA[214],DATA[213],DATA[212],DATA[211],
                      DATA[210],DATA[209],DATA[208]}), .EN (nx23596), .F ({
                      ImgReg5IN_223,ImgReg5IN_222,ImgReg5IN_221,ImgReg5IN_220,
                      ImgReg5IN_219,ImgReg5IN_218,ImgReg5IN_217,ImgReg5IN_216,
                      ImgReg5IN_215,ImgReg5IN_214,ImgReg5IN_213,ImgReg5IN_212,
                      ImgReg5IN_211,ImgReg5IN_210,ImgReg5IN_209,ImgReg5IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState0U (.D ({OutputImg1[223],OutputImg1[222],
                      OutputImg1[221],OutputImg1[220],OutputImg1[219],
                      OutputImg1[218],OutputImg1[217],OutputImg1[216],
                      OutputImg1[215],OutputImg1[214],OutputImg1[213],
                      OutputImg1[212],OutputImg1[211],OutputImg1[210],
                      OutputImg1[209],OutputImg1[208]}), .EN (nx23804), .F ({
                      ImgReg0IN_223,ImgReg0IN_222,ImgReg0IN_221,ImgReg0IN_220,
                      ImgReg0IN_219,ImgReg0IN_218,ImgReg0IN_217,ImgReg0IN_216,
                      ImgReg0IN_215,ImgReg0IN_214,ImgReg0IN_213,ImgReg0IN_212,
                      ImgReg0IN_211,ImgReg0IN_210,ImgReg0IN_209,ImgReg0IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState1U (.D ({OutputImg2[223],OutputImg2[222],
                      OutputImg2[221],OutputImg2[220],OutputImg2[219],
                      OutputImg2[218],OutputImg2[217],OutputImg2[216],
                      OutputImg2[215],OutputImg2[214],OutputImg2[213],
                      OutputImg2[212],OutputImg2[211],OutputImg2[210],
                      OutputImg2[209],OutputImg2[208]}), .EN (nx23804), .F ({
                      ImgReg1IN_223,ImgReg1IN_222,ImgReg1IN_221,ImgReg1IN_220,
                      ImgReg1IN_219,ImgReg1IN_218,ImgReg1IN_217,ImgReg1IN_216,
                      ImgReg1IN_215,ImgReg1IN_214,ImgReg1IN_213,ImgReg1IN_212,
                      ImgReg1IN_211,ImgReg1IN_210,ImgReg1IN_209,ImgReg1IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState2U (.D ({OutputImg3[223],OutputImg3[222],
                      OutputImg3[221],OutputImg3[220],OutputImg3[219],
                      OutputImg3[218],OutputImg3[217],OutputImg3[216],
                      OutputImg3[215],OutputImg3[214],OutputImg3[213],
                      OutputImg3[212],OutputImg3[211],OutputImg3[210],
                      OutputImg3[209],OutputImg3[208]}), .EN (nx23804), .F ({
                      ImgReg2IN_223,ImgReg2IN_222,ImgReg2IN_221,ImgReg2IN_220,
                      ImgReg2IN_219,ImgReg2IN_218,ImgReg2IN_217,ImgReg2IN_216,
                      ImgReg2IN_215,ImgReg2IN_214,ImgReg2IN_213,ImgReg2IN_212,
                      ImgReg2IN_211,ImgReg2IN_210,ImgReg2IN_209,ImgReg2IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState3U (.D ({OutputImg4[223],OutputImg4[222],
                      OutputImg4[221],OutputImg4[220],OutputImg4[219],
                      OutputImg4[218],OutputImg4[217],OutputImg4[216],
                      OutputImg4[215],OutputImg4[214],OutputImg4[213],
                      OutputImg4[212],OutputImg4[211],OutputImg4[210],
                      OutputImg4[209],OutputImg4[208]}), .EN (nx23804), .F ({
                      ImgReg3IN_223,ImgReg3IN_222,ImgReg3IN_221,ImgReg3IN_220,
                      ImgReg3IN_219,ImgReg3IN_218,ImgReg3IN_217,ImgReg3IN_216,
                      ImgReg3IN_215,ImgReg3IN_214,ImgReg3IN_213,ImgReg3IN_212,
                      ImgReg3IN_211,ImgReg3IN_210,ImgReg3IN_209,ImgReg3IN_208})
                      ) ;
    triStateBuffer_16 loop3_13_TriState4U (.D ({OutputImg5[223],OutputImg5[222],
                      OutputImg5[221],OutputImg5[220],OutputImg5[219],
                      OutputImg5[218],OutputImg5[217],OutputImg5[216],
                      OutputImg5[215],OutputImg5[214],OutputImg5[213],
                      OutputImg5[212],OutputImg5[211],OutputImg5[210],
                      OutputImg5[209],OutputImg5[208]}), .EN (nx23804), .F ({
                      ImgReg4IN_223,ImgReg4IN_222,ImgReg4IN_221,ImgReg4IN_220,
                      ImgReg4IN_219,ImgReg4IN_218,ImgReg4IN_217,ImgReg4IN_216,
                      ImgReg4IN_215,ImgReg4IN_214,ImgReg4IN_213,ImgReg4IN_212,
                      ImgReg4IN_211,ImgReg4IN_210,ImgReg4IN_209,ImgReg4IN_208})
                      ) ;
    nBitRegister_16 loop3_13_reg1 (.D ({ImgReg0IN_223,ImgReg0IN_222,
                    ImgReg0IN_221,ImgReg0IN_220,ImgReg0IN_219,ImgReg0IN_218,
                    ImgReg0IN_217,ImgReg0IN_216,ImgReg0IN_215,ImgReg0IN_214,
                    ImgReg0IN_213,ImgReg0IN_212,ImgReg0IN_211,ImgReg0IN_210,
                    ImgReg0IN_209,ImgReg0IN_208}), .CLK (nx23906), .RST (RST), .EN (
                    nx23720), .Q ({OutputImg0[223],OutputImg0[222],
                    OutputImg0[221],OutputImg0[220],OutputImg0[219],
                    OutputImg0[218],OutputImg0[217],OutputImg0[216],
                    OutputImg0[215],OutputImg0[214],OutputImg0[213],
                    OutputImg0[212],OutputImg0[211],OutputImg0[210],
                    OutputImg0[209],OutputImg0[208]})) ;
    nBitRegister_16 loop3_13_reg2 (.D ({ImgReg1IN_223,ImgReg1IN_222,
                    ImgReg1IN_221,ImgReg1IN_220,ImgReg1IN_219,ImgReg1IN_218,
                    ImgReg1IN_217,ImgReg1IN_216,ImgReg1IN_215,ImgReg1IN_214,
                    ImgReg1IN_213,ImgReg1IN_212,ImgReg1IN_211,ImgReg1IN_210,
                    ImgReg1IN_209,ImgReg1IN_208}), .CLK (nx23908), .RST (RST), .EN (
                    nx23730), .Q ({OutputImg1[223],OutputImg1[222],
                    OutputImg1[221],OutputImg1[220],OutputImg1[219],
                    OutputImg1[218],OutputImg1[217],OutputImg1[216],
                    OutputImg1[215],OutputImg1[214],OutputImg1[213],
                    OutputImg1[212],OutputImg1[211],OutputImg1[210],
                    OutputImg1[209],OutputImg1[208]})) ;
    nBitRegister_16 loop3_13_reg3 (.D ({ImgReg2IN_223,ImgReg2IN_222,
                    ImgReg2IN_221,ImgReg2IN_220,ImgReg2IN_219,ImgReg2IN_218,
                    ImgReg2IN_217,ImgReg2IN_216,ImgReg2IN_215,ImgReg2IN_214,
                    ImgReg2IN_213,ImgReg2IN_212,ImgReg2IN_211,ImgReg2IN_210,
                    ImgReg2IN_209,ImgReg2IN_208}), .CLK (nx23908), .RST (RST), .EN (
                    nx23740), .Q ({OutputImg2[223],OutputImg2[222],
                    OutputImg2[221],OutputImg2[220],OutputImg2[219],
                    OutputImg2[218],OutputImg2[217],OutputImg2[216],
                    OutputImg2[215],OutputImg2[214],OutputImg2[213],
                    OutputImg2[212],OutputImg2[211],OutputImg2[210],
                    OutputImg2[209],OutputImg2[208]})) ;
    nBitRegister_16 loop3_13_reg4 (.D ({ImgReg3IN_223,ImgReg3IN_222,
                    ImgReg3IN_221,ImgReg3IN_220,ImgReg3IN_219,ImgReg3IN_218,
                    ImgReg3IN_217,ImgReg3IN_216,ImgReg3IN_215,ImgReg3IN_214,
                    ImgReg3IN_213,ImgReg3IN_212,ImgReg3IN_211,ImgReg3IN_210,
                    ImgReg3IN_209,ImgReg3IN_208}), .CLK (nx23910), .RST (RST), .EN (
                    nx23750), .Q ({OutputImg3[223],OutputImg3[222],
                    OutputImg3[221],OutputImg3[220],OutputImg3[219],
                    OutputImg3[218],OutputImg3[217],OutputImg3[216],
                    OutputImg3[215],OutputImg3[214],OutputImg3[213],
                    OutputImg3[212],OutputImg3[211],OutputImg3[210],
                    OutputImg3[209],OutputImg3[208]})) ;
    nBitRegister_16 loop3_13_reg5 (.D ({ImgReg4IN_223,ImgReg4IN_222,
                    ImgReg4IN_221,ImgReg4IN_220,ImgReg4IN_219,ImgReg4IN_218,
                    ImgReg4IN_217,ImgReg4IN_216,ImgReg4IN_215,ImgReg4IN_214,
                    ImgReg4IN_213,ImgReg4IN_212,ImgReg4IN_211,ImgReg4IN_210,
                    ImgReg4IN_209,ImgReg4IN_208}), .CLK (nx23910), .RST (RST), .EN (
                    nx23760), .Q ({OutputImg4[223],OutputImg4[222],
                    OutputImg4[221],OutputImg4[220],OutputImg4[219],
                    OutputImg4[218],OutputImg4[217],OutputImg4[216],
                    OutputImg4[215],OutputImg4[214],OutputImg4[213],
                    OutputImg4[212],OutputImg4[211],OutputImg4[210],
                    OutputImg4[209],OutputImg4[208]})) ;
    nBitRegister_16 loop3_13_reg6 (.D ({ImgReg5IN_223,ImgReg5IN_222,
                    ImgReg5IN_221,ImgReg5IN_220,ImgReg5IN_219,ImgReg5IN_218,
                    ImgReg5IN_217,ImgReg5IN_216,ImgReg5IN_215,ImgReg5IN_214,
                    ImgReg5IN_213,ImgReg5IN_212,ImgReg5IN_211,ImgReg5IN_210,
                    ImgReg5IN_209,ImgReg5IN_208}), .CLK (nx23912), .RST (RST), .EN (
                    nx23770), .Q ({OutputImg5[223],OutputImg5[222],
                    OutputImg5[221],OutputImg5[220],OutputImg5[219],
                    OutputImg5[218],OutputImg5[217],OutputImg5[216],
                    OutputImg5[215],OutputImg5[214],OutputImg5[213],
                    OutputImg5[212],OutputImg5[211],OutputImg5[210],
                    OutputImg5[209],OutputImg5[208]})) ;
    triStateBuffer_16 loop3_14_TriState0L (.D ({OutputImg0[255],OutputImg0[254],
                      OutputImg0[253],OutputImg0[252],OutputImg0[251],
                      OutputImg0[250],OutputImg0[249],OutputImg0[248],
                      OutputImg0[247],OutputImg0[246],OutputImg0[245],
                      OutputImg0[244],OutputImg0[243],OutputImg0[242],
                      OutputImg0[241],OutputImg0[240]}), .EN (nx23690), .F ({
                      ImgReg0IN_239,ImgReg0IN_238,ImgReg0IN_237,ImgReg0IN_236,
                      ImgReg0IN_235,ImgReg0IN_234,ImgReg0IN_233,ImgReg0IN_232,
                      ImgReg0IN_231,ImgReg0IN_230,ImgReg0IN_229,ImgReg0IN_228,
                      ImgReg0IN_227,ImgReg0IN_226,ImgReg0IN_225,ImgReg0IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState1L (.D ({OutputImg1[255],OutputImg1[254],
                      OutputImg1[253],OutputImg1[252],OutputImg1[251],
                      OutputImg1[250],OutputImg1[249],OutputImg1[248],
                      OutputImg1[247],OutputImg1[246],OutputImg1[245],
                      OutputImg1[244],OutputImg1[243],OutputImg1[242],
                      OutputImg1[241],OutputImg1[240]}), .EN (nx23690), .F ({
                      ImgReg1IN_239,ImgReg1IN_238,ImgReg1IN_237,ImgReg1IN_236,
                      ImgReg1IN_235,ImgReg1IN_234,ImgReg1IN_233,ImgReg1IN_232,
                      ImgReg1IN_231,ImgReg1IN_230,ImgReg1IN_229,ImgReg1IN_228,
                      ImgReg1IN_227,ImgReg1IN_226,ImgReg1IN_225,ImgReg1IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState2L (.D ({OutputImg2[255],OutputImg2[254],
                      OutputImg2[253],OutputImg2[252],OutputImg2[251],
                      OutputImg2[250],OutputImg2[249],OutputImg2[248],
                      OutputImg2[247],OutputImg2[246],OutputImg2[245],
                      OutputImg2[244],OutputImg2[243],OutputImg2[242],
                      OutputImg2[241],OutputImg2[240]}), .EN (nx23690), .F ({
                      ImgReg2IN_239,ImgReg2IN_238,ImgReg2IN_237,ImgReg2IN_236,
                      ImgReg2IN_235,ImgReg2IN_234,ImgReg2IN_233,ImgReg2IN_232,
                      ImgReg2IN_231,ImgReg2IN_230,ImgReg2IN_229,ImgReg2IN_228,
                      ImgReg2IN_227,ImgReg2IN_226,ImgReg2IN_225,ImgReg2IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState3L (.D ({OutputImg3[255],OutputImg3[254],
                      OutputImg3[253],OutputImg3[252],OutputImg3[251],
                      OutputImg3[250],OutputImg3[249],OutputImg3[248],
                      OutputImg3[247],OutputImg3[246],OutputImg3[245],
                      OutputImg3[244],OutputImg3[243],OutputImg3[242],
                      OutputImg3[241],OutputImg3[240]}), .EN (nx23690), .F ({
                      ImgReg3IN_239,ImgReg3IN_238,ImgReg3IN_237,ImgReg3IN_236,
                      ImgReg3IN_235,ImgReg3IN_234,ImgReg3IN_233,ImgReg3IN_232,
                      ImgReg3IN_231,ImgReg3IN_230,ImgReg3IN_229,ImgReg3IN_228,
                      ImgReg3IN_227,ImgReg3IN_226,ImgReg3IN_225,ImgReg3IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState4L (.D ({OutputImg4[255],OutputImg4[254],
                      OutputImg4[253],OutputImg4[252],OutputImg4[251],
                      OutputImg4[250],OutputImg4[249],OutputImg4[248],
                      OutputImg4[247],OutputImg4[246],OutputImg4[245],
                      OutputImg4[244],OutputImg4[243],OutputImg4[242],
                      OutputImg4[241],OutputImg4[240]}), .EN (nx23690), .F ({
                      ImgReg4IN_239,ImgReg4IN_238,ImgReg4IN_237,ImgReg4IN_236,
                      ImgReg4IN_235,ImgReg4IN_234,ImgReg4IN_233,ImgReg4IN_232,
                      ImgReg4IN_231,ImgReg4IN_230,ImgReg4IN_229,ImgReg4IN_228,
                      ImgReg4IN_227,ImgReg4IN_226,ImgReg4IN_225,ImgReg4IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState5L (.D ({OutputImg5[255],OutputImg5[254],
                      OutputImg5[253],OutputImg5[252],OutputImg5[251],
                      OutputImg5[250],OutputImg5[249],OutputImg5[248],
                      OutputImg5[247],OutputImg5[246],OutputImg5[245],
                      OutputImg5[244],OutputImg5[243],OutputImg5[242],
                      OutputImg5[241],OutputImg5[240]}), .EN (nx23690), .F ({
                      ImgReg5IN_239,ImgReg5IN_238,ImgReg5IN_237,ImgReg5IN_236,
                      ImgReg5IN_235,ImgReg5IN_234,ImgReg5IN_233,ImgReg5IN_232,
                      ImgReg5IN_231,ImgReg5IN_230,ImgReg5IN_229,ImgReg5IN_228,
                      ImgReg5IN_227,ImgReg5IN_226,ImgReg5IN_225,ImgReg5IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState0N (.D ({DATA[239],DATA[238],DATA[237],
                      DATA[236],DATA[235],DATA[234],DATA[233],DATA[232],
                      DATA[231],DATA[230],DATA[229],DATA[228],DATA[227],
                      DATA[226],DATA[225],DATA[224]}), .EN (nx23658), .F ({
                      ImgReg0IN_239,ImgReg0IN_238,ImgReg0IN_237,ImgReg0IN_236,
                      ImgReg0IN_235,ImgReg0IN_234,ImgReg0IN_233,ImgReg0IN_232,
                      ImgReg0IN_231,ImgReg0IN_230,ImgReg0IN_229,ImgReg0IN_228,
                      ImgReg0IN_227,ImgReg0IN_226,ImgReg0IN_225,ImgReg0IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState1N (.D ({DATA[239],DATA[238],DATA[237],
                      DATA[236],DATA[235],DATA[234],DATA[233],DATA[232],
                      DATA[231],DATA[230],DATA[229],DATA[228],DATA[227],
                      DATA[226],DATA[225],DATA[224]}), .EN (nx23646), .F ({
                      ImgReg1IN_239,ImgReg1IN_238,ImgReg1IN_237,ImgReg1IN_236,
                      ImgReg1IN_235,ImgReg1IN_234,ImgReg1IN_233,ImgReg1IN_232,
                      ImgReg1IN_231,ImgReg1IN_230,ImgReg1IN_229,ImgReg1IN_228,
                      ImgReg1IN_227,ImgReg1IN_226,ImgReg1IN_225,ImgReg1IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState2N (.D ({DATA[239],DATA[238],DATA[237],
                      DATA[236],DATA[235],DATA[234],DATA[233],DATA[232],
                      DATA[231],DATA[230],DATA[229],DATA[228],DATA[227],
                      DATA[226],DATA[225],DATA[224]}), .EN (nx23634), .F ({
                      ImgReg2IN_239,ImgReg2IN_238,ImgReg2IN_237,ImgReg2IN_236,
                      ImgReg2IN_235,ImgReg2IN_234,ImgReg2IN_233,ImgReg2IN_232,
                      ImgReg2IN_231,ImgReg2IN_230,ImgReg2IN_229,ImgReg2IN_228,
                      ImgReg2IN_227,ImgReg2IN_226,ImgReg2IN_225,ImgReg2IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState3N (.D ({DATA[239],DATA[238],DATA[237],
                      DATA[236],DATA[235],DATA[234],DATA[233],DATA[232],
                      DATA[231],DATA[230],DATA[229],DATA[228],DATA[227],
                      DATA[226],DATA[225],DATA[224]}), .EN (nx23622), .F ({
                      ImgReg3IN_239,ImgReg3IN_238,ImgReg3IN_237,ImgReg3IN_236,
                      ImgReg3IN_235,ImgReg3IN_234,ImgReg3IN_233,ImgReg3IN_232,
                      ImgReg3IN_231,ImgReg3IN_230,ImgReg3IN_229,ImgReg3IN_228,
                      ImgReg3IN_227,ImgReg3IN_226,ImgReg3IN_225,ImgReg3IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState4N (.D ({DATA[239],DATA[238],DATA[237],
                      DATA[236],DATA[235],DATA[234],DATA[233],DATA[232],
                      DATA[231],DATA[230],DATA[229],DATA[228],DATA[227],
                      DATA[226],DATA[225],DATA[224]}), .EN (nx23610), .F ({
                      ImgReg4IN_239,ImgReg4IN_238,ImgReg4IN_237,ImgReg4IN_236,
                      ImgReg4IN_235,ImgReg4IN_234,ImgReg4IN_233,ImgReg4IN_232,
                      ImgReg4IN_231,ImgReg4IN_230,ImgReg4IN_229,ImgReg4IN_228,
                      ImgReg4IN_227,ImgReg4IN_226,ImgReg4IN_225,ImgReg4IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState5N (.D ({DATA[239],DATA[238],DATA[237],
                      DATA[236],DATA[235],DATA[234],DATA[233],DATA[232],
                      DATA[231],DATA[230],DATA[229],DATA[228],DATA[227],
                      DATA[226],DATA[225],DATA[224]}), .EN (nx23598), .F ({
                      ImgReg5IN_239,ImgReg5IN_238,ImgReg5IN_237,ImgReg5IN_236,
                      ImgReg5IN_235,ImgReg5IN_234,ImgReg5IN_233,ImgReg5IN_232,
                      ImgReg5IN_231,ImgReg5IN_230,ImgReg5IN_229,ImgReg5IN_228,
                      ImgReg5IN_227,ImgReg5IN_226,ImgReg5IN_225,ImgReg5IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState0U (.D ({OutputImg1[239],OutputImg1[238],
                      OutputImg1[237],OutputImg1[236],OutputImg1[235],
                      OutputImg1[234],OutputImg1[233],OutputImg1[232],
                      OutputImg1[231],OutputImg1[230],OutputImg1[229],
                      OutputImg1[228],OutputImg1[227],OutputImg1[226],
                      OutputImg1[225],OutputImg1[224]}), .EN (nx23806), .F ({
                      ImgReg0IN_239,ImgReg0IN_238,ImgReg0IN_237,ImgReg0IN_236,
                      ImgReg0IN_235,ImgReg0IN_234,ImgReg0IN_233,ImgReg0IN_232,
                      ImgReg0IN_231,ImgReg0IN_230,ImgReg0IN_229,ImgReg0IN_228,
                      ImgReg0IN_227,ImgReg0IN_226,ImgReg0IN_225,ImgReg0IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState1U (.D ({OutputImg2[239],OutputImg2[238],
                      OutputImg2[237],OutputImg2[236],OutputImg2[235],
                      OutputImg2[234],OutputImg2[233],OutputImg2[232],
                      OutputImg2[231],OutputImg2[230],OutputImg2[229],
                      OutputImg2[228],OutputImg2[227],OutputImg2[226],
                      OutputImg2[225],OutputImg2[224]}), .EN (nx23806), .F ({
                      ImgReg1IN_239,ImgReg1IN_238,ImgReg1IN_237,ImgReg1IN_236,
                      ImgReg1IN_235,ImgReg1IN_234,ImgReg1IN_233,ImgReg1IN_232,
                      ImgReg1IN_231,ImgReg1IN_230,ImgReg1IN_229,ImgReg1IN_228,
                      ImgReg1IN_227,ImgReg1IN_226,ImgReg1IN_225,ImgReg1IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState2U (.D ({OutputImg3[239],OutputImg3[238],
                      OutputImg3[237],OutputImg3[236],OutputImg3[235],
                      OutputImg3[234],OutputImg3[233],OutputImg3[232],
                      OutputImg3[231],OutputImg3[230],OutputImg3[229],
                      OutputImg3[228],OutputImg3[227],OutputImg3[226],
                      OutputImg3[225],OutputImg3[224]}), .EN (nx23806), .F ({
                      ImgReg2IN_239,ImgReg2IN_238,ImgReg2IN_237,ImgReg2IN_236,
                      ImgReg2IN_235,ImgReg2IN_234,ImgReg2IN_233,ImgReg2IN_232,
                      ImgReg2IN_231,ImgReg2IN_230,ImgReg2IN_229,ImgReg2IN_228,
                      ImgReg2IN_227,ImgReg2IN_226,ImgReg2IN_225,ImgReg2IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState3U (.D ({OutputImg4[239],OutputImg4[238],
                      OutputImg4[237],OutputImg4[236],OutputImg4[235],
                      OutputImg4[234],OutputImg4[233],OutputImg4[232],
                      OutputImg4[231],OutputImg4[230],OutputImg4[229],
                      OutputImg4[228],OutputImg4[227],OutputImg4[226],
                      OutputImg4[225],OutputImg4[224]}), .EN (nx23806), .F ({
                      ImgReg3IN_239,ImgReg3IN_238,ImgReg3IN_237,ImgReg3IN_236,
                      ImgReg3IN_235,ImgReg3IN_234,ImgReg3IN_233,ImgReg3IN_232,
                      ImgReg3IN_231,ImgReg3IN_230,ImgReg3IN_229,ImgReg3IN_228,
                      ImgReg3IN_227,ImgReg3IN_226,ImgReg3IN_225,ImgReg3IN_224})
                      ) ;
    triStateBuffer_16 loop3_14_TriState4U (.D ({OutputImg5[239],OutputImg5[238],
                      OutputImg5[237],OutputImg5[236],OutputImg5[235],
                      OutputImg5[234],OutputImg5[233],OutputImg5[232],
                      OutputImg5[231],OutputImg5[230],OutputImg5[229],
                      OutputImg5[228],OutputImg5[227],OutputImg5[226],
                      OutputImg5[225],OutputImg5[224]}), .EN (nx23806), .F ({
                      ImgReg4IN_239,ImgReg4IN_238,ImgReg4IN_237,ImgReg4IN_236,
                      ImgReg4IN_235,ImgReg4IN_234,ImgReg4IN_233,ImgReg4IN_232,
                      ImgReg4IN_231,ImgReg4IN_230,ImgReg4IN_229,ImgReg4IN_228,
                      ImgReg4IN_227,ImgReg4IN_226,ImgReg4IN_225,ImgReg4IN_224})
                      ) ;
    nBitRegister_16 loop3_14_reg1 (.D ({ImgReg0IN_239,ImgReg0IN_238,
                    ImgReg0IN_237,ImgReg0IN_236,ImgReg0IN_235,ImgReg0IN_234,
                    ImgReg0IN_233,ImgReg0IN_232,ImgReg0IN_231,ImgReg0IN_230,
                    ImgReg0IN_229,ImgReg0IN_228,ImgReg0IN_227,ImgReg0IN_226,
                    ImgReg0IN_225,ImgReg0IN_224}), .CLK (nx23912), .RST (RST), .EN (
                    nx23722), .Q ({OutputImg0[239],OutputImg0[238],
                    OutputImg0[237],OutputImg0[236],OutputImg0[235],
                    OutputImg0[234],OutputImg0[233],OutputImg0[232],
                    OutputImg0[231],OutputImg0[230],OutputImg0[229],
                    OutputImg0[228],OutputImg0[227],OutputImg0[226],
                    OutputImg0[225],OutputImg0[224]})) ;
    nBitRegister_16 loop3_14_reg2 (.D ({ImgReg1IN_239,ImgReg1IN_238,
                    ImgReg1IN_237,ImgReg1IN_236,ImgReg1IN_235,ImgReg1IN_234,
                    ImgReg1IN_233,ImgReg1IN_232,ImgReg1IN_231,ImgReg1IN_230,
                    ImgReg1IN_229,ImgReg1IN_228,ImgReg1IN_227,ImgReg1IN_226,
                    ImgReg1IN_225,ImgReg1IN_224}), .CLK (nx23914), .RST (RST), .EN (
                    nx23732), .Q ({OutputImg1[239],OutputImg1[238],
                    OutputImg1[237],OutputImg1[236],OutputImg1[235],
                    OutputImg1[234],OutputImg1[233],OutputImg1[232],
                    OutputImg1[231],OutputImg1[230],OutputImg1[229],
                    OutputImg1[228],OutputImg1[227],OutputImg1[226],
                    OutputImg1[225],OutputImg1[224]})) ;
    nBitRegister_16 loop3_14_reg3 (.D ({ImgReg2IN_239,ImgReg2IN_238,
                    ImgReg2IN_237,ImgReg2IN_236,ImgReg2IN_235,ImgReg2IN_234,
                    ImgReg2IN_233,ImgReg2IN_232,ImgReg2IN_231,ImgReg2IN_230,
                    ImgReg2IN_229,ImgReg2IN_228,ImgReg2IN_227,ImgReg2IN_226,
                    ImgReg2IN_225,ImgReg2IN_224}), .CLK (nx23914), .RST (RST), .EN (
                    nx23742), .Q ({OutputImg2[239],OutputImg2[238],
                    OutputImg2[237],OutputImg2[236],OutputImg2[235],
                    OutputImg2[234],OutputImg2[233],OutputImg2[232],
                    OutputImg2[231],OutputImg2[230],OutputImg2[229],
                    OutputImg2[228],OutputImg2[227],OutputImg2[226],
                    OutputImg2[225],OutputImg2[224]})) ;
    nBitRegister_16 loop3_14_reg4 (.D ({ImgReg3IN_239,ImgReg3IN_238,
                    ImgReg3IN_237,ImgReg3IN_236,ImgReg3IN_235,ImgReg3IN_234,
                    ImgReg3IN_233,ImgReg3IN_232,ImgReg3IN_231,ImgReg3IN_230,
                    ImgReg3IN_229,ImgReg3IN_228,ImgReg3IN_227,ImgReg3IN_226,
                    ImgReg3IN_225,ImgReg3IN_224}), .CLK (nx23916), .RST (RST), .EN (
                    nx23752), .Q ({OutputImg3[239],OutputImg3[238],
                    OutputImg3[237],OutputImg3[236],OutputImg3[235],
                    OutputImg3[234],OutputImg3[233],OutputImg3[232],
                    OutputImg3[231],OutputImg3[230],OutputImg3[229],
                    OutputImg3[228],OutputImg3[227],OutputImg3[226],
                    OutputImg3[225],OutputImg3[224]})) ;
    nBitRegister_16 loop3_14_reg5 (.D ({ImgReg4IN_239,ImgReg4IN_238,
                    ImgReg4IN_237,ImgReg4IN_236,ImgReg4IN_235,ImgReg4IN_234,
                    ImgReg4IN_233,ImgReg4IN_232,ImgReg4IN_231,ImgReg4IN_230,
                    ImgReg4IN_229,ImgReg4IN_228,ImgReg4IN_227,ImgReg4IN_226,
                    ImgReg4IN_225,ImgReg4IN_224}), .CLK (nx23916), .RST (RST), .EN (
                    nx23762), .Q ({OutputImg4[239],OutputImg4[238],
                    OutputImg4[237],OutputImg4[236],OutputImg4[235],
                    OutputImg4[234],OutputImg4[233],OutputImg4[232],
                    OutputImg4[231],OutputImg4[230],OutputImg4[229],
                    OutputImg4[228],OutputImg4[227],OutputImg4[226],
                    OutputImg4[225],OutputImg4[224]})) ;
    nBitRegister_16 loop3_14_reg6 (.D ({ImgReg5IN_239,ImgReg5IN_238,
                    ImgReg5IN_237,ImgReg5IN_236,ImgReg5IN_235,ImgReg5IN_234,
                    ImgReg5IN_233,ImgReg5IN_232,ImgReg5IN_231,ImgReg5IN_230,
                    ImgReg5IN_229,ImgReg5IN_228,ImgReg5IN_227,ImgReg5IN_226,
                    ImgReg5IN_225,ImgReg5IN_224}), .CLK (nx23918), .RST (RST), .EN (
                    nx23772), .Q ({OutputImg5[239],OutputImg5[238],
                    OutputImg5[237],OutputImg5[236],OutputImg5[235],
                    OutputImg5[234],OutputImg5[233],OutputImg5[232],
                    OutputImg5[231],OutputImg5[230],OutputImg5[229],
                    OutputImg5[228],OutputImg5[227],OutputImg5[226],
                    OutputImg5[225],OutputImg5[224]})) ;
    triStateBuffer_16 loop3_15_TriState0L (.D ({OutputImg0[271],OutputImg0[270],
                      OutputImg0[269],OutputImg0[268],OutputImg0[267],
                      OutputImg0[266],OutputImg0[265],OutputImg0[264],
                      OutputImg0[263],OutputImg0[262],OutputImg0[261],
                      OutputImg0[260],OutputImg0[259],OutputImg0[258],
                      OutputImg0[257],OutputImg0[256]}), .EN (nx23690), .F ({
                      ImgReg0IN_255,ImgReg0IN_254,ImgReg0IN_253,ImgReg0IN_252,
                      ImgReg0IN_251,ImgReg0IN_250,ImgReg0IN_249,ImgReg0IN_248,
                      ImgReg0IN_247,ImgReg0IN_246,ImgReg0IN_245,ImgReg0IN_244,
                      ImgReg0IN_243,ImgReg0IN_242,ImgReg0IN_241,ImgReg0IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState1L (.D ({OutputImg1[271],OutputImg1[270],
                      OutputImg1[269],OutputImg1[268],OutputImg1[267],
                      OutputImg1[266],OutputImg1[265],OutputImg1[264],
                      OutputImg1[263],OutputImg1[262],OutputImg1[261],
                      OutputImg1[260],OutputImg1[259],OutputImg1[258],
                      OutputImg1[257],OutputImg1[256]}), .EN (nx23692), .F ({
                      ImgReg1IN_255,ImgReg1IN_254,ImgReg1IN_253,ImgReg1IN_252,
                      ImgReg1IN_251,ImgReg1IN_250,ImgReg1IN_249,ImgReg1IN_248,
                      ImgReg1IN_247,ImgReg1IN_246,ImgReg1IN_245,ImgReg1IN_244,
                      ImgReg1IN_243,ImgReg1IN_242,ImgReg1IN_241,ImgReg1IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState2L (.D ({OutputImg2[271],OutputImg2[270],
                      OutputImg2[269],OutputImg2[268],OutputImg2[267],
                      OutputImg2[266],OutputImg2[265],OutputImg2[264],
                      OutputImg2[263],OutputImg2[262],OutputImg2[261],
                      OutputImg2[260],OutputImg2[259],OutputImg2[258],
                      OutputImg2[257],OutputImg2[256]}), .EN (nx23692), .F ({
                      ImgReg2IN_255,ImgReg2IN_254,ImgReg2IN_253,ImgReg2IN_252,
                      ImgReg2IN_251,ImgReg2IN_250,ImgReg2IN_249,ImgReg2IN_248,
                      ImgReg2IN_247,ImgReg2IN_246,ImgReg2IN_245,ImgReg2IN_244,
                      ImgReg2IN_243,ImgReg2IN_242,ImgReg2IN_241,ImgReg2IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState3L (.D ({OutputImg3[271],OutputImg3[270],
                      OutputImg3[269],OutputImg3[268],OutputImg3[267],
                      OutputImg3[266],OutputImg3[265],OutputImg3[264],
                      OutputImg3[263],OutputImg3[262],OutputImg3[261],
                      OutputImg3[260],OutputImg3[259],OutputImg3[258],
                      OutputImg3[257],OutputImg3[256]}), .EN (nx23692), .F ({
                      ImgReg3IN_255,ImgReg3IN_254,ImgReg3IN_253,ImgReg3IN_252,
                      ImgReg3IN_251,ImgReg3IN_250,ImgReg3IN_249,ImgReg3IN_248,
                      ImgReg3IN_247,ImgReg3IN_246,ImgReg3IN_245,ImgReg3IN_244,
                      ImgReg3IN_243,ImgReg3IN_242,ImgReg3IN_241,ImgReg3IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState4L (.D ({OutputImg4[271],OutputImg4[270],
                      OutputImg4[269],OutputImg4[268],OutputImg4[267],
                      OutputImg4[266],OutputImg4[265],OutputImg4[264],
                      OutputImg4[263],OutputImg4[262],OutputImg4[261],
                      OutputImg4[260],OutputImg4[259],OutputImg4[258],
                      OutputImg4[257],OutputImg4[256]}), .EN (nx23692), .F ({
                      ImgReg4IN_255,ImgReg4IN_254,ImgReg4IN_253,ImgReg4IN_252,
                      ImgReg4IN_251,ImgReg4IN_250,ImgReg4IN_249,ImgReg4IN_248,
                      ImgReg4IN_247,ImgReg4IN_246,ImgReg4IN_245,ImgReg4IN_244,
                      ImgReg4IN_243,ImgReg4IN_242,ImgReg4IN_241,ImgReg4IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState5L (.D ({OutputImg5[271],OutputImg5[270],
                      OutputImg5[269],OutputImg5[268],OutputImg5[267],
                      OutputImg5[266],OutputImg5[265],OutputImg5[264],
                      OutputImg5[263],OutputImg5[262],OutputImg5[261],
                      OutputImg5[260],OutputImg5[259],OutputImg5[258],
                      OutputImg5[257],OutputImg5[256]}), .EN (nx23692), .F ({
                      ImgReg5IN_255,ImgReg5IN_254,ImgReg5IN_253,ImgReg5IN_252,
                      ImgReg5IN_251,ImgReg5IN_250,ImgReg5IN_249,ImgReg5IN_248,
                      ImgReg5IN_247,ImgReg5IN_246,ImgReg5IN_245,ImgReg5IN_244,
                      ImgReg5IN_243,ImgReg5IN_242,ImgReg5IN_241,ImgReg5IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState0N (.D ({DATA[255],DATA[254],DATA[253],
                      DATA[252],DATA[251],DATA[250],DATA[249],DATA[248],
                      DATA[247],DATA[246],DATA[245],DATA[244],DATA[243],
                      DATA[242],DATA[241],DATA[240]}), .EN (nx23658), .F ({
                      ImgReg0IN_255,ImgReg0IN_254,ImgReg0IN_253,ImgReg0IN_252,
                      ImgReg0IN_251,ImgReg0IN_250,ImgReg0IN_249,ImgReg0IN_248,
                      ImgReg0IN_247,ImgReg0IN_246,ImgReg0IN_245,ImgReg0IN_244,
                      ImgReg0IN_243,ImgReg0IN_242,ImgReg0IN_241,ImgReg0IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState1N (.D ({DATA[255],DATA[254],DATA[253],
                      DATA[252],DATA[251],DATA[250],DATA[249],DATA[248],
                      DATA[247],DATA[246],DATA[245],DATA[244],DATA[243],
                      DATA[242],DATA[241],DATA[240]}), .EN (nx23646), .F ({
                      ImgReg1IN_255,ImgReg1IN_254,ImgReg1IN_253,ImgReg1IN_252,
                      ImgReg1IN_251,ImgReg1IN_250,ImgReg1IN_249,ImgReg1IN_248,
                      ImgReg1IN_247,ImgReg1IN_246,ImgReg1IN_245,ImgReg1IN_244,
                      ImgReg1IN_243,ImgReg1IN_242,ImgReg1IN_241,ImgReg1IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState2N (.D ({DATA[255],DATA[254],DATA[253],
                      DATA[252],DATA[251],DATA[250],DATA[249],DATA[248],
                      DATA[247],DATA[246],DATA[245],DATA[244],DATA[243],
                      DATA[242],DATA[241],DATA[240]}), .EN (nx23634), .F ({
                      ImgReg2IN_255,ImgReg2IN_254,ImgReg2IN_253,ImgReg2IN_252,
                      ImgReg2IN_251,ImgReg2IN_250,ImgReg2IN_249,ImgReg2IN_248,
                      ImgReg2IN_247,ImgReg2IN_246,ImgReg2IN_245,ImgReg2IN_244,
                      ImgReg2IN_243,ImgReg2IN_242,ImgReg2IN_241,ImgReg2IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState3N (.D ({DATA[255],DATA[254],DATA[253],
                      DATA[252],DATA[251],DATA[250],DATA[249],DATA[248],
                      DATA[247],DATA[246],DATA[245],DATA[244],DATA[243],
                      DATA[242],DATA[241],DATA[240]}), .EN (nx23622), .F ({
                      ImgReg3IN_255,ImgReg3IN_254,ImgReg3IN_253,ImgReg3IN_252,
                      ImgReg3IN_251,ImgReg3IN_250,ImgReg3IN_249,ImgReg3IN_248,
                      ImgReg3IN_247,ImgReg3IN_246,ImgReg3IN_245,ImgReg3IN_244,
                      ImgReg3IN_243,ImgReg3IN_242,ImgReg3IN_241,ImgReg3IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState4N (.D ({DATA[255],DATA[254],DATA[253],
                      DATA[252],DATA[251],DATA[250],DATA[249],DATA[248],
                      DATA[247],DATA[246],DATA[245],DATA[244],DATA[243],
                      DATA[242],DATA[241],DATA[240]}), .EN (nx23610), .F ({
                      ImgReg4IN_255,ImgReg4IN_254,ImgReg4IN_253,ImgReg4IN_252,
                      ImgReg4IN_251,ImgReg4IN_250,ImgReg4IN_249,ImgReg4IN_248,
                      ImgReg4IN_247,ImgReg4IN_246,ImgReg4IN_245,ImgReg4IN_244,
                      ImgReg4IN_243,ImgReg4IN_242,ImgReg4IN_241,ImgReg4IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState5N (.D ({DATA[255],DATA[254],DATA[253],
                      DATA[252],DATA[251],DATA[250],DATA[249],DATA[248],
                      DATA[247],DATA[246],DATA[245],DATA[244],DATA[243],
                      DATA[242],DATA[241],DATA[240]}), .EN (nx23598), .F ({
                      ImgReg5IN_255,ImgReg5IN_254,ImgReg5IN_253,ImgReg5IN_252,
                      ImgReg5IN_251,ImgReg5IN_250,ImgReg5IN_249,ImgReg5IN_248,
                      ImgReg5IN_247,ImgReg5IN_246,ImgReg5IN_245,ImgReg5IN_244,
                      ImgReg5IN_243,ImgReg5IN_242,ImgReg5IN_241,ImgReg5IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState0U (.D ({OutputImg1[255],OutputImg1[254],
                      OutputImg1[253],OutputImg1[252],OutputImg1[251],
                      OutputImg1[250],OutputImg1[249],OutputImg1[248],
                      OutputImg1[247],OutputImg1[246],OutputImg1[245],
                      OutputImg1[244],OutputImg1[243],OutputImg1[242],
                      OutputImg1[241],OutputImg1[240]}), .EN (nx23806), .F ({
                      ImgReg0IN_255,ImgReg0IN_254,ImgReg0IN_253,ImgReg0IN_252,
                      ImgReg0IN_251,ImgReg0IN_250,ImgReg0IN_249,ImgReg0IN_248,
                      ImgReg0IN_247,ImgReg0IN_246,ImgReg0IN_245,ImgReg0IN_244,
                      ImgReg0IN_243,ImgReg0IN_242,ImgReg0IN_241,ImgReg0IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState1U (.D ({OutputImg2[255],OutputImg2[254],
                      OutputImg2[253],OutputImg2[252],OutputImg2[251],
                      OutputImg2[250],OutputImg2[249],OutputImg2[248],
                      OutputImg2[247],OutputImg2[246],OutputImg2[245],
                      OutputImg2[244],OutputImg2[243],OutputImg2[242],
                      OutputImg2[241],OutputImg2[240]}), .EN (nx23806), .F ({
                      ImgReg1IN_255,ImgReg1IN_254,ImgReg1IN_253,ImgReg1IN_252,
                      ImgReg1IN_251,ImgReg1IN_250,ImgReg1IN_249,ImgReg1IN_248,
                      ImgReg1IN_247,ImgReg1IN_246,ImgReg1IN_245,ImgReg1IN_244,
                      ImgReg1IN_243,ImgReg1IN_242,ImgReg1IN_241,ImgReg1IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState2U (.D ({OutputImg3[255],OutputImg3[254],
                      OutputImg3[253],OutputImg3[252],OutputImg3[251],
                      OutputImg3[250],OutputImg3[249],OutputImg3[248],
                      OutputImg3[247],OutputImg3[246],OutputImg3[245],
                      OutputImg3[244],OutputImg3[243],OutputImg3[242],
                      OutputImg3[241],OutputImg3[240]}), .EN (nx23808), .F ({
                      ImgReg2IN_255,ImgReg2IN_254,ImgReg2IN_253,ImgReg2IN_252,
                      ImgReg2IN_251,ImgReg2IN_250,ImgReg2IN_249,ImgReg2IN_248,
                      ImgReg2IN_247,ImgReg2IN_246,ImgReg2IN_245,ImgReg2IN_244,
                      ImgReg2IN_243,ImgReg2IN_242,ImgReg2IN_241,ImgReg2IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState3U (.D ({OutputImg4[255],OutputImg4[254],
                      OutputImg4[253],OutputImg4[252],OutputImg4[251],
                      OutputImg4[250],OutputImg4[249],OutputImg4[248],
                      OutputImg4[247],OutputImg4[246],OutputImg4[245],
                      OutputImg4[244],OutputImg4[243],OutputImg4[242],
                      OutputImg4[241],OutputImg4[240]}), .EN (nx23808), .F ({
                      ImgReg3IN_255,ImgReg3IN_254,ImgReg3IN_253,ImgReg3IN_252,
                      ImgReg3IN_251,ImgReg3IN_250,ImgReg3IN_249,ImgReg3IN_248,
                      ImgReg3IN_247,ImgReg3IN_246,ImgReg3IN_245,ImgReg3IN_244,
                      ImgReg3IN_243,ImgReg3IN_242,ImgReg3IN_241,ImgReg3IN_240})
                      ) ;
    triStateBuffer_16 loop3_15_TriState4U (.D ({OutputImg5[255],OutputImg5[254],
                      OutputImg5[253],OutputImg5[252],OutputImg5[251],
                      OutputImg5[250],OutputImg5[249],OutputImg5[248],
                      OutputImg5[247],OutputImg5[246],OutputImg5[245],
                      OutputImg5[244],OutputImg5[243],OutputImg5[242],
                      OutputImg5[241],OutputImg5[240]}), .EN (nx23808), .F ({
                      ImgReg4IN_255,ImgReg4IN_254,ImgReg4IN_253,ImgReg4IN_252,
                      ImgReg4IN_251,ImgReg4IN_250,ImgReg4IN_249,ImgReg4IN_248,
                      ImgReg4IN_247,ImgReg4IN_246,ImgReg4IN_245,ImgReg4IN_244,
                      ImgReg4IN_243,ImgReg4IN_242,ImgReg4IN_241,ImgReg4IN_240})
                      ) ;
    nBitRegister_16 loop3_15_reg1 (.D ({ImgReg0IN_255,ImgReg0IN_254,
                    ImgReg0IN_253,ImgReg0IN_252,ImgReg0IN_251,ImgReg0IN_250,
                    ImgReg0IN_249,ImgReg0IN_248,ImgReg0IN_247,ImgReg0IN_246,
                    ImgReg0IN_245,ImgReg0IN_244,ImgReg0IN_243,ImgReg0IN_242,
                    ImgReg0IN_241,ImgReg0IN_240}), .CLK (nx23918), .RST (RST), .EN (
                    nx23722), .Q ({OutputImg0[255],OutputImg0[254],
                    OutputImg0[253],OutputImg0[252],OutputImg0[251],
                    OutputImg0[250],OutputImg0[249],OutputImg0[248],
                    OutputImg0[247],OutputImg0[246],OutputImg0[245],
                    OutputImg0[244],OutputImg0[243],OutputImg0[242],
                    OutputImg0[241],OutputImg0[240]})) ;
    nBitRegister_16 loop3_15_reg2 (.D ({ImgReg1IN_255,ImgReg1IN_254,
                    ImgReg1IN_253,ImgReg1IN_252,ImgReg1IN_251,ImgReg1IN_250,
                    ImgReg1IN_249,ImgReg1IN_248,ImgReg1IN_247,ImgReg1IN_246,
                    ImgReg1IN_245,ImgReg1IN_244,ImgReg1IN_243,ImgReg1IN_242,
                    ImgReg1IN_241,ImgReg1IN_240}), .CLK (nx23920), .RST (RST), .EN (
                    nx23732), .Q ({OutputImg1[255],OutputImg1[254],
                    OutputImg1[253],OutputImg1[252],OutputImg1[251],
                    OutputImg1[250],OutputImg1[249],OutputImg1[248],
                    OutputImg1[247],OutputImg1[246],OutputImg1[245],
                    OutputImg1[244],OutputImg1[243],OutputImg1[242],
                    OutputImg1[241],OutputImg1[240]})) ;
    nBitRegister_16 loop3_15_reg3 (.D ({ImgReg2IN_255,ImgReg2IN_254,
                    ImgReg2IN_253,ImgReg2IN_252,ImgReg2IN_251,ImgReg2IN_250,
                    ImgReg2IN_249,ImgReg2IN_248,ImgReg2IN_247,ImgReg2IN_246,
                    ImgReg2IN_245,ImgReg2IN_244,ImgReg2IN_243,ImgReg2IN_242,
                    ImgReg2IN_241,ImgReg2IN_240}), .CLK (nx23920), .RST (RST), .EN (
                    nx23742), .Q ({OutputImg2[255],OutputImg2[254],
                    OutputImg2[253],OutputImg2[252],OutputImg2[251],
                    OutputImg2[250],OutputImg2[249],OutputImg2[248],
                    OutputImg2[247],OutputImg2[246],OutputImg2[245],
                    OutputImg2[244],OutputImg2[243],OutputImg2[242],
                    OutputImg2[241],OutputImg2[240]})) ;
    nBitRegister_16 loop3_15_reg4 (.D ({ImgReg3IN_255,ImgReg3IN_254,
                    ImgReg3IN_253,ImgReg3IN_252,ImgReg3IN_251,ImgReg3IN_250,
                    ImgReg3IN_249,ImgReg3IN_248,ImgReg3IN_247,ImgReg3IN_246,
                    ImgReg3IN_245,ImgReg3IN_244,ImgReg3IN_243,ImgReg3IN_242,
                    ImgReg3IN_241,ImgReg3IN_240}), .CLK (nx23922), .RST (RST), .EN (
                    nx23752), .Q ({OutputImg3[255],OutputImg3[254],
                    OutputImg3[253],OutputImg3[252],OutputImg3[251],
                    OutputImg3[250],OutputImg3[249],OutputImg3[248],
                    OutputImg3[247],OutputImg3[246],OutputImg3[245],
                    OutputImg3[244],OutputImg3[243],OutputImg3[242],
                    OutputImg3[241],OutputImg3[240]})) ;
    nBitRegister_16 loop3_15_reg5 (.D ({ImgReg4IN_255,ImgReg4IN_254,
                    ImgReg4IN_253,ImgReg4IN_252,ImgReg4IN_251,ImgReg4IN_250,
                    ImgReg4IN_249,ImgReg4IN_248,ImgReg4IN_247,ImgReg4IN_246,
                    ImgReg4IN_245,ImgReg4IN_244,ImgReg4IN_243,ImgReg4IN_242,
                    ImgReg4IN_241,ImgReg4IN_240}), .CLK (nx23922), .RST (RST), .EN (
                    nx23762), .Q ({OutputImg4[255],OutputImg4[254],
                    OutputImg4[253],OutputImg4[252],OutputImg4[251],
                    OutputImg4[250],OutputImg4[249],OutputImg4[248],
                    OutputImg4[247],OutputImg4[246],OutputImg4[245],
                    OutputImg4[244],OutputImg4[243],OutputImg4[242],
                    OutputImg4[241],OutputImg4[240]})) ;
    nBitRegister_16 loop3_15_reg6 (.D ({ImgReg5IN_255,ImgReg5IN_254,
                    ImgReg5IN_253,ImgReg5IN_252,ImgReg5IN_251,ImgReg5IN_250,
                    ImgReg5IN_249,ImgReg5IN_248,ImgReg5IN_247,ImgReg5IN_246,
                    ImgReg5IN_245,ImgReg5IN_244,ImgReg5IN_243,ImgReg5IN_242,
                    ImgReg5IN_241,ImgReg5IN_240}), .CLK (nx23924), .RST (RST), .EN (
                    nx23772), .Q ({OutputImg5[255],OutputImg5[254],
                    OutputImg5[253],OutputImg5[252],OutputImg5[251],
                    OutputImg5[250],OutputImg5[249],OutputImg5[248],
                    OutputImg5[247],OutputImg5[246],OutputImg5[245],
                    OutputImg5[244],OutputImg5[243],OutputImg5[242],
                    OutputImg5[241],OutputImg5[240]})) ;
    triStateBuffer_16 loop3_16_TriState0L (.D ({OutputImg0[287],OutputImg0[286],
                      OutputImg0[285],OutputImg0[284],OutputImg0[283],
                      OutputImg0[282],OutputImg0[281],OutputImg0[280],
                      OutputImg0[279],OutputImg0[278],OutputImg0[277],
                      OutputImg0[276],OutputImg0[275],OutputImg0[274],
                      OutputImg0[273],OutputImg0[272]}), .EN (nx23692), .F ({
                      ImgReg0IN_271,ImgReg0IN_270,ImgReg0IN_269,ImgReg0IN_268,
                      ImgReg0IN_267,ImgReg0IN_266,ImgReg0IN_265,ImgReg0IN_264,
                      ImgReg0IN_263,ImgReg0IN_262,ImgReg0IN_261,ImgReg0IN_260,
                      ImgReg0IN_259,ImgReg0IN_258,ImgReg0IN_257,ImgReg0IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState1L (.D ({OutputImg1[287],OutputImg1[286],
                      OutputImg1[285],OutputImg1[284],OutputImg1[283],
                      OutputImg1[282],OutputImg1[281],OutputImg1[280],
                      OutputImg1[279],OutputImg1[278],OutputImg1[277],
                      OutputImg1[276],OutputImg1[275],OutputImg1[274],
                      OutputImg1[273],OutputImg1[272]}), .EN (nx23692), .F ({
                      ImgReg1IN_271,ImgReg1IN_270,ImgReg1IN_269,ImgReg1IN_268,
                      ImgReg1IN_267,ImgReg1IN_266,ImgReg1IN_265,ImgReg1IN_264,
                      ImgReg1IN_263,ImgReg1IN_262,ImgReg1IN_261,ImgReg1IN_260,
                      ImgReg1IN_259,ImgReg1IN_258,ImgReg1IN_257,ImgReg1IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState2L (.D ({OutputImg2[287],OutputImg2[286],
                      OutputImg2[285],OutputImg2[284],OutputImg2[283],
                      OutputImg2[282],OutputImg2[281],OutputImg2[280],
                      OutputImg2[279],OutputImg2[278],OutputImg2[277],
                      OutputImg2[276],OutputImg2[275],OutputImg2[274],
                      OutputImg2[273],OutputImg2[272]}), .EN (nx23694), .F ({
                      ImgReg2IN_271,ImgReg2IN_270,ImgReg2IN_269,ImgReg2IN_268,
                      ImgReg2IN_267,ImgReg2IN_266,ImgReg2IN_265,ImgReg2IN_264,
                      ImgReg2IN_263,ImgReg2IN_262,ImgReg2IN_261,ImgReg2IN_260,
                      ImgReg2IN_259,ImgReg2IN_258,ImgReg2IN_257,ImgReg2IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState3L (.D ({OutputImg3[287],OutputImg3[286],
                      OutputImg3[285],OutputImg3[284],OutputImg3[283],
                      OutputImg3[282],OutputImg3[281],OutputImg3[280],
                      OutputImg3[279],OutputImg3[278],OutputImg3[277],
                      OutputImg3[276],OutputImg3[275],OutputImg3[274],
                      OutputImg3[273],OutputImg3[272]}), .EN (nx23694), .F ({
                      ImgReg3IN_271,ImgReg3IN_270,ImgReg3IN_269,ImgReg3IN_268,
                      ImgReg3IN_267,ImgReg3IN_266,ImgReg3IN_265,ImgReg3IN_264,
                      ImgReg3IN_263,ImgReg3IN_262,ImgReg3IN_261,ImgReg3IN_260,
                      ImgReg3IN_259,ImgReg3IN_258,ImgReg3IN_257,ImgReg3IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState4L (.D ({OutputImg4[287],OutputImg4[286],
                      OutputImg4[285],OutputImg4[284],OutputImg4[283],
                      OutputImg4[282],OutputImg4[281],OutputImg4[280],
                      OutputImg4[279],OutputImg4[278],OutputImg4[277],
                      OutputImg4[276],OutputImg4[275],OutputImg4[274],
                      OutputImg4[273],OutputImg4[272]}), .EN (nx23694), .F ({
                      ImgReg4IN_271,ImgReg4IN_270,ImgReg4IN_269,ImgReg4IN_268,
                      ImgReg4IN_267,ImgReg4IN_266,ImgReg4IN_265,ImgReg4IN_264,
                      ImgReg4IN_263,ImgReg4IN_262,ImgReg4IN_261,ImgReg4IN_260,
                      ImgReg4IN_259,ImgReg4IN_258,ImgReg4IN_257,ImgReg4IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState5L (.D ({OutputImg5[287],OutputImg5[286],
                      OutputImg5[285],OutputImg5[284],OutputImg5[283],
                      OutputImg5[282],OutputImg5[281],OutputImg5[280],
                      OutputImg5[279],OutputImg5[278],OutputImg5[277],
                      OutputImg5[276],OutputImg5[275],OutputImg5[274],
                      OutputImg5[273],OutputImg5[272]}), .EN (nx23694), .F ({
                      ImgReg5IN_271,ImgReg5IN_270,ImgReg5IN_269,ImgReg5IN_268,
                      ImgReg5IN_267,ImgReg5IN_266,ImgReg5IN_265,ImgReg5IN_264,
                      ImgReg5IN_263,ImgReg5IN_262,ImgReg5IN_261,ImgReg5IN_260,
                      ImgReg5IN_259,ImgReg5IN_258,ImgReg5IN_257,ImgReg5IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState0N (.D ({DATA[271],DATA[270],DATA[269],
                      DATA[268],DATA[267],DATA[266],DATA[265],DATA[264],
                      DATA[263],DATA[262],DATA[261],DATA[260],DATA[259],
                      DATA[258],DATA[257],DATA[256]}), .EN (nx23658), .F ({
                      ImgReg0IN_271,ImgReg0IN_270,ImgReg0IN_269,ImgReg0IN_268,
                      ImgReg0IN_267,ImgReg0IN_266,ImgReg0IN_265,ImgReg0IN_264,
                      ImgReg0IN_263,ImgReg0IN_262,ImgReg0IN_261,ImgReg0IN_260,
                      ImgReg0IN_259,ImgReg0IN_258,ImgReg0IN_257,ImgReg0IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState1N (.D ({DATA[271],DATA[270],DATA[269],
                      DATA[268],DATA[267],DATA[266],DATA[265],DATA[264],
                      DATA[263],DATA[262],DATA[261],DATA[260],DATA[259],
                      DATA[258],DATA[257],DATA[256]}), .EN (nx23646), .F ({
                      ImgReg1IN_271,ImgReg1IN_270,ImgReg1IN_269,ImgReg1IN_268,
                      ImgReg1IN_267,ImgReg1IN_266,ImgReg1IN_265,ImgReg1IN_264,
                      ImgReg1IN_263,ImgReg1IN_262,ImgReg1IN_261,ImgReg1IN_260,
                      ImgReg1IN_259,ImgReg1IN_258,ImgReg1IN_257,ImgReg1IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState2N (.D ({DATA[271],DATA[270],DATA[269],
                      DATA[268],DATA[267],DATA[266],DATA[265],DATA[264],
                      DATA[263],DATA[262],DATA[261],DATA[260],DATA[259],
                      DATA[258],DATA[257],DATA[256]}), .EN (nx23634), .F ({
                      ImgReg2IN_271,ImgReg2IN_270,ImgReg2IN_269,ImgReg2IN_268,
                      ImgReg2IN_267,ImgReg2IN_266,ImgReg2IN_265,ImgReg2IN_264,
                      ImgReg2IN_263,ImgReg2IN_262,ImgReg2IN_261,ImgReg2IN_260,
                      ImgReg2IN_259,ImgReg2IN_258,ImgReg2IN_257,ImgReg2IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState3N (.D ({DATA[271],DATA[270],DATA[269],
                      DATA[268],DATA[267],DATA[266],DATA[265],DATA[264],
                      DATA[263],DATA[262],DATA[261],DATA[260],DATA[259],
                      DATA[258],DATA[257],DATA[256]}), .EN (nx23622), .F ({
                      ImgReg3IN_271,ImgReg3IN_270,ImgReg3IN_269,ImgReg3IN_268,
                      ImgReg3IN_267,ImgReg3IN_266,ImgReg3IN_265,ImgReg3IN_264,
                      ImgReg3IN_263,ImgReg3IN_262,ImgReg3IN_261,ImgReg3IN_260,
                      ImgReg3IN_259,ImgReg3IN_258,ImgReg3IN_257,ImgReg3IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState4N (.D ({DATA[271],DATA[270],DATA[269],
                      DATA[268],DATA[267],DATA[266],DATA[265],DATA[264],
                      DATA[263],DATA[262],DATA[261],DATA[260],DATA[259],
                      DATA[258],DATA[257],DATA[256]}), .EN (nx23610), .F ({
                      ImgReg4IN_271,ImgReg4IN_270,ImgReg4IN_269,ImgReg4IN_268,
                      ImgReg4IN_267,ImgReg4IN_266,ImgReg4IN_265,ImgReg4IN_264,
                      ImgReg4IN_263,ImgReg4IN_262,ImgReg4IN_261,ImgReg4IN_260,
                      ImgReg4IN_259,ImgReg4IN_258,ImgReg4IN_257,ImgReg4IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState5N (.D ({DATA[271],DATA[270],DATA[269],
                      DATA[268],DATA[267],DATA[266],DATA[265],DATA[264],
                      DATA[263],DATA[262],DATA[261],DATA[260],DATA[259],
                      DATA[258],DATA[257],DATA[256]}), .EN (nx23598), .F ({
                      ImgReg5IN_271,ImgReg5IN_270,ImgReg5IN_269,ImgReg5IN_268,
                      ImgReg5IN_267,ImgReg5IN_266,ImgReg5IN_265,ImgReg5IN_264,
                      ImgReg5IN_263,ImgReg5IN_262,ImgReg5IN_261,ImgReg5IN_260,
                      ImgReg5IN_259,ImgReg5IN_258,ImgReg5IN_257,ImgReg5IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState0U (.D ({OutputImg1[271],OutputImg1[270],
                      OutputImg1[269],OutputImg1[268],OutputImg1[267],
                      OutputImg1[266],OutputImg1[265],OutputImg1[264],
                      OutputImg1[263],OutputImg1[262],OutputImg1[261],
                      OutputImg1[260],OutputImg1[259],OutputImg1[258],
                      OutputImg1[257],OutputImg1[256]}), .EN (nx23808), .F ({
                      ImgReg0IN_271,ImgReg0IN_270,ImgReg0IN_269,ImgReg0IN_268,
                      ImgReg0IN_267,ImgReg0IN_266,ImgReg0IN_265,ImgReg0IN_264,
                      ImgReg0IN_263,ImgReg0IN_262,ImgReg0IN_261,ImgReg0IN_260,
                      ImgReg0IN_259,ImgReg0IN_258,ImgReg0IN_257,ImgReg0IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState1U (.D ({OutputImg2[271],OutputImg2[270],
                      OutputImg2[269],OutputImg2[268],OutputImg2[267],
                      OutputImg2[266],OutputImg2[265],OutputImg2[264],
                      OutputImg2[263],OutputImg2[262],OutputImg2[261],
                      OutputImg2[260],OutputImg2[259],OutputImg2[258],
                      OutputImg2[257],OutputImg2[256]}), .EN (nx23808), .F ({
                      ImgReg1IN_271,ImgReg1IN_270,ImgReg1IN_269,ImgReg1IN_268,
                      ImgReg1IN_267,ImgReg1IN_266,ImgReg1IN_265,ImgReg1IN_264,
                      ImgReg1IN_263,ImgReg1IN_262,ImgReg1IN_261,ImgReg1IN_260,
                      ImgReg1IN_259,ImgReg1IN_258,ImgReg1IN_257,ImgReg1IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState2U (.D ({OutputImg3[271],OutputImg3[270],
                      OutputImg3[269],OutputImg3[268],OutputImg3[267],
                      OutputImg3[266],OutputImg3[265],OutputImg3[264],
                      OutputImg3[263],OutputImg3[262],OutputImg3[261],
                      OutputImg3[260],OutputImg3[259],OutputImg3[258],
                      OutputImg3[257],OutputImg3[256]}), .EN (nx23808), .F ({
                      ImgReg2IN_271,ImgReg2IN_270,ImgReg2IN_269,ImgReg2IN_268,
                      ImgReg2IN_267,ImgReg2IN_266,ImgReg2IN_265,ImgReg2IN_264,
                      ImgReg2IN_263,ImgReg2IN_262,ImgReg2IN_261,ImgReg2IN_260,
                      ImgReg2IN_259,ImgReg2IN_258,ImgReg2IN_257,ImgReg2IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState3U (.D ({OutputImg4[271],OutputImg4[270],
                      OutputImg4[269],OutputImg4[268],OutputImg4[267],
                      OutputImg4[266],OutputImg4[265],OutputImg4[264],
                      OutputImg4[263],OutputImg4[262],OutputImg4[261],
                      OutputImg4[260],OutputImg4[259],OutputImg4[258],
                      OutputImg4[257],OutputImg4[256]}), .EN (nx23808), .F ({
                      ImgReg3IN_271,ImgReg3IN_270,ImgReg3IN_269,ImgReg3IN_268,
                      ImgReg3IN_267,ImgReg3IN_266,ImgReg3IN_265,ImgReg3IN_264,
                      ImgReg3IN_263,ImgReg3IN_262,ImgReg3IN_261,ImgReg3IN_260,
                      ImgReg3IN_259,ImgReg3IN_258,ImgReg3IN_257,ImgReg3IN_256})
                      ) ;
    triStateBuffer_16 loop3_16_TriState4U (.D ({OutputImg5[271],OutputImg5[270],
                      OutputImg5[269],OutputImg5[268],OutputImg5[267],
                      OutputImg5[266],OutputImg5[265],OutputImg5[264],
                      OutputImg5[263],OutputImg5[262],OutputImg5[261],
                      OutputImg5[260],OutputImg5[259],OutputImg5[258],
                      OutputImg5[257],OutputImg5[256]}), .EN (nx23810), .F ({
                      ImgReg4IN_271,ImgReg4IN_270,ImgReg4IN_269,ImgReg4IN_268,
                      ImgReg4IN_267,ImgReg4IN_266,ImgReg4IN_265,ImgReg4IN_264,
                      ImgReg4IN_263,ImgReg4IN_262,ImgReg4IN_261,ImgReg4IN_260,
                      ImgReg4IN_259,ImgReg4IN_258,ImgReg4IN_257,ImgReg4IN_256})
                      ) ;
    nBitRegister_16 loop3_16_reg1 (.D ({ImgReg0IN_271,ImgReg0IN_270,
                    ImgReg0IN_269,ImgReg0IN_268,ImgReg0IN_267,ImgReg0IN_266,
                    ImgReg0IN_265,ImgReg0IN_264,ImgReg0IN_263,ImgReg0IN_262,
                    ImgReg0IN_261,ImgReg0IN_260,ImgReg0IN_259,ImgReg0IN_258,
                    ImgReg0IN_257,ImgReg0IN_256}), .CLK (nx23924), .RST (RST), .EN (
                    nx23722), .Q ({OutputImg0[271],OutputImg0[270],
                    OutputImg0[269],OutputImg0[268],OutputImg0[267],
                    OutputImg0[266],OutputImg0[265],OutputImg0[264],
                    OutputImg0[263],OutputImg0[262],OutputImg0[261],
                    OutputImg0[260],OutputImg0[259],OutputImg0[258],
                    OutputImg0[257],OutputImg0[256]})) ;
    nBitRegister_16 loop3_16_reg2 (.D ({ImgReg1IN_271,ImgReg1IN_270,
                    ImgReg1IN_269,ImgReg1IN_268,ImgReg1IN_267,ImgReg1IN_266,
                    ImgReg1IN_265,ImgReg1IN_264,ImgReg1IN_263,ImgReg1IN_262,
                    ImgReg1IN_261,ImgReg1IN_260,ImgReg1IN_259,ImgReg1IN_258,
                    ImgReg1IN_257,ImgReg1IN_256}), .CLK (nx23926), .RST (RST), .EN (
                    nx23732), .Q ({OutputImg1[271],OutputImg1[270],
                    OutputImg1[269],OutputImg1[268],OutputImg1[267],
                    OutputImg1[266],OutputImg1[265],OutputImg1[264],
                    OutputImg1[263],OutputImg1[262],OutputImg1[261],
                    OutputImg1[260],OutputImg1[259],OutputImg1[258],
                    OutputImg1[257],OutputImg1[256]})) ;
    nBitRegister_16 loop3_16_reg3 (.D ({ImgReg2IN_271,ImgReg2IN_270,
                    ImgReg2IN_269,ImgReg2IN_268,ImgReg2IN_267,ImgReg2IN_266,
                    ImgReg2IN_265,ImgReg2IN_264,ImgReg2IN_263,ImgReg2IN_262,
                    ImgReg2IN_261,ImgReg2IN_260,ImgReg2IN_259,ImgReg2IN_258,
                    ImgReg2IN_257,ImgReg2IN_256}), .CLK (nx23926), .RST (RST), .EN (
                    nx23742), .Q ({OutputImg2[271],OutputImg2[270],
                    OutputImg2[269],OutputImg2[268],OutputImg2[267],
                    OutputImg2[266],OutputImg2[265],OutputImg2[264],
                    OutputImg2[263],OutputImg2[262],OutputImg2[261],
                    OutputImg2[260],OutputImg2[259],OutputImg2[258],
                    OutputImg2[257],OutputImg2[256]})) ;
    nBitRegister_16 loop3_16_reg4 (.D ({ImgReg3IN_271,ImgReg3IN_270,
                    ImgReg3IN_269,ImgReg3IN_268,ImgReg3IN_267,ImgReg3IN_266,
                    ImgReg3IN_265,ImgReg3IN_264,ImgReg3IN_263,ImgReg3IN_262,
                    ImgReg3IN_261,ImgReg3IN_260,ImgReg3IN_259,ImgReg3IN_258,
                    ImgReg3IN_257,ImgReg3IN_256}), .CLK (nx23928), .RST (RST), .EN (
                    nx23752), .Q ({OutputImg3[271],OutputImg3[270],
                    OutputImg3[269],OutputImg3[268],OutputImg3[267],
                    OutputImg3[266],OutputImg3[265],OutputImg3[264],
                    OutputImg3[263],OutputImg3[262],OutputImg3[261],
                    OutputImg3[260],OutputImg3[259],OutputImg3[258],
                    OutputImg3[257],OutputImg3[256]})) ;
    nBitRegister_16 loop3_16_reg5 (.D ({ImgReg4IN_271,ImgReg4IN_270,
                    ImgReg4IN_269,ImgReg4IN_268,ImgReg4IN_267,ImgReg4IN_266,
                    ImgReg4IN_265,ImgReg4IN_264,ImgReg4IN_263,ImgReg4IN_262,
                    ImgReg4IN_261,ImgReg4IN_260,ImgReg4IN_259,ImgReg4IN_258,
                    ImgReg4IN_257,ImgReg4IN_256}), .CLK (nx23928), .RST (RST), .EN (
                    nx23762), .Q ({OutputImg4[271],OutputImg4[270],
                    OutputImg4[269],OutputImg4[268],OutputImg4[267],
                    OutputImg4[266],OutputImg4[265],OutputImg4[264],
                    OutputImg4[263],OutputImg4[262],OutputImg4[261],
                    OutputImg4[260],OutputImg4[259],OutputImg4[258],
                    OutputImg4[257],OutputImg4[256]})) ;
    nBitRegister_16 loop3_16_reg6 (.D ({ImgReg5IN_271,ImgReg5IN_270,
                    ImgReg5IN_269,ImgReg5IN_268,ImgReg5IN_267,ImgReg5IN_266,
                    ImgReg5IN_265,ImgReg5IN_264,ImgReg5IN_263,ImgReg5IN_262,
                    ImgReg5IN_261,ImgReg5IN_260,ImgReg5IN_259,ImgReg5IN_258,
                    ImgReg5IN_257,ImgReg5IN_256}), .CLK (nx23930), .RST (RST), .EN (
                    nx23772), .Q ({OutputImg5[271],OutputImg5[270],
                    OutputImg5[269],OutputImg5[268],OutputImg5[267],
                    OutputImg5[266],OutputImg5[265],OutputImg5[264],
                    OutputImg5[263],OutputImg5[262],OutputImg5[261],
                    OutputImg5[260],OutputImg5[259],OutputImg5[258],
                    OutputImg5[257],OutputImg5[256]})) ;
    triStateBuffer_16 loop3_17_TriState0L (.D ({OutputImg0[303],OutputImg0[302],
                      OutputImg0[301],OutputImg0[300],OutputImg0[299],
                      OutputImg0[298],OutputImg0[297],OutputImg0[296],
                      OutputImg0[295],OutputImg0[294],OutputImg0[293],
                      OutputImg0[292],OutputImg0[291],OutputImg0[290],
                      OutputImg0[289],OutputImg0[288]}), .EN (nx23694), .F ({
                      ImgReg0IN_287,ImgReg0IN_286,ImgReg0IN_285,ImgReg0IN_284,
                      ImgReg0IN_283,ImgReg0IN_282,ImgReg0IN_281,ImgReg0IN_280,
                      ImgReg0IN_279,ImgReg0IN_278,ImgReg0IN_277,ImgReg0IN_276,
                      ImgReg0IN_275,ImgReg0IN_274,ImgReg0IN_273,ImgReg0IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState1L (.D ({OutputImg1[303],OutputImg1[302],
                      OutputImg1[301],OutputImg1[300],OutputImg1[299],
                      OutputImg1[298],OutputImg1[297],OutputImg1[296],
                      OutputImg1[295],OutputImg1[294],OutputImg1[293],
                      OutputImg1[292],OutputImg1[291],OutputImg1[290],
                      OutputImg1[289],OutputImg1[288]}), .EN (nx23694), .F ({
                      ImgReg1IN_287,ImgReg1IN_286,ImgReg1IN_285,ImgReg1IN_284,
                      ImgReg1IN_283,ImgReg1IN_282,ImgReg1IN_281,ImgReg1IN_280,
                      ImgReg1IN_279,ImgReg1IN_278,ImgReg1IN_277,ImgReg1IN_276,
                      ImgReg1IN_275,ImgReg1IN_274,ImgReg1IN_273,ImgReg1IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState2L (.D ({OutputImg2[303],OutputImg2[302],
                      OutputImg2[301],OutputImg2[300],OutputImg2[299],
                      OutputImg2[298],OutputImg2[297],OutputImg2[296],
                      OutputImg2[295],OutputImg2[294],OutputImg2[293],
                      OutputImg2[292],OutputImg2[291],OutputImg2[290],
                      OutputImg2[289],OutputImg2[288]}), .EN (nx23694), .F ({
                      ImgReg2IN_287,ImgReg2IN_286,ImgReg2IN_285,ImgReg2IN_284,
                      ImgReg2IN_283,ImgReg2IN_282,ImgReg2IN_281,ImgReg2IN_280,
                      ImgReg2IN_279,ImgReg2IN_278,ImgReg2IN_277,ImgReg2IN_276,
                      ImgReg2IN_275,ImgReg2IN_274,ImgReg2IN_273,ImgReg2IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState3L (.D ({OutputImg3[303],OutputImg3[302],
                      OutputImg3[301],OutputImg3[300],OutputImg3[299],
                      OutputImg3[298],OutputImg3[297],OutputImg3[296],
                      OutputImg3[295],OutputImg3[294],OutputImg3[293],
                      OutputImg3[292],OutputImg3[291],OutputImg3[290],
                      OutputImg3[289],OutputImg3[288]}), .EN (nx23696), .F ({
                      ImgReg3IN_287,ImgReg3IN_286,ImgReg3IN_285,ImgReg3IN_284,
                      ImgReg3IN_283,ImgReg3IN_282,ImgReg3IN_281,ImgReg3IN_280,
                      ImgReg3IN_279,ImgReg3IN_278,ImgReg3IN_277,ImgReg3IN_276,
                      ImgReg3IN_275,ImgReg3IN_274,ImgReg3IN_273,ImgReg3IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState4L (.D ({OutputImg4[303],OutputImg4[302],
                      OutputImg4[301],OutputImg4[300],OutputImg4[299],
                      OutputImg4[298],OutputImg4[297],OutputImg4[296],
                      OutputImg4[295],OutputImg4[294],OutputImg4[293],
                      OutputImg4[292],OutputImg4[291],OutputImg4[290],
                      OutputImg4[289],OutputImg4[288]}), .EN (nx23696), .F ({
                      ImgReg4IN_287,ImgReg4IN_286,ImgReg4IN_285,ImgReg4IN_284,
                      ImgReg4IN_283,ImgReg4IN_282,ImgReg4IN_281,ImgReg4IN_280,
                      ImgReg4IN_279,ImgReg4IN_278,ImgReg4IN_277,ImgReg4IN_276,
                      ImgReg4IN_275,ImgReg4IN_274,ImgReg4IN_273,ImgReg4IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState5L (.D ({OutputImg5[303],OutputImg5[302],
                      OutputImg5[301],OutputImg5[300],OutputImg5[299],
                      OutputImg5[298],OutputImg5[297],OutputImg5[296],
                      OutputImg5[295],OutputImg5[294],OutputImg5[293],
                      OutputImg5[292],OutputImg5[291],OutputImg5[290],
                      OutputImg5[289],OutputImg5[288]}), .EN (nx23696), .F ({
                      ImgReg5IN_287,ImgReg5IN_286,ImgReg5IN_285,ImgReg5IN_284,
                      ImgReg5IN_283,ImgReg5IN_282,ImgReg5IN_281,ImgReg5IN_280,
                      ImgReg5IN_279,ImgReg5IN_278,ImgReg5IN_277,ImgReg5IN_276,
                      ImgReg5IN_275,ImgReg5IN_274,ImgReg5IN_273,ImgReg5IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState0N (.D ({DATA[287],DATA[286],DATA[285],
                      DATA[284],DATA[283],DATA[282],DATA[281],DATA[280],
                      DATA[279],DATA[278],DATA[277],DATA[276],DATA[275],
                      DATA[274],DATA[273],DATA[272]}), .EN (nx23658), .F ({
                      ImgReg0IN_287,ImgReg0IN_286,ImgReg0IN_285,ImgReg0IN_284,
                      ImgReg0IN_283,ImgReg0IN_282,ImgReg0IN_281,ImgReg0IN_280,
                      ImgReg0IN_279,ImgReg0IN_278,ImgReg0IN_277,ImgReg0IN_276,
                      ImgReg0IN_275,ImgReg0IN_274,ImgReg0IN_273,ImgReg0IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState1N (.D ({DATA[287],DATA[286],DATA[285],
                      DATA[284],DATA[283],DATA[282],DATA[281],DATA[280],
                      DATA[279],DATA[278],DATA[277],DATA[276],DATA[275],
                      DATA[274],DATA[273],DATA[272]}), .EN (nx23646), .F ({
                      ImgReg1IN_287,ImgReg1IN_286,ImgReg1IN_285,ImgReg1IN_284,
                      ImgReg1IN_283,ImgReg1IN_282,ImgReg1IN_281,ImgReg1IN_280,
                      ImgReg1IN_279,ImgReg1IN_278,ImgReg1IN_277,ImgReg1IN_276,
                      ImgReg1IN_275,ImgReg1IN_274,ImgReg1IN_273,ImgReg1IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState2N (.D ({DATA[287],DATA[286],DATA[285],
                      DATA[284],DATA[283],DATA[282],DATA[281],DATA[280],
                      DATA[279],DATA[278],DATA[277],DATA[276],DATA[275],
                      DATA[274],DATA[273],DATA[272]}), .EN (nx23634), .F ({
                      ImgReg2IN_287,ImgReg2IN_286,ImgReg2IN_285,ImgReg2IN_284,
                      ImgReg2IN_283,ImgReg2IN_282,ImgReg2IN_281,ImgReg2IN_280,
                      ImgReg2IN_279,ImgReg2IN_278,ImgReg2IN_277,ImgReg2IN_276,
                      ImgReg2IN_275,ImgReg2IN_274,ImgReg2IN_273,ImgReg2IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState3N (.D ({DATA[287],DATA[286],DATA[285],
                      DATA[284],DATA[283],DATA[282],DATA[281],DATA[280],
                      DATA[279],DATA[278],DATA[277],DATA[276],DATA[275],
                      DATA[274],DATA[273],DATA[272]}), .EN (nx23622), .F ({
                      ImgReg3IN_287,ImgReg3IN_286,ImgReg3IN_285,ImgReg3IN_284,
                      ImgReg3IN_283,ImgReg3IN_282,ImgReg3IN_281,ImgReg3IN_280,
                      ImgReg3IN_279,ImgReg3IN_278,ImgReg3IN_277,ImgReg3IN_276,
                      ImgReg3IN_275,ImgReg3IN_274,ImgReg3IN_273,ImgReg3IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState4N (.D ({DATA[287],DATA[286],DATA[285],
                      DATA[284],DATA[283],DATA[282],DATA[281],DATA[280],
                      DATA[279],DATA[278],DATA[277],DATA[276],DATA[275],
                      DATA[274],DATA[273],DATA[272]}), .EN (nx23610), .F ({
                      ImgReg4IN_287,ImgReg4IN_286,ImgReg4IN_285,ImgReg4IN_284,
                      ImgReg4IN_283,ImgReg4IN_282,ImgReg4IN_281,ImgReg4IN_280,
                      ImgReg4IN_279,ImgReg4IN_278,ImgReg4IN_277,ImgReg4IN_276,
                      ImgReg4IN_275,ImgReg4IN_274,ImgReg4IN_273,ImgReg4IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState5N (.D ({DATA[287],DATA[286],DATA[285],
                      DATA[284],DATA[283],DATA[282],DATA[281],DATA[280],
                      DATA[279],DATA[278],DATA[277],DATA[276],DATA[275],
                      DATA[274],DATA[273],DATA[272]}), .EN (nx23598), .F ({
                      ImgReg5IN_287,ImgReg5IN_286,ImgReg5IN_285,ImgReg5IN_284,
                      ImgReg5IN_283,ImgReg5IN_282,ImgReg5IN_281,ImgReg5IN_280,
                      ImgReg5IN_279,ImgReg5IN_278,ImgReg5IN_277,ImgReg5IN_276,
                      ImgReg5IN_275,ImgReg5IN_274,ImgReg5IN_273,ImgReg5IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState0U (.D ({OutputImg1[287],OutputImg1[286],
                      OutputImg1[285],OutputImg1[284],OutputImg1[283],
                      OutputImg1[282],OutputImg1[281],OutputImg1[280],
                      OutputImg1[279],OutputImg1[278],OutputImg1[277],
                      OutputImg1[276],OutputImg1[275],OutputImg1[274],
                      OutputImg1[273],OutputImg1[272]}), .EN (nx23810), .F ({
                      ImgReg0IN_287,ImgReg0IN_286,ImgReg0IN_285,ImgReg0IN_284,
                      ImgReg0IN_283,ImgReg0IN_282,ImgReg0IN_281,ImgReg0IN_280,
                      ImgReg0IN_279,ImgReg0IN_278,ImgReg0IN_277,ImgReg0IN_276,
                      ImgReg0IN_275,ImgReg0IN_274,ImgReg0IN_273,ImgReg0IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState1U (.D ({OutputImg2[287],OutputImg2[286],
                      OutputImg2[285],OutputImg2[284],OutputImg2[283],
                      OutputImg2[282],OutputImg2[281],OutputImg2[280],
                      OutputImg2[279],OutputImg2[278],OutputImg2[277],
                      OutputImg2[276],OutputImg2[275],OutputImg2[274],
                      OutputImg2[273],OutputImg2[272]}), .EN (nx23810), .F ({
                      ImgReg1IN_287,ImgReg1IN_286,ImgReg1IN_285,ImgReg1IN_284,
                      ImgReg1IN_283,ImgReg1IN_282,ImgReg1IN_281,ImgReg1IN_280,
                      ImgReg1IN_279,ImgReg1IN_278,ImgReg1IN_277,ImgReg1IN_276,
                      ImgReg1IN_275,ImgReg1IN_274,ImgReg1IN_273,ImgReg1IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState2U (.D ({OutputImg3[287],OutputImg3[286],
                      OutputImg3[285],OutputImg3[284],OutputImg3[283],
                      OutputImg3[282],OutputImg3[281],OutputImg3[280],
                      OutputImg3[279],OutputImg3[278],OutputImg3[277],
                      OutputImg3[276],OutputImg3[275],OutputImg3[274],
                      OutputImg3[273],OutputImg3[272]}), .EN (nx23810), .F ({
                      ImgReg2IN_287,ImgReg2IN_286,ImgReg2IN_285,ImgReg2IN_284,
                      ImgReg2IN_283,ImgReg2IN_282,ImgReg2IN_281,ImgReg2IN_280,
                      ImgReg2IN_279,ImgReg2IN_278,ImgReg2IN_277,ImgReg2IN_276,
                      ImgReg2IN_275,ImgReg2IN_274,ImgReg2IN_273,ImgReg2IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState3U (.D ({OutputImg4[287],OutputImg4[286],
                      OutputImg4[285],OutputImg4[284],OutputImg4[283],
                      OutputImg4[282],OutputImg4[281],OutputImg4[280],
                      OutputImg4[279],OutputImg4[278],OutputImg4[277],
                      OutputImg4[276],OutputImg4[275],OutputImg4[274],
                      OutputImg4[273],OutputImg4[272]}), .EN (nx23810), .F ({
                      ImgReg3IN_287,ImgReg3IN_286,ImgReg3IN_285,ImgReg3IN_284,
                      ImgReg3IN_283,ImgReg3IN_282,ImgReg3IN_281,ImgReg3IN_280,
                      ImgReg3IN_279,ImgReg3IN_278,ImgReg3IN_277,ImgReg3IN_276,
                      ImgReg3IN_275,ImgReg3IN_274,ImgReg3IN_273,ImgReg3IN_272})
                      ) ;
    triStateBuffer_16 loop3_17_TriState4U (.D ({OutputImg5[287],OutputImg5[286],
                      OutputImg5[285],OutputImg5[284],OutputImg5[283],
                      OutputImg5[282],OutputImg5[281],OutputImg5[280],
                      OutputImg5[279],OutputImg5[278],OutputImg5[277],
                      OutputImg5[276],OutputImg5[275],OutputImg5[274],
                      OutputImg5[273],OutputImg5[272]}), .EN (nx23810), .F ({
                      ImgReg4IN_287,ImgReg4IN_286,ImgReg4IN_285,ImgReg4IN_284,
                      ImgReg4IN_283,ImgReg4IN_282,ImgReg4IN_281,ImgReg4IN_280,
                      ImgReg4IN_279,ImgReg4IN_278,ImgReg4IN_277,ImgReg4IN_276,
                      ImgReg4IN_275,ImgReg4IN_274,ImgReg4IN_273,ImgReg4IN_272})
                      ) ;
    nBitRegister_16 loop3_17_reg1 (.D ({ImgReg0IN_287,ImgReg0IN_286,
                    ImgReg0IN_285,ImgReg0IN_284,ImgReg0IN_283,ImgReg0IN_282,
                    ImgReg0IN_281,ImgReg0IN_280,ImgReg0IN_279,ImgReg0IN_278,
                    ImgReg0IN_277,ImgReg0IN_276,ImgReg0IN_275,ImgReg0IN_274,
                    ImgReg0IN_273,ImgReg0IN_272}), .CLK (nx23930), .RST (RST), .EN (
                    nx23722), .Q ({OutputImg0[287],OutputImg0[286],
                    OutputImg0[285],OutputImg0[284],OutputImg0[283],
                    OutputImg0[282],OutputImg0[281],OutputImg0[280],
                    OutputImg0[279],OutputImg0[278],OutputImg0[277],
                    OutputImg0[276],OutputImg0[275],OutputImg0[274],
                    OutputImg0[273],OutputImg0[272]})) ;
    nBitRegister_16 loop3_17_reg2 (.D ({ImgReg1IN_287,ImgReg1IN_286,
                    ImgReg1IN_285,ImgReg1IN_284,ImgReg1IN_283,ImgReg1IN_282,
                    ImgReg1IN_281,ImgReg1IN_280,ImgReg1IN_279,ImgReg1IN_278,
                    ImgReg1IN_277,ImgReg1IN_276,ImgReg1IN_275,ImgReg1IN_274,
                    ImgReg1IN_273,ImgReg1IN_272}), .CLK (nx23932), .RST (RST), .EN (
                    nx23732), .Q ({OutputImg1[287],OutputImg1[286],
                    OutputImg1[285],OutputImg1[284],OutputImg1[283],
                    OutputImg1[282],OutputImg1[281],OutputImg1[280],
                    OutputImg1[279],OutputImg1[278],OutputImg1[277],
                    OutputImg1[276],OutputImg1[275],OutputImg1[274],
                    OutputImg1[273],OutputImg1[272]})) ;
    nBitRegister_16 loop3_17_reg3 (.D ({ImgReg2IN_287,ImgReg2IN_286,
                    ImgReg2IN_285,ImgReg2IN_284,ImgReg2IN_283,ImgReg2IN_282,
                    ImgReg2IN_281,ImgReg2IN_280,ImgReg2IN_279,ImgReg2IN_278,
                    ImgReg2IN_277,ImgReg2IN_276,ImgReg2IN_275,ImgReg2IN_274,
                    ImgReg2IN_273,ImgReg2IN_272}), .CLK (nx23932), .RST (RST), .EN (
                    nx23742), .Q ({OutputImg2[287],OutputImg2[286],
                    OutputImg2[285],OutputImg2[284],OutputImg2[283],
                    OutputImg2[282],OutputImg2[281],OutputImg2[280],
                    OutputImg2[279],OutputImg2[278],OutputImg2[277],
                    OutputImg2[276],OutputImg2[275],OutputImg2[274],
                    OutputImg2[273],OutputImg2[272]})) ;
    nBitRegister_16 loop3_17_reg4 (.D ({ImgReg3IN_287,ImgReg3IN_286,
                    ImgReg3IN_285,ImgReg3IN_284,ImgReg3IN_283,ImgReg3IN_282,
                    ImgReg3IN_281,ImgReg3IN_280,ImgReg3IN_279,ImgReg3IN_278,
                    ImgReg3IN_277,ImgReg3IN_276,ImgReg3IN_275,ImgReg3IN_274,
                    ImgReg3IN_273,ImgReg3IN_272}), .CLK (nx23934), .RST (RST), .EN (
                    nx23752), .Q ({OutputImg3[287],OutputImg3[286],
                    OutputImg3[285],OutputImg3[284],OutputImg3[283],
                    OutputImg3[282],OutputImg3[281],OutputImg3[280],
                    OutputImg3[279],OutputImg3[278],OutputImg3[277],
                    OutputImg3[276],OutputImg3[275],OutputImg3[274],
                    OutputImg3[273],OutputImg3[272]})) ;
    nBitRegister_16 loop3_17_reg5 (.D ({ImgReg4IN_287,ImgReg4IN_286,
                    ImgReg4IN_285,ImgReg4IN_284,ImgReg4IN_283,ImgReg4IN_282,
                    ImgReg4IN_281,ImgReg4IN_280,ImgReg4IN_279,ImgReg4IN_278,
                    ImgReg4IN_277,ImgReg4IN_276,ImgReg4IN_275,ImgReg4IN_274,
                    ImgReg4IN_273,ImgReg4IN_272}), .CLK (nx23934), .RST (RST), .EN (
                    nx23762), .Q ({OutputImg4[287],OutputImg4[286],
                    OutputImg4[285],OutputImg4[284],OutputImg4[283],
                    OutputImg4[282],OutputImg4[281],OutputImg4[280],
                    OutputImg4[279],OutputImg4[278],OutputImg4[277],
                    OutputImg4[276],OutputImg4[275],OutputImg4[274],
                    OutputImg4[273],OutputImg4[272]})) ;
    nBitRegister_16 loop3_17_reg6 (.D ({ImgReg5IN_287,ImgReg5IN_286,
                    ImgReg5IN_285,ImgReg5IN_284,ImgReg5IN_283,ImgReg5IN_282,
                    ImgReg5IN_281,ImgReg5IN_280,ImgReg5IN_279,ImgReg5IN_278,
                    ImgReg5IN_277,ImgReg5IN_276,ImgReg5IN_275,ImgReg5IN_274,
                    ImgReg5IN_273,ImgReg5IN_272}), .CLK (nx23936), .RST (RST), .EN (
                    nx23772), .Q ({OutputImg5[287],OutputImg5[286],
                    OutputImg5[285],OutputImg5[284],OutputImg5[283],
                    OutputImg5[282],OutputImg5[281],OutputImg5[280],
                    OutputImg5[279],OutputImg5[278],OutputImg5[277],
                    OutputImg5[276],OutputImg5[275],OutputImg5[274],
                    OutputImg5[273],OutputImg5[272]})) ;
    triStateBuffer_16 loop3_18_TriState0L (.D ({OutputImg0[319],OutputImg0[318],
                      OutputImg0[317],OutputImg0[316],OutputImg0[315],
                      OutputImg0[314],OutputImg0[313],OutputImg0[312],
                      OutputImg0[311],OutputImg0[310],OutputImg0[309],
                      OutputImg0[308],OutputImg0[307],OutputImg0[306],
                      OutputImg0[305],OutputImg0[304]}), .EN (nx23696), .F ({
                      ImgReg0IN_303,ImgReg0IN_302,ImgReg0IN_301,ImgReg0IN_300,
                      ImgReg0IN_299,ImgReg0IN_298,ImgReg0IN_297,ImgReg0IN_296,
                      ImgReg0IN_295,ImgReg0IN_294,ImgReg0IN_293,ImgReg0IN_292,
                      ImgReg0IN_291,ImgReg0IN_290,ImgReg0IN_289,ImgReg0IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState1L (.D ({OutputImg1[319],OutputImg1[318],
                      OutputImg1[317],OutputImg1[316],OutputImg1[315],
                      OutputImg1[314],OutputImg1[313],OutputImg1[312],
                      OutputImg1[311],OutputImg1[310],OutputImg1[309],
                      OutputImg1[308],OutputImg1[307],OutputImg1[306],
                      OutputImg1[305],OutputImg1[304]}), .EN (nx23696), .F ({
                      ImgReg1IN_303,ImgReg1IN_302,ImgReg1IN_301,ImgReg1IN_300,
                      ImgReg1IN_299,ImgReg1IN_298,ImgReg1IN_297,ImgReg1IN_296,
                      ImgReg1IN_295,ImgReg1IN_294,ImgReg1IN_293,ImgReg1IN_292,
                      ImgReg1IN_291,ImgReg1IN_290,ImgReg1IN_289,ImgReg1IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState2L (.D ({OutputImg2[319],OutputImg2[318],
                      OutputImg2[317],OutputImg2[316],OutputImg2[315],
                      OutputImg2[314],OutputImg2[313],OutputImg2[312],
                      OutputImg2[311],OutputImg2[310],OutputImg2[309],
                      OutputImg2[308],OutputImg2[307],OutputImg2[306],
                      OutputImg2[305],OutputImg2[304]}), .EN (nx23696), .F ({
                      ImgReg2IN_303,ImgReg2IN_302,ImgReg2IN_301,ImgReg2IN_300,
                      ImgReg2IN_299,ImgReg2IN_298,ImgReg2IN_297,ImgReg2IN_296,
                      ImgReg2IN_295,ImgReg2IN_294,ImgReg2IN_293,ImgReg2IN_292,
                      ImgReg2IN_291,ImgReg2IN_290,ImgReg2IN_289,ImgReg2IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState3L (.D ({OutputImg3[319],OutputImg3[318],
                      OutputImg3[317],OutputImg3[316],OutputImg3[315],
                      OutputImg3[314],OutputImg3[313],OutputImg3[312],
                      OutputImg3[311],OutputImg3[310],OutputImg3[309],
                      OutputImg3[308],OutputImg3[307],OutputImg3[306],
                      OutputImg3[305],OutputImg3[304]}), .EN (nx23696), .F ({
                      ImgReg3IN_303,ImgReg3IN_302,ImgReg3IN_301,ImgReg3IN_300,
                      ImgReg3IN_299,ImgReg3IN_298,ImgReg3IN_297,ImgReg3IN_296,
                      ImgReg3IN_295,ImgReg3IN_294,ImgReg3IN_293,ImgReg3IN_292,
                      ImgReg3IN_291,ImgReg3IN_290,ImgReg3IN_289,ImgReg3IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState4L (.D ({OutputImg4[319],OutputImg4[318],
                      OutputImg4[317],OutputImg4[316],OutputImg4[315],
                      OutputImg4[314],OutputImg4[313],OutputImg4[312],
                      OutputImg4[311],OutputImg4[310],OutputImg4[309],
                      OutputImg4[308],OutputImg4[307],OutputImg4[306],
                      OutputImg4[305],OutputImg4[304]}), .EN (nx23698), .F ({
                      ImgReg4IN_303,ImgReg4IN_302,ImgReg4IN_301,ImgReg4IN_300,
                      ImgReg4IN_299,ImgReg4IN_298,ImgReg4IN_297,ImgReg4IN_296,
                      ImgReg4IN_295,ImgReg4IN_294,ImgReg4IN_293,ImgReg4IN_292,
                      ImgReg4IN_291,ImgReg4IN_290,ImgReg4IN_289,ImgReg4IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState5L (.D ({OutputImg5[319],OutputImg5[318],
                      OutputImg5[317],OutputImg5[316],OutputImg5[315],
                      OutputImg5[314],OutputImg5[313],OutputImg5[312],
                      OutputImg5[311],OutputImg5[310],OutputImg5[309],
                      OutputImg5[308],OutputImg5[307],OutputImg5[306],
                      OutputImg5[305],OutputImg5[304]}), .EN (nx23698), .F ({
                      ImgReg5IN_303,ImgReg5IN_302,ImgReg5IN_301,ImgReg5IN_300,
                      ImgReg5IN_299,ImgReg5IN_298,ImgReg5IN_297,ImgReg5IN_296,
                      ImgReg5IN_295,ImgReg5IN_294,ImgReg5IN_293,ImgReg5IN_292,
                      ImgReg5IN_291,ImgReg5IN_290,ImgReg5IN_289,ImgReg5IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState0N (.D ({DATA[303],DATA[302],DATA[301],
                      DATA[300],DATA[299],DATA[298],DATA[297],DATA[296],
                      DATA[295],DATA[294],DATA[293],DATA[292],DATA[291],
                      DATA[290],DATA[289],DATA[288]}), .EN (nx23658), .F ({
                      ImgReg0IN_303,ImgReg0IN_302,ImgReg0IN_301,ImgReg0IN_300,
                      ImgReg0IN_299,ImgReg0IN_298,ImgReg0IN_297,ImgReg0IN_296,
                      ImgReg0IN_295,ImgReg0IN_294,ImgReg0IN_293,ImgReg0IN_292,
                      ImgReg0IN_291,ImgReg0IN_290,ImgReg0IN_289,ImgReg0IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState1N (.D ({DATA[303],DATA[302],DATA[301],
                      DATA[300],DATA[299],DATA[298],DATA[297],DATA[296],
                      DATA[295],DATA[294],DATA[293],DATA[292],DATA[291],
                      DATA[290],DATA[289],DATA[288]}), .EN (nx23646), .F ({
                      ImgReg1IN_303,ImgReg1IN_302,ImgReg1IN_301,ImgReg1IN_300,
                      ImgReg1IN_299,ImgReg1IN_298,ImgReg1IN_297,ImgReg1IN_296,
                      ImgReg1IN_295,ImgReg1IN_294,ImgReg1IN_293,ImgReg1IN_292,
                      ImgReg1IN_291,ImgReg1IN_290,ImgReg1IN_289,ImgReg1IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState2N (.D ({DATA[303],DATA[302],DATA[301],
                      DATA[300],DATA[299],DATA[298],DATA[297],DATA[296],
                      DATA[295],DATA[294],DATA[293],DATA[292],DATA[291],
                      DATA[290],DATA[289],DATA[288]}), .EN (nx23634), .F ({
                      ImgReg2IN_303,ImgReg2IN_302,ImgReg2IN_301,ImgReg2IN_300,
                      ImgReg2IN_299,ImgReg2IN_298,ImgReg2IN_297,ImgReg2IN_296,
                      ImgReg2IN_295,ImgReg2IN_294,ImgReg2IN_293,ImgReg2IN_292,
                      ImgReg2IN_291,ImgReg2IN_290,ImgReg2IN_289,ImgReg2IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState3N (.D ({DATA[303],DATA[302],DATA[301],
                      DATA[300],DATA[299],DATA[298],DATA[297],DATA[296],
                      DATA[295],DATA[294],DATA[293],DATA[292],DATA[291],
                      DATA[290],DATA[289],DATA[288]}), .EN (nx23622), .F ({
                      ImgReg3IN_303,ImgReg3IN_302,ImgReg3IN_301,ImgReg3IN_300,
                      ImgReg3IN_299,ImgReg3IN_298,ImgReg3IN_297,ImgReg3IN_296,
                      ImgReg3IN_295,ImgReg3IN_294,ImgReg3IN_293,ImgReg3IN_292,
                      ImgReg3IN_291,ImgReg3IN_290,ImgReg3IN_289,ImgReg3IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState4N (.D ({DATA[303],DATA[302],DATA[301],
                      DATA[300],DATA[299],DATA[298],DATA[297],DATA[296],
                      DATA[295],DATA[294],DATA[293],DATA[292],DATA[291],
                      DATA[290],DATA[289],DATA[288]}), .EN (nx23610), .F ({
                      ImgReg4IN_303,ImgReg4IN_302,ImgReg4IN_301,ImgReg4IN_300,
                      ImgReg4IN_299,ImgReg4IN_298,ImgReg4IN_297,ImgReg4IN_296,
                      ImgReg4IN_295,ImgReg4IN_294,ImgReg4IN_293,ImgReg4IN_292,
                      ImgReg4IN_291,ImgReg4IN_290,ImgReg4IN_289,ImgReg4IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState5N (.D ({DATA[303],DATA[302],DATA[301],
                      DATA[300],DATA[299],DATA[298],DATA[297],DATA[296],
                      DATA[295],DATA[294],DATA[293],DATA[292],DATA[291],
                      DATA[290],DATA[289],DATA[288]}), .EN (nx23598), .F ({
                      ImgReg5IN_303,ImgReg5IN_302,ImgReg5IN_301,ImgReg5IN_300,
                      ImgReg5IN_299,ImgReg5IN_298,ImgReg5IN_297,ImgReg5IN_296,
                      ImgReg5IN_295,ImgReg5IN_294,ImgReg5IN_293,ImgReg5IN_292,
                      ImgReg5IN_291,ImgReg5IN_290,ImgReg5IN_289,ImgReg5IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState0U (.D ({OutputImg1[303],OutputImg1[302],
                      OutputImg1[301],OutputImg1[300],OutputImg1[299],
                      OutputImg1[298],OutputImg1[297],OutputImg1[296],
                      OutputImg1[295],OutputImg1[294],OutputImg1[293],
                      OutputImg1[292],OutputImg1[291],OutputImg1[290],
                      OutputImg1[289],OutputImg1[288]}), .EN (nx23810), .F ({
                      ImgReg0IN_303,ImgReg0IN_302,ImgReg0IN_301,ImgReg0IN_300,
                      ImgReg0IN_299,ImgReg0IN_298,ImgReg0IN_297,ImgReg0IN_296,
                      ImgReg0IN_295,ImgReg0IN_294,ImgReg0IN_293,ImgReg0IN_292,
                      ImgReg0IN_291,ImgReg0IN_290,ImgReg0IN_289,ImgReg0IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState1U (.D ({OutputImg2[303],OutputImg2[302],
                      OutputImg2[301],OutputImg2[300],OutputImg2[299],
                      OutputImg2[298],OutputImg2[297],OutputImg2[296],
                      OutputImg2[295],OutputImg2[294],OutputImg2[293],
                      OutputImg2[292],OutputImg2[291],OutputImg2[290],
                      OutputImg2[289],OutputImg2[288]}), .EN (nx23812), .F ({
                      ImgReg1IN_303,ImgReg1IN_302,ImgReg1IN_301,ImgReg1IN_300,
                      ImgReg1IN_299,ImgReg1IN_298,ImgReg1IN_297,ImgReg1IN_296,
                      ImgReg1IN_295,ImgReg1IN_294,ImgReg1IN_293,ImgReg1IN_292,
                      ImgReg1IN_291,ImgReg1IN_290,ImgReg1IN_289,ImgReg1IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState2U (.D ({OutputImg3[303],OutputImg3[302],
                      OutputImg3[301],OutputImg3[300],OutputImg3[299],
                      OutputImg3[298],OutputImg3[297],OutputImg3[296],
                      OutputImg3[295],OutputImg3[294],OutputImg3[293],
                      OutputImg3[292],OutputImg3[291],OutputImg3[290],
                      OutputImg3[289],OutputImg3[288]}), .EN (nx23812), .F ({
                      ImgReg2IN_303,ImgReg2IN_302,ImgReg2IN_301,ImgReg2IN_300,
                      ImgReg2IN_299,ImgReg2IN_298,ImgReg2IN_297,ImgReg2IN_296,
                      ImgReg2IN_295,ImgReg2IN_294,ImgReg2IN_293,ImgReg2IN_292,
                      ImgReg2IN_291,ImgReg2IN_290,ImgReg2IN_289,ImgReg2IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState3U (.D ({OutputImg4[303],OutputImg4[302],
                      OutputImg4[301],OutputImg4[300],OutputImg4[299],
                      OutputImg4[298],OutputImg4[297],OutputImg4[296],
                      OutputImg4[295],OutputImg4[294],OutputImg4[293],
                      OutputImg4[292],OutputImg4[291],OutputImg4[290],
                      OutputImg4[289],OutputImg4[288]}), .EN (nx23812), .F ({
                      ImgReg3IN_303,ImgReg3IN_302,ImgReg3IN_301,ImgReg3IN_300,
                      ImgReg3IN_299,ImgReg3IN_298,ImgReg3IN_297,ImgReg3IN_296,
                      ImgReg3IN_295,ImgReg3IN_294,ImgReg3IN_293,ImgReg3IN_292,
                      ImgReg3IN_291,ImgReg3IN_290,ImgReg3IN_289,ImgReg3IN_288})
                      ) ;
    triStateBuffer_16 loop3_18_TriState4U (.D ({OutputImg5[303],OutputImg5[302],
                      OutputImg5[301],OutputImg5[300],OutputImg5[299],
                      OutputImg5[298],OutputImg5[297],OutputImg5[296],
                      OutputImg5[295],OutputImg5[294],OutputImg5[293],
                      OutputImg5[292],OutputImg5[291],OutputImg5[290],
                      OutputImg5[289],OutputImg5[288]}), .EN (nx23812), .F ({
                      ImgReg4IN_303,ImgReg4IN_302,ImgReg4IN_301,ImgReg4IN_300,
                      ImgReg4IN_299,ImgReg4IN_298,ImgReg4IN_297,ImgReg4IN_296,
                      ImgReg4IN_295,ImgReg4IN_294,ImgReg4IN_293,ImgReg4IN_292,
                      ImgReg4IN_291,ImgReg4IN_290,ImgReg4IN_289,ImgReg4IN_288})
                      ) ;
    nBitRegister_16 loop3_18_reg1 (.D ({ImgReg0IN_303,ImgReg0IN_302,
                    ImgReg0IN_301,ImgReg0IN_300,ImgReg0IN_299,ImgReg0IN_298,
                    ImgReg0IN_297,ImgReg0IN_296,ImgReg0IN_295,ImgReg0IN_294,
                    ImgReg0IN_293,ImgReg0IN_292,ImgReg0IN_291,ImgReg0IN_290,
                    ImgReg0IN_289,ImgReg0IN_288}), .CLK (nx23936), .RST (RST), .EN (
                    nx23722), .Q ({OutputImg0[303],OutputImg0[302],
                    OutputImg0[301],OutputImg0[300],OutputImg0[299],
                    OutputImg0[298],OutputImg0[297],OutputImg0[296],
                    OutputImg0[295],OutputImg0[294],OutputImg0[293],
                    OutputImg0[292],OutputImg0[291],OutputImg0[290],
                    OutputImg0[289],OutputImg0[288]})) ;
    nBitRegister_16 loop3_18_reg2 (.D ({ImgReg1IN_303,ImgReg1IN_302,
                    ImgReg1IN_301,ImgReg1IN_300,ImgReg1IN_299,ImgReg1IN_298,
                    ImgReg1IN_297,ImgReg1IN_296,ImgReg1IN_295,ImgReg1IN_294,
                    ImgReg1IN_293,ImgReg1IN_292,ImgReg1IN_291,ImgReg1IN_290,
                    ImgReg1IN_289,ImgReg1IN_288}), .CLK (nx23938), .RST (RST), .EN (
                    nx23732), .Q ({OutputImg1[303],OutputImg1[302],
                    OutputImg1[301],OutputImg1[300],OutputImg1[299],
                    OutputImg1[298],OutputImg1[297],OutputImg1[296],
                    OutputImg1[295],OutputImg1[294],OutputImg1[293],
                    OutputImg1[292],OutputImg1[291],OutputImg1[290],
                    OutputImg1[289],OutputImg1[288]})) ;
    nBitRegister_16 loop3_18_reg3 (.D ({ImgReg2IN_303,ImgReg2IN_302,
                    ImgReg2IN_301,ImgReg2IN_300,ImgReg2IN_299,ImgReg2IN_298,
                    ImgReg2IN_297,ImgReg2IN_296,ImgReg2IN_295,ImgReg2IN_294,
                    ImgReg2IN_293,ImgReg2IN_292,ImgReg2IN_291,ImgReg2IN_290,
                    ImgReg2IN_289,ImgReg2IN_288}), .CLK (nx23938), .RST (RST), .EN (
                    nx23742), .Q ({OutputImg2[303],OutputImg2[302],
                    OutputImg2[301],OutputImg2[300],OutputImg2[299],
                    OutputImg2[298],OutputImg2[297],OutputImg2[296],
                    OutputImg2[295],OutputImg2[294],OutputImg2[293],
                    OutputImg2[292],OutputImg2[291],OutputImg2[290],
                    OutputImg2[289],OutputImg2[288]})) ;
    nBitRegister_16 loop3_18_reg4 (.D ({ImgReg3IN_303,ImgReg3IN_302,
                    ImgReg3IN_301,ImgReg3IN_300,ImgReg3IN_299,ImgReg3IN_298,
                    ImgReg3IN_297,ImgReg3IN_296,ImgReg3IN_295,ImgReg3IN_294,
                    ImgReg3IN_293,ImgReg3IN_292,ImgReg3IN_291,ImgReg3IN_290,
                    ImgReg3IN_289,ImgReg3IN_288}), .CLK (nx23940), .RST (RST), .EN (
                    nx23752), .Q ({OutputImg3[303],OutputImg3[302],
                    OutputImg3[301],OutputImg3[300],OutputImg3[299],
                    OutputImg3[298],OutputImg3[297],OutputImg3[296],
                    OutputImg3[295],OutputImg3[294],OutputImg3[293],
                    OutputImg3[292],OutputImg3[291],OutputImg3[290],
                    OutputImg3[289],OutputImg3[288]})) ;
    nBitRegister_16 loop3_18_reg5 (.D ({ImgReg4IN_303,ImgReg4IN_302,
                    ImgReg4IN_301,ImgReg4IN_300,ImgReg4IN_299,ImgReg4IN_298,
                    ImgReg4IN_297,ImgReg4IN_296,ImgReg4IN_295,ImgReg4IN_294,
                    ImgReg4IN_293,ImgReg4IN_292,ImgReg4IN_291,ImgReg4IN_290,
                    ImgReg4IN_289,ImgReg4IN_288}), .CLK (nx23940), .RST (RST), .EN (
                    nx23762), .Q ({OutputImg4[303],OutputImg4[302],
                    OutputImg4[301],OutputImg4[300],OutputImg4[299],
                    OutputImg4[298],OutputImg4[297],OutputImg4[296],
                    OutputImg4[295],OutputImg4[294],OutputImg4[293],
                    OutputImg4[292],OutputImg4[291],OutputImg4[290],
                    OutputImg4[289],OutputImg4[288]})) ;
    nBitRegister_16 loop3_18_reg6 (.D ({ImgReg5IN_303,ImgReg5IN_302,
                    ImgReg5IN_301,ImgReg5IN_300,ImgReg5IN_299,ImgReg5IN_298,
                    ImgReg5IN_297,ImgReg5IN_296,ImgReg5IN_295,ImgReg5IN_294,
                    ImgReg5IN_293,ImgReg5IN_292,ImgReg5IN_291,ImgReg5IN_290,
                    ImgReg5IN_289,ImgReg5IN_288}), .CLK (nx23942), .RST (RST), .EN (
                    nx23772), .Q ({OutputImg5[303],OutputImg5[302],
                    OutputImg5[301],OutputImg5[300],OutputImg5[299],
                    OutputImg5[298],OutputImg5[297],OutputImg5[296],
                    OutputImg5[295],OutputImg5[294],OutputImg5[293],
                    OutputImg5[292],OutputImg5[291],OutputImg5[290],
                    OutputImg5[289],OutputImg5[288]})) ;
    triStateBuffer_16 loop3_19_TriState0L (.D ({OutputImg0[335],OutputImg0[334],
                      OutputImg0[333],OutputImg0[332],OutputImg0[331],
                      OutputImg0[330],OutputImg0[329],OutputImg0[328],
                      OutputImg0[327],OutputImg0[326],OutputImg0[325],
                      OutputImg0[324],OutputImg0[323],OutputImg0[322],
                      OutputImg0[321],OutputImg0[320]}), .EN (nx23698), .F ({
                      ImgReg0IN_319,ImgReg0IN_318,ImgReg0IN_317,ImgReg0IN_316,
                      ImgReg0IN_315,ImgReg0IN_314,ImgReg0IN_313,ImgReg0IN_312,
                      ImgReg0IN_311,ImgReg0IN_310,ImgReg0IN_309,ImgReg0IN_308,
                      ImgReg0IN_307,ImgReg0IN_306,ImgReg0IN_305,ImgReg0IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState1L (.D ({OutputImg1[335],OutputImg1[334],
                      OutputImg1[333],OutputImg1[332],OutputImg1[331],
                      OutputImg1[330],OutputImg1[329],OutputImg1[328],
                      OutputImg1[327],OutputImg1[326],OutputImg1[325],
                      OutputImg1[324],OutputImg1[323],OutputImg1[322],
                      OutputImg1[321],OutputImg1[320]}), .EN (nx23698), .F ({
                      ImgReg1IN_319,ImgReg1IN_318,ImgReg1IN_317,ImgReg1IN_316,
                      ImgReg1IN_315,ImgReg1IN_314,ImgReg1IN_313,ImgReg1IN_312,
                      ImgReg1IN_311,ImgReg1IN_310,ImgReg1IN_309,ImgReg1IN_308,
                      ImgReg1IN_307,ImgReg1IN_306,ImgReg1IN_305,ImgReg1IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState2L (.D ({OutputImg2[335],OutputImg2[334],
                      OutputImg2[333],OutputImg2[332],OutputImg2[331],
                      OutputImg2[330],OutputImg2[329],OutputImg2[328],
                      OutputImg2[327],OutputImg2[326],OutputImg2[325],
                      OutputImg2[324],OutputImg2[323],OutputImg2[322],
                      OutputImg2[321],OutputImg2[320]}), .EN (nx23698), .F ({
                      ImgReg2IN_319,ImgReg2IN_318,ImgReg2IN_317,ImgReg2IN_316,
                      ImgReg2IN_315,ImgReg2IN_314,ImgReg2IN_313,ImgReg2IN_312,
                      ImgReg2IN_311,ImgReg2IN_310,ImgReg2IN_309,ImgReg2IN_308,
                      ImgReg2IN_307,ImgReg2IN_306,ImgReg2IN_305,ImgReg2IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState3L (.D ({OutputImg3[335],OutputImg3[334],
                      OutputImg3[333],OutputImg3[332],OutputImg3[331],
                      OutputImg3[330],OutputImg3[329],OutputImg3[328],
                      OutputImg3[327],OutputImg3[326],OutputImg3[325],
                      OutputImg3[324],OutputImg3[323],OutputImg3[322],
                      OutputImg3[321],OutputImg3[320]}), .EN (nx23698), .F ({
                      ImgReg3IN_319,ImgReg3IN_318,ImgReg3IN_317,ImgReg3IN_316,
                      ImgReg3IN_315,ImgReg3IN_314,ImgReg3IN_313,ImgReg3IN_312,
                      ImgReg3IN_311,ImgReg3IN_310,ImgReg3IN_309,ImgReg3IN_308,
                      ImgReg3IN_307,ImgReg3IN_306,ImgReg3IN_305,ImgReg3IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState4L (.D ({OutputImg4[335],OutputImg4[334],
                      OutputImg4[333],OutputImg4[332],OutputImg4[331],
                      OutputImg4[330],OutputImg4[329],OutputImg4[328],
                      OutputImg4[327],OutputImg4[326],OutputImg4[325],
                      OutputImg4[324],OutputImg4[323],OutputImg4[322],
                      OutputImg4[321],OutputImg4[320]}), .EN (nx23698), .F ({
                      ImgReg4IN_319,ImgReg4IN_318,ImgReg4IN_317,ImgReg4IN_316,
                      ImgReg4IN_315,ImgReg4IN_314,ImgReg4IN_313,ImgReg4IN_312,
                      ImgReg4IN_311,ImgReg4IN_310,ImgReg4IN_309,ImgReg4IN_308,
                      ImgReg4IN_307,ImgReg4IN_306,ImgReg4IN_305,ImgReg4IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState5L (.D ({OutputImg5[335],OutputImg5[334],
                      OutputImg5[333],OutputImg5[332],OutputImg5[331],
                      OutputImg5[330],OutputImg5[329],OutputImg5[328],
                      OutputImg5[327],OutputImg5[326],OutputImg5[325],
                      OutputImg5[324],OutputImg5[323],OutputImg5[322],
                      OutputImg5[321],OutputImg5[320]}), .EN (nx23700), .F ({
                      ImgReg5IN_319,ImgReg5IN_318,ImgReg5IN_317,ImgReg5IN_316,
                      ImgReg5IN_315,ImgReg5IN_314,ImgReg5IN_313,ImgReg5IN_312,
                      ImgReg5IN_311,ImgReg5IN_310,ImgReg5IN_309,ImgReg5IN_308,
                      ImgReg5IN_307,ImgReg5IN_306,ImgReg5IN_305,ImgReg5IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState0N (.D ({DATA[319],DATA[318],DATA[317],
                      DATA[316],DATA[315],DATA[314],DATA[313],DATA[312],
                      DATA[311],DATA[310],DATA[309],DATA[308],DATA[307],
                      DATA[306],DATA[305],DATA[304]}), .EN (nx23658), .F ({
                      ImgReg0IN_319,ImgReg0IN_318,ImgReg0IN_317,ImgReg0IN_316,
                      ImgReg0IN_315,ImgReg0IN_314,ImgReg0IN_313,ImgReg0IN_312,
                      ImgReg0IN_311,ImgReg0IN_310,ImgReg0IN_309,ImgReg0IN_308,
                      ImgReg0IN_307,ImgReg0IN_306,ImgReg0IN_305,ImgReg0IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState1N (.D ({DATA[319],DATA[318],DATA[317],
                      DATA[316],DATA[315],DATA[314],DATA[313],DATA[312],
                      DATA[311],DATA[310],DATA[309],DATA[308],DATA[307],
                      DATA[306],DATA[305],DATA[304]}), .EN (nx23646), .F ({
                      ImgReg1IN_319,ImgReg1IN_318,ImgReg1IN_317,ImgReg1IN_316,
                      ImgReg1IN_315,ImgReg1IN_314,ImgReg1IN_313,ImgReg1IN_312,
                      ImgReg1IN_311,ImgReg1IN_310,ImgReg1IN_309,ImgReg1IN_308,
                      ImgReg1IN_307,ImgReg1IN_306,ImgReg1IN_305,ImgReg1IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState2N (.D ({DATA[319],DATA[318],DATA[317],
                      DATA[316],DATA[315],DATA[314],DATA[313],DATA[312],
                      DATA[311],DATA[310],DATA[309],DATA[308],DATA[307],
                      DATA[306],DATA[305],DATA[304]}), .EN (nx23634), .F ({
                      ImgReg2IN_319,ImgReg2IN_318,ImgReg2IN_317,ImgReg2IN_316,
                      ImgReg2IN_315,ImgReg2IN_314,ImgReg2IN_313,ImgReg2IN_312,
                      ImgReg2IN_311,ImgReg2IN_310,ImgReg2IN_309,ImgReg2IN_308,
                      ImgReg2IN_307,ImgReg2IN_306,ImgReg2IN_305,ImgReg2IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState3N (.D ({DATA[319],DATA[318],DATA[317],
                      DATA[316],DATA[315],DATA[314],DATA[313],DATA[312],
                      DATA[311],DATA[310],DATA[309],DATA[308],DATA[307],
                      DATA[306],DATA[305],DATA[304]}), .EN (nx23622), .F ({
                      ImgReg3IN_319,ImgReg3IN_318,ImgReg3IN_317,ImgReg3IN_316,
                      ImgReg3IN_315,ImgReg3IN_314,ImgReg3IN_313,ImgReg3IN_312,
                      ImgReg3IN_311,ImgReg3IN_310,ImgReg3IN_309,ImgReg3IN_308,
                      ImgReg3IN_307,ImgReg3IN_306,ImgReg3IN_305,ImgReg3IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState4N (.D ({DATA[319],DATA[318],DATA[317],
                      DATA[316],DATA[315],DATA[314],DATA[313],DATA[312],
                      DATA[311],DATA[310],DATA[309],DATA[308],DATA[307],
                      DATA[306],DATA[305],DATA[304]}), .EN (nx23610), .F ({
                      ImgReg4IN_319,ImgReg4IN_318,ImgReg4IN_317,ImgReg4IN_316,
                      ImgReg4IN_315,ImgReg4IN_314,ImgReg4IN_313,ImgReg4IN_312,
                      ImgReg4IN_311,ImgReg4IN_310,ImgReg4IN_309,ImgReg4IN_308,
                      ImgReg4IN_307,ImgReg4IN_306,ImgReg4IN_305,ImgReg4IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState5N (.D ({DATA[319],DATA[318],DATA[317],
                      DATA[316],DATA[315],DATA[314],DATA[313],DATA[312],
                      DATA[311],DATA[310],DATA[309],DATA[308],DATA[307],
                      DATA[306],DATA[305],DATA[304]}), .EN (nx23598), .F ({
                      ImgReg5IN_319,ImgReg5IN_318,ImgReg5IN_317,ImgReg5IN_316,
                      ImgReg5IN_315,ImgReg5IN_314,ImgReg5IN_313,ImgReg5IN_312,
                      ImgReg5IN_311,ImgReg5IN_310,ImgReg5IN_309,ImgReg5IN_308,
                      ImgReg5IN_307,ImgReg5IN_306,ImgReg5IN_305,ImgReg5IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState0U (.D ({OutputImg1[319],OutputImg1[318],
                      OutputImg1[317],OutputImg1[316],OutputImg1[315],
                      OutputImg1[314],OutputImg1[313],OutputImg1[312],
                      OutputImg1[311],OutputImg1[310],OutputImg1[309],
                      OutputImg1[308],OutputImg1[307],OutputImg1[306],
                      OutputImg1[305],OutputImg1[304]}), .EN (nx23812), .F ({
                      ImgReg0IN_319,ImgReg0IN_318,ImgReg0IN_317,ImgReg0IN_316,
                      ImgReg0IN_315,ImgReg0IN_314,ImgReg0IN_313,ImgReg0IN_312,
                      ImgReg0IN_311,ImgReg0IN_310,ImgReg0IN_309,ImgReg0IN_308,
                      ImgReg0IN_307,ImgReg0IN_306,ImgReg0IN_305,ImgReg0IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState1U (.D ({OutputImg2[319],OutputImg2[318],
                      OutputImg2[317],OutputImg2[316],OutputImg2[315],
                      OutputImg2[314],OutputImg2[313],OutputImg2[312],
                      OutputImg2[311],OutputImg2[310],OutputImg2[309],
                      OutputImg2[308],OutputImg2[307],OutputImg2[306],
                      OutputImg2[305],OutputImg2[304]}), .EN (nx23812), .F ({
                      ImgReg1IN_319,ImgReg1IN_318,ImgReg1IN_317,ImgReg1IN_316,
                      ImgReg1IN_315,ImgReg1IN_314,ImgReg1IN_313,ImgReg1IN_312,
                      ImgReg1IN_311,ImgReg1IN_310,ImgReg1IN_309,ImgReg1IN_308,
                      ImgReg1IN_307,ImgReg1IN_306,ImgReg1IN_305,ImgReg1IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState2U (.D ({OutputImg3[319],OutputImg3[318],
                      OutputImg3[317],OutputImg3[316],OutputImg3[315],
                      OutputImg3[314],OutputImg3[313],OutputImg3[312],
                      OutputImg3[311],OutputImg3[310],OutputImg3[309],
                      OutputImg3[308],OutputImg3[307],OutputImg3[306],
                      OutputImg3[305],OutputImg3[304]}), .EN (nx23812), .F ({
                      ImgReg2IN_319,ImgReg2IN_318,ImgReg2IN_317,ImgReg2IN_316,
                      ImgReg2IN_315,ImgReg2IN_314,ImgReg2IN_313,ImgReg2IN_312,
                      ImgReg2IN_311,ImgReg2IN_310,ImgReg2IN_309,ImgReg2IN_308,
                      ImgReg2IN_307,ImgReg2IN_306,ImgReg2IN_305,ImgReg2IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState3U (.D ({OutputImg4[319],OutputImg4[318],
                      OutputImg4[317],OutputImg4[316],OutputImg4[315],
                      OutputImg4[314],OutputImg4[313],OutputImg4[312],
                      OutputImg4[311],OutputImg4[310],OutputImg4[309],
                      OutputImg4[308],OutputImg4[307],OutputImg4[306],
                      OutputImg4[305],OutputImg4[304]}), .EN (nx23814), .F ({
                      ImgReg3IN_319,ImgReg3IN_318,ImgReg3IN_317,ImgReg3IN_316,
                      ImgReg3IN_315,ImgReg3IN_314,ImgReg3IN_313,ImgReg3IN_312,
                      ImgReg3IN_311,ImgReg3IN_310,ImgReg3IN_309,ImgReg3IN_308,
                      ImgReg3IN_307,ImgReg3IN_306,ImgReg3IN_305,ImgReg3IN_304})
                      ) ;
    triStateBuffer_16 loop3_19_TriState4U (.D ({OutputImg5[319],OutputImg5[318],
                      OutputImg5[317],OutputImg5[316],OutputImg5[315],
                      OutputImg5[314],OutputImg5[313],OutputImg5[312],
                      OutputImg5[311],OutputImg5[310],OutputImg5[309],
                      OutputImg5[308],OutputImg5[307],OutputImg5[306],
                      OutputImg5[305],OutputImg5[304]}), .EN (nx23814), .F ({
                      ImgReg4IN_319,ImgReg4IN_318,ImgReg4IN_317,ImgReg4IN_316,
                      ImgReg4IN_315,ImgReg4IN_314,ImgReg4IN_313,ImgReg4IN_312,
                      ImgReg4IN_311,ImgReg4IN_310,ImgReg4IN_309,ImgReg4IN_308,
                      ImgReg4IN_307,ImgReg4IN_306,ImgReg4IN_305,ImgReg4IN_304})
                      ) ;
    nBitRegister_16 loop3_19_reg1 (.D ({ImgReg0IN_319,ImgReg0IN_318,
                    ImgReg0IN_317,ImgReg0IN_316,ImgReg0IN_315,ImgReg0IN_314,
                    ImgReg0IN_313,ImgReg0IN_312,ImgReg0IN_311,ImgReg0IN_310,
                    ImgReg0IN_309,ImgReg0IN_308,ImgReg0IN_307,ImgReg0IN_306,
                    ImgReg0IN_305,ImgReg0IN_304}), .CLK (nx23942), .RST (RST), .EN (
                    nx23722), .Q ({OutputImg0[319],OutputImg0[318],
                    OutputImg0[317],OutputImg0[316],OutputImg0[315],
                    OutputImg0[314],OutputImg0[313],OutputImg0[312],
                    OutputImg0[311],OutputImg0[310],OutputImg0[309],
                    OutputImg0[308],OutputImg0[307],OutputImg0[306],
                    OutputImg0[305],OutputImg0[304]})) ;
    nBitRegister_16 loop3_19_reg2 (.D ({ImgReg1IN_319,ImgReg1IN_318,
                    ImgReg1IN_317,ImgReg1IN_316,ImgReg1IN_315,ImgReg1IN_314,
                    ImgReg1IN_313,ImgReg1IN_312,ImgReg1IN_311,ImgReg1IN_310,
                    ImgReg1IN_309,ImgReg1IN_308,ImgReg1IN_307,ImgReg1IN_306,
                    ImgReg1IN_305,ImgReg1IN_304}), .CLK (nx23944), .RST (RST), .EN (
                    nx23732), .Q ({OutputImg1[319],OutputImg1[318],
                    OutputImg1[317],OutputImg1[316],OutputImg1[315],
                    OutputImg1[314],OutputImg1[313],OutputImg1[312],
                    OutputImg1[311],OutputImg1[310],OutputImg1[309],
                    OutputImg1[308],OutputImg1[307],OutputImg1[306],
                    OutputImg1[305],OutputImg1[304]})) ;
    nBitRegister_16 loop3_19_reg3 (.D ({ImgReg2IN_319,ImgReg2IN_318,
                    ImgReg2IN_317,ImgReg2IN_316,ImgReg2IN_315,ImgReg2IN_314,
                    ImgReg2IN_313,ImgReg2IN_312,ImgReg2IN_311,ImgReg2IN_310,
                    ImgReg2IN_309,ImgReg2IN_308,ImgReg2IN_307,ImgReg2IN_306,
                    ImgReg2IN_305,ImgReg2IN_304}), .CLK (nx23944), .RST (RST), .EN (
                    nx23742), .Q ({OutputImg2[319],OutputImg2[318],
                    OutputImg2[317],OutputImg2[316],OutputImg2[315],
                    OutputImg2[314],OutputImg2[313],OutputImg2[312],
                    OutputImg2[311],OutputImg2[310],OutputImg2[309],
                    OutputImg2[308],OutputImg2[307],OutputImg2[306],
                    OutputImg2[305],OutputImg2[304]})) ;
    nBitRegister_16 loop3_19_reg4 (.D ({ImgReg3IN_319,ImgReg3IN_318,
                    ImgReg3IN_317,ImgReg3IN_316,ImgReg3IN_315,ImgReg3IN_314,
                    ImgReg3IN_313,ImgReg3IN_312,ImgReg3IN_311,ImgReg3IN_310,
                    ImgReg3IN_309,ImgReg3IN_308,ImgReg3IN_307,ImgReg3IN_306,
                    ImgReg3IN_305,ImgReg3IN_304}), .CLK (nx23946), .RST (RST), .EN (
                    nx23752), .Q ({OutputImg3[319],OutputImg3[318],
                    OutputImg3[317],OutputImg3[316],OutputImg3[315],
                    OutputImg3[314],OutputImg3[313],OutputImg3[312],
                    OutputImg3[311],OutputImg3[310],OutputImg3[309],
                    OutputImg3[308],OutputImg3[307],OutputImg3[306],
                    OutputImg3[305],OutputImg3[304]})) ;
    nBitRegister_16 loop3_19_reg5 (.D ({ImgReg4IN_319,ImgReg4IN_318,
                    ImgReg4IN_317,ImgReg4IN_316,ImgReg4IN_315,ImgReg4IN_314,
                    ImgReg4IN_313,ImgReg4IN_312,ImgReg4IN_311,ImgReg4IN_310,
                    ImgReg4IN_309,ImgReg4IN_308,ImgReg4IN_307,ImgReg4IN_306,
                    ImgReg4IN_305,ImgReg4IN_304}), .CLK (nx23946), .RST (RST), .EN (
                    nx23762), .Q ({OutputImg4[319],OutputImg4[318],
                    OutputImg4[317],OutputImg4[316],OutputImg4[315],
                    OutputImg4[314],OutputImg4[313],OutputImg4[312],
                    OutputImg4[311],OutputImg4[310],OutputImg4[309],
                    OutputImg4[308],OutputImg4[307],OutputImg4[306],
                    OutputImg4[305],OutputImg4[304]})) ;
    nBitRegister_16 loop3_19_reg6 (.D ({ImgReg5IN_319,ImgReg5IN_318,
                    ImgReg5IN_317,ImgReg5IN_316,ImgReg5IN_315,ImgReg5IN_314,
                    ImgReg5IN_313,ImgReg5IN_312,ImgReg5IN_311,ImgReg5IN_310,
                    ImgReg5IN_309,ImgReg5IN_308,ImgReg5IN_307,ImgReg5IN_306,
                    ImgReg5IN_305,ImgReg5IN_304}), .CLK (nx23948), .RST (RST), .EN (
                    nx23772), .Q ({OutputImg5[319],OutputImg5[318],
                    OutputImg5[317],OutputImg5[316],OutputImg5[315],
                    OutputImg5[314],OutputImg5[313],OutputImg5[312],
                    OutputImg5[311],OutputImg5[310],OutputImg5[309],
                    OutputImg5[308],OutputImg5[307],OutputImg5[306],
                    OutputImg5[305],OutputImg5[304]})) ;
    triStateBuffer_16 loop3_20_TriState0L (.D ({OutputImg0[351],OutputImg0[350],
                      OutputImg0[349],OutputImg0[348],OutputImg0[347],
                      OutputImg0[346],OutputImg0[345],OutputImg0[344],
                      OutputImg0[343],OutputImg0[342],OutputImg0[341],
                      OutputImg0[340],OutputImg0[339],OutputImg0[338],
                      OutputImg0[337],OutputImg0[336]}), .EN (nx23700), .F ({
                      ImgReg0IN_335,ImgReg0IN_334,ImgReg0IN_333,ImgReg0IN_332,
                      ImgReg0IN_331,ImgReg0IN_330,ImgReg0IN_329,ImgReg0IN_328,
                      ImgReg0IN_327,ImgReg0IN_326,ImgReg0IN_325,ImgReg0IN_324,
                      ImgReg0IN_323,ImgReg0IN_322,ImgReg0IN_321,ImgReg0IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState1L (.D ({OutputImg1[351],OutputImg1[350],
                      OutputImg1[349],OutputImg1[348],OutputImg1[347],
                      OutputImg1[346],OutputImg1[345],OutputImg1[344],
                      OutputImg1[343],OutputImg1[342],OutputImg1[341],
                      OutputImg1[340],OutputImg1[339],OutputImg1[338],
                      OutputImg1[337],OutputImg1[336]}), .EN (nx23700), .F ({
                      ImgReg1IN_335,ImgReg1IN_334,ImgReg1IN_333,ImgReg1IN_332,
                      ImgReg1IN_331,ImgReg1IN_330,ImgReg1IN_329,ImgReg1IN_328,
                      ImgReg1IN_327,ImgReg1IN_326,ImgReg1IN_325,ImgReg1IN_324,
                      ImgReg1IN_323,ImgReg1IN_322,ImgReg1IN_321,ImgReg1IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState2L (.D ({OutputImg2[351],OutputImg2[350],
                      OutputImg2[349],OutputImg2[348],OutputImg2[347],
                      OutputImg2[346],OutputImg2[345],OutputImg2[344],
                      OutputImg2[343],OutputImg2[342],OutputImg2[341],
                      OutputImg2[340],OutputImg2[339],OutputImg2[338],
                      OutputImg2[337],OutputImg2[336]}), .EN (nx23700), .F ({
                      ImgReg2IN_335,ImgReg2IN_334,ImgReg2IN_333,ImgReg2IN_332,
                      ImgReg2IN_331,ImgReg2IN_330,ImgReg2IN_329,ImgReg2IN_328,
                      ImgReg2IN_327,ImgReg2IN_326,ImgReg2IN_325,ImgReg2IN_324,
                      ImgReg2IN_323,ImgReg2IN_322,ImgReg2IN_321,ImgReg2IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState3L (.D ({OutputImg3[351],OutputImg3[350],
                      OutputImg3[349],OutputImg3[348],OutputImg3[347],
                      OutputImg3[346],OutputImg3[345],OutputImg3[344],
                      OutputImg3[343],OutputImg3[342],OutputImg3[341],
                      OutputImg3[340],OutputImg3[339],OutputImg3[338],
                      OutputImg3[337],OutputImg3[336]}), .EN (nx23700), .F ({
                      ImgReg3IN_335,ImgReg3IN_334,ImgReg3IN_333,ImgReg3IN_332,
                      ImgReg3IN_331,ImgReg3IN_330,ImgReg3IN_329,ImgReg3IN_328,
                      ImgReg3IN_327,ImgReg3IN_326,ImgReg3IN_325,ImgReg3IN_324,
                      ImgReg3IN_323,ImgReg3IN_322,ImgReg3IN_321,ImgReg3IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState4L (.D ({OutputImg4[351],OutputImg4[350],
                      OutputImg4[349],OutputImg4[348],OutputImg4[347],
                      OutputImg4[346],OutputImg4[345],OutputImg4[344],
                      OutputImg4[343],OutputImg4[342],OutputImg4[341],
                      OutputImg4[340],OutputImg4[339],OutputImg4[338],
                      OutputImg4[337],OutputImg4[336]}), .EN (nx23700), .F ({
                      ImgReg4IN_335,ImgReg4IN_334,ImgReg4IN_333,ImgReg4IN_332,
                      ImgReg4IN_331,ImgReg4IN_330,ImgReg4IN_329,ImgReg4IN_328,
                      ImgReg4IN_327,ImgReg4IN_326,ImgReg4IN_325,ImgReg4IN_324,
                      ImgReg4IN_323,ImgReg4IN_322,ImgReg4IN_321,ImgReg4IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState5L (.D ({OutputImg5[351],OutputImg5[350],
                      OutputImg5[349],OutputImg5[348],OutputImg5[347],
                      OutputImg5[346],OutputImg5[345],OutputImg5[344],
                      OutputImg5[343],OutputImg5[342],OutputImg5[341],
                      OutputImg5[340],OutputImg5[339],OutputImg5[338],
                      OutputImg5[337],OutputImg5[336]}), .EN (nx23700), .F ({
                      ImgReg5IN_335,ImgReg5IN_334,ImgReg5IN_333,ImgReg5IN_332,
                      ImgReg5IN_331,ImgReg5IN_330,ImgReg5IN_329,ImgReg5IN_328,
                      ImgReg5IN_327,ImgReg5IN_326,ImgReg5IN_325,ImgReg5IN_324,
                      ImgReg5IN_323,ImgReg5IN_322,ImgReg5IN_321,ImgReg5IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState0N (.D ({DATA[335],DATA[334],DATA[333],
                      DATA[332],DATA[331],DATA[330],DATA[329],DATA[328],
                      DATA[327],DATA[326],DATA[325],DATA[324],DATA[323],
                      DATA[322],DATA[321],DATA[320]}), .EN (nx23658), .F ({
                      ImgReg0IN_335,ImgReg0IN_334,ImgReg0IN_333,ImgReg0IN_332,
                      ImgReg0IN_331,ImgReg0IN_330,ImgReg0IN_329,ImgReg0IN_328,
                      ImgReg0IN_327,ImgReg0IN_326,ImgReg0IN_325,ImgReg0IN_324,
                      ImgReg0IN_323,ImgReg0IN_322,ImgReg0IN_321,ImgReg0IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState1N (.D ({DATA[335],DATA[334],DATA[333],
                      DATA[332],DATA[331],DATA[330],DATA[329],DATA[328],
                      DATA[327],DATA[326],DATA[325],DATA[324],DATA[323],
                      DATA[322],DATA[321],DATA[320]}), .EN (nx23646), .F ({
                      ImgReg1IN_335,ImgReg1IN_334,ImgReg1IN_333,ImgReg1IN_332,
                      ImgReg1IN_331,ImgReg1IN_330,ImgReg1IN_329,ImgReg1IN_328,
                      ImgReg1IN_327,ImgReg1IN_326,ImgReg1IN_325,ImgReg1IN_324,
                      ImgReg1IN_323,ImgReg1IN_322,ImgReg1IN_321,ImgReg1IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState2N (.D ({DATA[335],DATA[334],DATA[333],
                      DATA[332],DATA[331],DATA[330],DATA[329],DATA[328],
                      DATA[327],DATA[326],DATA[325],DATA[324],DATA[323],
                      DATA[322],DATA[321],DATA[320]}), .EN (nx23634), .F ({
                      ImgReg2IN_335,ImgReg2IN_334,ImgReg2IN_333,ImgReg2IN_332,
                      ImgReg2IN_331,ImgReg2IN_330,ImgReg2IN_329,ImgReg2IN_328,
                      ImgReg2IN_327,ImgReg2IN_326,ImgReg2IN_325,ImgReg2IN_324,
                      ImgReg2IN_323,ImgReg2IN_322,ImgReg2IN_321,ImgReg2IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState3N (.D ({DATA[335],DATA[334],DATA[333],
                      DATA[332],DATA[331],DATA[330],DATA[329],DATA[328],
                      DATA[327],DATA[326],DATA[325],DATA[324],DATA[323],
                      DATA[322],DATA[321],DATA[320]}), .EN (nx23622), .F ({
                      ImgReg3IN_335,ImgReg3IN_334,ImgReg3IN_333,ImgReg3IN_332,
                      ImgReg3IN_331,ImgReg3IN_330,ImgReg3IN_329,ImgReg3IN_328,
                      ImgReg3IN_327,ImgReg3IN_326,ImgReg3IN_325,ImgReg3IN_324,
                      ImgReg3IN_323,ImgReg3IN_322,ImgReg3IN_321,ImgReg3IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState4N (.D ({DATA[335],DATA[334],DATA[333],
                      DATA[332],DATA[331],DATA[330],DATA[329],DATA[328],
                      DATA[327],DATA[326],DATA[325],DATA[324],DATA[323],
                      DATA[322],DATA[321],DATA[320]}), .EN (nx23610), .F ({
                      ImgReg4IN_335,ImgReg4IN_334,ImgReg4IN_333,ImgReg4IN_332,
                      ImgReg4IN_331,ImgReg4IN_330,ImgReg4IN_329,ImgReg4IN_328,
                      ImgReg4IN_327,ImgReg4IN_326,ImgReg4IN_325,ImgReg4IN_324,
                      ImgReg4IN_323,ImgReg4IN_322,ImgReg4IN_321,ImgReg4IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState5N (.D ({DATA[335],DATA[334],DATA[333],
                      DATA[332],DATA[331],DATA[330],DATA[329],DATA[328],
                      DATA[327],DATA[326],DATA[325],DATA[324],DATA[323],
                      DATA[322],DATA[321],DATA[320]}), .EN (nx23598), .F ({
                      ImgReg5IN_335,ImgReg5IN_334,ImgReg5IN_333,ImgReg5IN_332,
                      ImgReg5IN_331,ImgReg5IN_330,ImgReg5IN_329,ImgReg5IN_328,
                      ImgReg5IN_327,ImgReg5IN_326,ImgReg5IN_325,ImgReg5IN_324,
                      ImgReg5IN_323,ImgReg5IN_322,ImgReg5IN_321,ImgReg5IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState0U (.D ({OutputImg1[335],OutputImg1[334],
                      OutputImg1[333],OutputImg1[332],OutputImg1[331],
                      OutputImg1[330],OutputImg1[329],OutputImg1[328],
                      OutputImg1[327],OutputImg1[326],OutputImg1[325],
                      OutputImg1[324],OutputImg1[323],OutputImg1[322],
                      OutputImg1[321],OutputImg1[320]}), .EN (nx23814), .F ({
                      ImgReg0IN_335,ImgReg0IN_334,ImgReg0IN_333,ImgReg0IN_332,
                      ImgReg0IN_331,ImgReg0IN_330,ImgReg0IN_329,ImgReg0IN_328,
                      ImgReg0IN_327,ImgReg0IN_326,ImgReg0IN_325,ImgReg0IN_324,
                      ImgReg0IN_323,ImgReg0IN_322,ImgReg0IN_321,ImgReg0IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState1U (.D ({OutputImg2[335],OutputImg2[334],
                      OutputImg2[333],OutputImg2[332],OutputImg2[331],
                      OutputImg2[330],OutputImg2[329],OutputImg2[328],
                      OutputImg2[327],OutputImg2[326],OutputImg2[325],
                      OutputImg2[324],OutputImg2[323],OutputImg2[322],
                      OutputImg2[321],OutputImg2[320]}), .EN (nx23814), .F ({
                      ImgReg1IN_335,ImgReg1IN_334,ImgReg1IN_333,ImgReg1IN_332,
                      ImgReg1IN_331,ImgReg1IN_330,ImgReg1IN_329,ImgReg1IN_328,
                      ImgReg1IN_327,ImgReg1IN_326,ImgReg1IN_325,ImgReg1IN_324,
                      ImgReg1IN_323,ImgReg1IN_322,ImgReg1IN_321,ImgReg1IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState2U (.D ({OutputImg3[335],OutputImg3[334],
                      OutputImg3[333],OutputImg3[332],OutputImg3[331],
                      OutputImg3[330],OutputImg3[329],OutputImg3[328],
                      OutputImg3[327],OutputImg3[326],OutputImg3[325],
                      OutputImg3[324],OutputImg3[323],OutputImg3[322],
                      OutputImg3[321],OutputImg3[320]}), .EN (nx23814), .F ({
                      ImgReg2IN_335,ImgReg2IN_334,ImgReg2IN_333,ImgReg2IN_332,
                      ImgReg2IN_331,ImgReg2IN_330,ImgReg2IN_329,ImgReg2IN_328,
                      ImgReg2IN_327,ImgReg2IN_326,ImgReg2IN_325,ImgReg2IN_324,
                      ImgReg2IN_323,ImgReg2IN_322,ImgReg2IN_321,ImgReg2IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState3U (.D ({OutputImg4[335],OutputImg4[334],
                      OutputImg4[333],OutputImg4[332],OutputImg4[331],
                      OutputImg4[330],OutputImg4[329],OutputImg4[328],
                      OutputImg4[327],OutputImg4[326],OutputImg4[325],
                      OutputImg4[324],OutputImg4[323],OutputImg4[322],
                      OutputImg4[321],OutputImg4[320]}), .EN (nx23814), .F ({
                      ImgReg3IN_335,ImgReg3IN_334,ImgReg3IN_333,ImgReg3IN_332,
                      ImgReg3IN_331,ImgReg3IN_330,ImgReg3IN_329,ImgReg3IN_328,
                      ImgReg3IN_327,ImgReg3IN_326,ImgReg3IN_325,ImgReg3IN_324,
                      ImgReg3IN_323,ImgReg3IN_322,ImgReg3IN_321,ImgReg3IN_320})
                      ) ;
    triStateBuffer_16 loop3_20_TriState4U (.D ({OutputImg5[335],OutputImg5[334],
                      OutputImg5[333],OutputImg5[332],OutputImg5[331],
                      OutputImg5[330],OutputImg5[329],OutputImg5[328],
                      OutputImg5[327],OutputImg5[326],OutputImg5[325],
                      OutputImg5[324],OutputImg5[323],OutputImg5[322],
                      OutputImg5[321],OutputImg5[320]}), .EN (nx23814), .F ({
                      ImgReg4IN_335,ImgReg4IN_334,ImgReg4IN_333,ImgReg4IN_332,
                      ImgReg4IN_331,ImgReg4IN_330,ImgReg4IN_329,ImgReg4IN_328,
                      ImgReg4IN_327,ImgReg4IN_326,ImgReg4IN_325,ImgReg4IN_324,
                      ImgReg4IN_323,ImgReg4IN_322,ImgReg4IN_321,ImgReg4IN_320})
                      ) ;
    nBitRegister_16 loop3_20_reg1 (.D ({ImgReg0IN_335,ImgReg0IN_334,
                    ImgReg0IN_333,ImgReg0IN_332,ImgReg0IN_331,ImgReg0IN_330,
                    ImgReg0IN_329,ImgReg0IN_328,ImgReg0IN_327,ImgReg0IN_326,
                    ImgReg0IN_325,ImgReg0IN_324,ImgReg0IN_323,ImgReg0IN_322,
                    ImgReg0IN_321,ImgReg0IN_320}), .CLK (nx23948), .RST (RST), .EN (
                    nx23722), .Q ({OutputImg0[335],OutputImg0[334],
                    OutputImg0[333],OutputImg0[332],OutputImg0[331],
                    OutputImg0[330],OutputImg0[329],OutputImg0[328],
                    OutputImg0[327],OutputImg0[326],OutputImg0[325],
                    OutputImg0[324],OutputImg0[323],OutputImg0[322],
                    OutputImg0[321],OutputImg0[320]})) ;
    nBitRegister_16 loop3_20_reg2 (.D ({ImgReg1IN_335,ImgReg1IN_334,
                    ImgReg1IN_333,ImgReg1IN_332,ImgReg1IN_331,ImgReg1IN_330,
                    ImgReg1IN_329,ImgReg1IN_328,ImgReg1IN_327,ImgReg1IN_326,
                    ImgReg1IN_325,ImgReg1IN_324,ImgReg1IN_323,ImgReg1IN_322,
                    ImgReg1IN_321,ImgReg1IN_320}), .CLK (nx23950), .RST (RST), .EN (
                    nx23732), .Q ({OutputImg1[335],OutputImg1[334],
                    OutputImg1[333],OutputImg1[332],OutputImg1[331],
                    OutputImg1[330],OutputImg1[329],OutputImg1[328],
                    OutputImg1[327],OutputImg1[326],OutputImg1[325],
                    OutputImg1[324],OutputImg1[323],OutputImg1[322],
                    OutputImg1[321],OutputImg1[320]})) ;
    nBitRegister_16 loop3_20_reg3 (.D ({ImgReg2IN_335,ImgReg2IN_334,
                    ImgReg2IN_333,ImgReg2IN_332,ImgReg2IN_331,ImgReg2IN_330,
                    ImgReg2IN_329,ImgReg2IN_328,ImgReg2IN_327,ImgReg2IN_326,
                    ImgReg2IN_325,ImgReg2IN_324,ImgReg2IN_323,ImgReg2IN_322,
                    ImgReg2IN_321,ImgReg2IN_320}), .CLK (nx23950), .RST (RST), .EN (
                    nx23742), .Q ({OutputImg2[335],OutputImg2[334],
                    OutputImg2[333],OutputImg2[332],OutputImg2[331],
                    OutputImg2[330],OutputImg2[329],OutputImg2[328],
                    OutputImg2[327],OutputImg2[326],OutputImg2[325],
                    OutputImg2[324],OutputImg2[323],OutputImg2[322],
                    OutputImg2[321],OutputImg2[320]})) ;
    nBitRegister_16 loop3_20_reg4 (.D ({ImgReg3IN_335,ImgReg3IN_334,
                    ImgReg3IN_333,ImgReg3IN_332,ImgReg3IN_331,ImgReg3IN_330,
                    ImgReg3IN_329,ImgReg3IN_328,ImgReg3IN_327,ImgReg3IN_326,
                    ImgReg3IN_325,ImgReg3IN_324,ImgReg3IN_323,ImgReg3IN_322,
                    ImgReg3IN_321,ImgReg3IN_320}), .CLK (nx23952), .RST (RST), .EN (
                    nx23752), .Q ({OutputImg3[335],OutputImg3[334],
                    OutputImg3[333],OutputImg3[332],OutputImg3[331],
                    OutputImg3[330],OutputImg3[329],OutputImg3[328],
                    OutputImg3[327],OutputImg3[326],OutputImg3[325],
                    OutputImg3[324],OutputImg3[323],OutputImg3[322],
                    OutputImg3[321],OutputImg3[320]})) ;
    nBitRegister_16 loop3_20_reg5 (.D ({ImgReg4IN_335,ImgReg4IN_334,
                    ImgReg4IN_333,ImgReg4IN_332,ImgReg4IN_331,ImgReg4IN_330,
                    ImgReg4IN_329,ImgReg4IN_328,ImgReg4IN_327,ImgReg4IN_326,
                    ImgReg4IN_325,ImgReg4IN_324,ImgReg4IN_323,ImgReg4IN_322,
                    ImgReg4IN_321,ImgReg4IN_320}), .CLK (nx23952), .RST (RST), .EN (
                    nx23762), .Q ({OutputImg4[335],OutputImg4[334],
                    OutputImg4[333],OutputImg4[332],OutputImg4[331],
                    OutputImg4[330],OutputImg4[329],OutputImg4[328],
                    OutputImg4[327],OutputImg4[326],OutputImg4[325],
                    OutputImg4[324],OutputImg4[323],OutputImg4[322],
                    OutputImg4[321],OutputImg4[320]})) ;
    nBitRegister_16 loop3_20_reg6 (.D ({ImgReg5IN_335,ImgReg5IN_334,
                    ImgReg5IN_333,ImgReg5IN_332,ImgReg5IN_331,ImgReg5IN_330,
                    ImgReg5IN_329,ImgReg5IN_328,ImgReg5IN_327,ImgReg5IN_326,
                    ImgReg5IN_325,ImgReg5IN_324,ImgReg5IN_323,ImgReg5IN_322,
                    ImgReg5IN_321,ImgReg5IN_320}), .CLK (nx23954), .RST (RST), .EN (
                    nx23772), .Q ({OutputImg5[335],OutputImg5[334],
                    OutputImg5[333],OutputImg5[332],OutputImg5[331],
                    OutputImg5[330],OutputImg5[329],OutputImg5[328],
                    OutputImg5[327],OutputImg5[326],OutputImg5[325],
                    OutputImg5[324],OutputImg5[323],OutputImg5[322],
                    OutputImg5[321],OutputImg5[320]})) ;
    triStateBuffer_16 loop3_21_TriState0L (.D ({OutputImg0[367],OutputImg0[366],
                      OutputImg0[365],OutputImg0[364],OutputImg0[363],
                      OutputImg0[362],OutputImg0[361],OutputImg0[360],
                      OutputImg0[359],OutputImg0[358],OutputImg0[357],
                      OutputImg0[356],OutputImg0[355],OutputImg0[354],
                      OutputImg0[353],OutputImg0[352]}), .EN (nx23702), .F ({
                      ImgReg0IN_351,ImgReg0IN_350,ImgReg0IN_349,ImgReg0IN_348,
                      ImgReg0IN_347,ImgReg0IN_346,ImgReg0IN_345,ImgReg0IN_344,
                      ImgReg0IN_343,ImgReg0IN_342,ImgReg0IN_341,ImgReg0IN_340,
                      ImgReg0IN_339,ImgReg0IN_338,ImgReg0IN_337,ImgReg0IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState1L (.D ({OutputImg1[367],OutputImg1[366],
                      OutputImg1[365],OutputImg1[364],OutputImg1[363],
                      OutputImg1[362],OutputImg1[361],OutputImg1[360],
                      OutputImg1[359],OutputImg1[358],OutputImg1[357],
                      OutputImg1[356],OutputImg1[355],OutputImg1[354],
                      OutputImg1[353],OutputImg1[352]}), .EN (nx23702), .F ({
                      ImgReg1IN_351,ImgReg1IN_350,ImgReg1IN_349,ImgReg1IN_348,
                      ImgReg1IN_347,ImgReg1IN_346,ImgReg1IN_345,ImgReg1IN_344,
                      ImgReg1IN_343,ImgReg1IN_342,ImgReg1IN_341,ImgReg1IN_340,
                      ImgReg1IN_339,ImgReg1IN_338,ImgReg1IN_337,ImgReg1IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState2L (.D ({OutputImg2[367],OutputImg2[366],
                      OutputImg2[365],OutputImg2[364],OutputImg2[363],
                      OutputImg2[362],OutputImg2[361],OutputImg2[360],
                      OutputImg2[359],OutputImg2[358],OutputImg2[357],
                      OutputImg2[356],OutputImg2[355],OutputImg2[354],
                      OutputImg2[353],OutputImg2[352]}), .EN (nx23702), .F ({
                      ImgReg2IN_351,ImgReg2IN_350,ImgReg2IN_349,ImgReg2IN_348,
                      ImgReg2IN_347,ImgReg2IN_346,ImgReg2IN_345,ImgReg2IN_344,
                      ImgReg2IN_343,ImgReg2IN_342,ImgReg2IN_341,ImgReg2IN_340,
                      ImgReg2IN_339,ImgReg2IN_338,ImgReg2IN_337,ImgReg2IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState3L (.D ({OutputImg3[367],OutputImg3[366],
                      OutputImg3[365],OutputImg3[364],OutputImg3[363],
                      OutputImg3[362],OutputImg3[361],OutputImg3[360],
                      OutputImg3[359],OutputImg3[358],OutputImg3[357],
                      OutputImg3[356],OutputImg3[355],OutputImg3[354],
                      OutputImg3[353],OutputImg3[352]}), .EN (nx23702), .F ({
                      ImgReg3IN_351,ImgReg3IN_350,ImgReg3IN_349,ImgReg3IN_348,
                      ImgReg3IN_347,ImgReg3IN_346,ImgReg3IN_345,ImgReg3IN_344,
                      ImgReg3IN_343,ImgReg3IN_342,ImgReg3IN_341,ImgReg3IN_340,
                      ImgReg3IN_339,ImgReg3IN_338,ImgReg3IN_337,ImgReg3IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState4L (.D ({OutputImg4[367],OutputImg4[366],
                      OutputImg4[365],OutputImg4[364],OutputImg4[363],
                      OutputImg4[362],OutputImg4[361],OutputImg4[360],
                      OutputImg4[359],OutputImg4[358],OutputImg4[357],
                      OutputImg4[356],OutputImg4[355],OutputImg4[354],
                      OutputImg4[353],OutputImg4[352]}), .EN (nx23702), .F ({
                      ImgReg4IN_351,ImgReg4IN_350,ImgReg4IN_349,ImgReg4IN_348,
                      ImgReg4IN_347,ImgReg4IN_346,ImgReg4IN_345,ImgReg4IN_344,
                      ImgReg4IN_343,ImgReg4IN_342,ImgReg4IN_341,ImgReg4IN_340,
                      ImgReg4IN_339,ImgReg4IN_338,ImgReg4IN_337,ImgReg4IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState5L (.D ({OutputImg5[367],OutputImg5[366],
                      OutputImg5[365],OutputImg5[364],OutputImg5[363],
                      OutputImg5[362],OutputImg5[361],OutputImg5[360],
                      OutputImg5[359],OutputImg5[358],OutputImg5[357],
                      OutputImg5[356],OutputImg5[355],OutputImg5[354],
                      OutputImg5[353],OutputImg5[352]}), .EN (nx23702), .F ({
                      ImgReg5IN_351,ImgReg5IN_350,ImgReg5IN_349,ImgReg5IN_348,
                      ImgReg5IN_347,ImgReg5IN_346,ImgReg5IN_345,ImgReg5IN_344,
                      ImgReg5IN_343,ImgReg5IN_342,ImgReg5IN_341,ImgReg5IN_340,
                      ImgReg5IN_339,ImgReg5IN_338,ImgReg5IN_337,ImgReg5IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState0N (.D ({DATA[351],DATA[350],DATA[349],
                      DATA[348],DATA[347],DATA[346],DATA[345],DATA[344],
                      DATA[343],DATA[342],DATA[341],DATA[340],DATA[339],
                      DATA[338],DATA[337],DATA[336]}), .EN (nx23660), .F ({
                      ImgReg0IN_351,ImgReg0IN_350,ImgReg0IN_349,ImgReg0IN_348,
                      ImgReg0IN_347,ImgReg0IN_346,ImgReg0IN_345,ImgReg0IN_344,
                      ImgReg0IN_343,ImgReg0IN_342,ImgReg0IN_341,ImgReg0IN_340,
                      ImgReg0IN_339,ImgReg0IN_338,ImgReg0IN_337,ImgReg0IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState1N (.D ({DATA[351],DATA[350],DATA[349],
                      DATA[348],DATA[347],DATA[346],DATA[345],DATA[344],
                      DATA[343],DATA[342],DATA[341],DATA[340],DATA[339],
                      DATA[338],DATA[337],DATA[336]}), .EN (nx23648), .F ({
                      ImgReg1IN_351,ImgReg1IN_350,ImgReg1IN_349,ImgReg1IN_348,
                      ImgReg1IN_347,ImgReg1IN_346,ImgReg1IN_345,ImgReg1IN_344,
                      ImgReg1IN_343,ImgReg1IN_342,ImgReg1IN_341,ImgReg1IN_340,
                      ImgReg1IN_339,ImgReg1IN_338,ImgReg1IN_337,ImgReg1IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState2N (.D ({DATA[351],DATA[350],DATA[349],
                      DATA[348],DATA[347],DATA[346],DATA[345],DATA[344],
                      DATA[343],DATA[342],DATA[341],DATA[340],DATA[339],
                      DATA[338],DATA[337],DATA[336]}), .EN (nx23636), .F ({
                      ImgReg2IN_351,ImgReg2IN_350,ImgReg2IN_349,ImgReg2IN_348,
                      ImgReg2IN_347,ImgReg2IN_346,ImgReg2IN_345,ImgReg2IN_344,
                      ImgReg2IN_343,ImgReg2IN_342,ImgReg2IN_341,ImgReg2IN_340,
                      ImgReg2IN_339,ImgReg2IN_338,ImgReg2IN_337,ImgReg2IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState3N (.D ({DATA[351],DATA[350],DATA[349],
                      DATA[348],DATA[347],DATA[346],DATA[345],DATA[344],
                      DATA[343],DATA[342],DATA[341],DATA[340],DATA[339],
                      DATA[338],DATA[337],DATA[336]}), .EN (nx23624), .F ({
                      ImgReg3IN_351,ImgReg3IN_350,ImgReg3IN_349,ImgReg3IN_348,
                      ImgReg3IN_347,ImgReg3IN_346,ImgReg3IN_345,ImgReg3IN_344,
                      ImgReg3IN_343,ImgReg3IN_342,ImgReg3IN_341,ImgReg3IN_340,
                      ImgReg3IN_339,ImgReg3IN_338,ImgReg3IN_337,ImgReg3IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState4N (.D ({DATA[351],DATA[350],DATA[349],
                      DATA[348],DATA[347],DATA[346],DATA[345],DATA[344],
                      DATA[343],DATA[342],DATA[341],DATA[340],DATA[339],
                      DATA[338],DATA[337],DATA[336]}), .EN (nx23612), .F ({
                      ImgReg4IN_351,ImgReg4IN_350,ImgReg4IN_349,ImgReg4IN_348,
                      ImgReg4IN_347,ImgReg4IN_346,ImgReg4IN_345,ImgReg4IN_344,
                      ImgReg4IN_343,ImgReg4IN_342,ImgReg4IN_341,ImgReg4IN_340,
                      ImgReg4IN_339,ImgReg4IN_338,ImgReg4IN_337,ImgReg4IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState5N (.D ({DATA[351],DATA[350],DATA[349],
                      DATA[348],DATA[347],DATA[346],DATA[345],DATA[344],
                      DATA[343],DATA[342],DATA[341],DATA[340],DATA[339],
                      DATA[338],DATA[337],DATA[336]}), .EN (nx23600), .F ({
                      ImgReg5IN_351,ImgReg5IN_350,ImgReg5IN_349,ImgReg5IN_348,
                      ImgReg5IN_347,ImgReg5IN_346,ImgReg5IN_345,ImgReg5IN_344,
                      ImgReg5IN_343,ImgReg5IN_342,ImgReg5IN_341,ImgReg5IN_340,
                      ImgReg5IN_339,ImgReg5IN_338,ImgReg5IN_337,ImgReg5IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState0U (.D ({OutputImg1[351],OutputImg1[350],
                      OutputImg1[349],OutputImg1[348],OutputImg1[347],
                      OutputImg1[346],OutputImg1[345],OutputImg1[344],
                      OutputImg1[343],OutputImg1[342],OutputImg1[341],
                      OutputImg1[340],OutputImg1[339],OutputImg1[338],
                      OutputImg1[337],OutputImg1[336]}), .EN (nx23816), .F ({
                      ImgReg0IN_351,ImgReg0IN_350,ImgReg0IN_349,ImgReg0IN_348,
                      ImgReg0IN_347,ImgReg0IN_346,ImgReg0IN_345,ImgReg0IN_344,
                      ImgReg0IN_343,ImgReg0IN_342,ImgReg0IN_341,ImgReg0IN_340,
                      ImgReg0IN_339,ImgReg0IN_338,ImgReg0IN_337,ImgReg0IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState1U (.D ({OutputImg2[351],OutputImg2[350],
                      OutputImg2[349],OutputImg2[348],OutputImg2[347],
                      OutputImg2[346],OutputImg2[345],OutputImg2[344],
                      OutputImg2[343],OutputImg2[342],OutputImg2[341],
                      OutputImg2[340],OutputImg2[339],OutputImg2[338],
                      OutputImg2[337],OutputImg2[336]}), .EN (nx23816), .F ({
                      ImgReg1IN_351,ImgReg1IN_350,ImgReg1IN_349,ImgReg1IN_348,
                      ImgReg1IN_347,ImgReg1IN_346,ImgReg1IN_345,ImgReg1IN_344,
                      ImgReg1IN_343,ImgReg1IN_342,ImgReg1IN_341,ImgReg1IN_340,
                      ImgReg1IN_339,ImgReg1IN_338,ImgReg1IN_337,ImgReg1IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState2U (.D ({OutputImg3[351],OutputImg3[350],
                      OutputImg3[349],OutputImg3[348],OutputImg3[347],
                      OutputImg3[346],OutputImg3[345],OutputImg3[344],
                      OutputImg3[343],OutputImg3[342],OutputImg3[341],
                      OutputImg3[340],OutputImg3[339],OutputImg3[338],
                      OutputImg3[337],OutputImg3[336]}), .EN (nx23816), .F ({
                      ImgReg2IN_351,ImgReg2IN_350,ImgReg2IN_349,ImgReg2IN_348,
                      ImgReg2IN_347,ImgReg2IN_346,ImgReg2IN_345,ImgReg2IN_344,
                      ImgReg2IN_343,ImgReg2IN_342,ImgReg2IN_341,ImgReg2IN_340,
                      ImgReg2IN_339,ImgReg2IN_338,ImgReg2IN_337,ImgReg2IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState3U (.D ({OutputImg4[351],OutputImg4[350],
                      OutputImg4[349],OutputImg4[348],OutputImg4[347],
                      OutputImg4[346],OutputImg4[345],OutputImg4[344],
                      OutputImg4[343],OutputImg4[342],OutputImg4[341],
                      OutputImg4[340],OutputImg4[339],OutputImg4[338],
                      OutputImg4[337],OutputImg4[336]}), .EN (nx23816), .F ({
                      ImgReg3IN_351,ImgReg3IN_350,ImgReg3IN_349,ImgReg3IN_348,
                      ImgReg3IN_347,ImgReg3IN_346,ImgReg3IN_345,ImgReg3IN_344,
                      ImgReg3IN_343,ImgReg3IN_342,ImgReg3IN_341,ImgReg3IN_340,
                      ImgReg3IN_339,ImgReg3IN_338,ImgReg3IN_337,ImgReg3IN_336})
                      ) ;
    triStateBuffer_16 loop3_21_TriState4U (.D ({OutputImg5[351],OutputImg5[350],
                      OutputImg5[349],OutputImg5[348],OutputImg5[347],
                      OutputImg5[346],OutputImg5[345],OutputImg5[344],
                      OutputImg5[343],OutputImg5[342],OutputImg5[341],
                      OutputImg5[340],OutputImg5[339],OutputImg5[338],
                      OutputImg5[337],OutputImg5[336]}), .EN (nx23816), .F ({
                      ImgReg4IN_351,ImgReg4IN_350,ImgReg4IN_349,ImgReg4IN_348,
                      ImgReg4IN_347,ImgReg4IN_346,ImgReg4IN_345,ImgReg4IN_344,
                      ImgReg4IN_343,ImgReg4IN_342,ImgReg4IN_341,ImgReg4IN_340,
                      ImgReg4IN_339,ImgReg4IN_338,ImgReg4IN_337,ImgReg4IN_336})
                      ) ;
    nBitRegister_16 loop3_21_reg1 (.D ({ImgReg0IN_351,ImgReg0IN_350,
                    ImgReg0IN_349,ImgReg0IN_348,ImgReg0IN_347,ImgReg0IN_346,
                    ImgReg0IN_345,ImgReg0IN_344,ImgReg0IN_343,ImgReg0IN_342,
                    ImgReg0IN_341,ImgReg0IN_340,ImgReg0IN_339,ImgReg0IN_338,
                    ImgReg0IN_337,ImgReg0IN_336}), .CLK (nx23954), .RST (RST), .EN (
                    nx23724), .Q ({OutputImg0[351],OutputImg0[350],
                    OutputImg0[349],OutputImg0[348],OutputImg0[347],
                    OutputImg0[346],OutputImg0[345],OutputImg0[344],
                    OutputImg0[343],OutputImg0[342],OutputImg0[341],
                    OutputImg0[340],OutputImg0[339],OutputImg0[338],
                    OutputImg0[337],OutputImg0[336]})) ;
    nBitRegister_16 loop3_21_reg2 (.D ({ImgReg1IN_351,ImgReg1IN_350,
                    ImgReg1IN_349,ImgReg1IN_348,ImgReg1IN_347,ImgReg1IN_346,
                    ImgReg1IN_345,ImgReg1IN_344,ImgReg1IN_343,ImgReg1IN_342,
                    ImgReg1IN_341,ImgReg1IN_340,ImgReg1IN_339,ImgReg1IN_338,
                    ImgReg1IN_337,ImgReg1IN_336}), .CLK (nx23956), .RST (RST), .EN (
                    nx23734), .Q ({OutputImg1[351],OutputImg1[350],
                    OutputImg1[349],OutputImg1[348],OutputImg1[347],
                    OutputImg1[346],OutputImg1[345],OutputImg1[344],
                    OutputImg1[343],OutputImg1[342],OutputImg1[341],
                    OutputImg1[340],OutputImg1[339],OutputImg1[338],
                    OutputImg1[337],OutputImg1[336]})) ;
    nBitRegister_16 loop3_21_reg3 (.D ({ImgReg2IN_351,ImgReg2IN_350,
                    ImgReg2IN_349,ImgReg2IN_348,ImgReg2IN_347,ImgReg2IN_346,
                    ImgReg2IN_345,ImgReg2IN_344,ImgReg2IN_343,ImgReg2IN_342,
                    ImgReg2IN_341,ImgReg2IN_340,ImgReg2IN_339,ImgReg2IN_338,
                    ImgReg2IN_337,ImgReg2IN_336}), .CLK (nx23956), .RST (RST), .EN (
                    nx23744), .Q ({OutputImg2[351],OutputImg2[350],
                    OutputImg2[349],OutputImg2[348],OutputImg2[347],
                    OutputImg2[346],OutputImg2[345],OutputImg2[344],
                    OutputImg2[343],OutputImg2[342],OutputImg2[341],
                    OutputImg2[340],OutputImg2[339],OutputImg2[338],
                    OutputImg2[337],OutputImg2[336]})) ;
    nBitRegister_16 loop3_21_reg4 (.D ({ImgReg3IN_351,ImgReg3IN_350,
                    ImgReg3IN_349,ImgReg3IN_348,ImgReg3IN_347,ImgReg3IN_346,
                    ImgReg3IN_345,ImgReg3IN_344,ImgReg3IN_343,ImgReg3IN_342,
                    ImgReg3IN_341,ImgReg3IN_340,ImgReg3IN_339,ImgReg3IN_338,
                    ImgReg3IN_337,ImgReg3IN_336}), .CLK (nx23958), .RST (RST), .EN (
                    nx23754), .Q ({OutputImg3[351],OutputImg3[350],
                    OutputImg3[349],OutputImg3[348],OutputImg3[347],
                    OutputImg3[346],OutputImg3[345],OutputImg3[344],
                    OutputImg3[343],OutputImg3[342],OutputImg3[341],
                    OutputImg3[340],OutputImg3[339],OutputImg3[338],
                    OutputImg3[337],OutputImg3[336]})) ;
    nBitRegister_16 loop3_21_reg5 (.D ({ImgReg4IN_351,ImgReg4IN_350,
                    ImgReg4IN_349,ImgReg4IN_348,ImgReg4IN_347,ImgReg4IN_346,
                    ImgReg4IN_345,ImgReg4IN_344,ImgReg4IN_343,ImgReg4IN_342,
                    ImgReg4IN_341,ImgReg4IN_340,ImgReg4IN_339,ImgReg4IN_338,
                    ImgReg4IN_337,ImgReg4IN_336}), .CLK (nx23958), .RST (RST), .EN (
                    nx23764), .Q ({OutputImg4[351],OutputImg4[350],
                    OutputImg4[349],OutputImg4[348],OutputImg4[347],
                    OutputImg4[346],OutputImg4[345],OutputImg4[344],
                    OutputImg4[343],OutputImg4[342],OutputImg4[341],
                    OutputImg4[340],OutputImg4[339],OutputImg4[338],
                    OutputImg4[337],OutputImg4[336]})) ;
    nBitRegister_16 loop3_21_reg6 (.D ({ImgReg5IN_351,ImgReg5IN_350,
                    ImgReg5IN_349,ImgReg5IN_348,ImgReg5IN_347,ImgReg5IN_346,
                    ImgReg5IN_345,ImgReg5IN_344,ImgReg5IN_343,ImgReg5IN_342,
                    ImgReg5IN_341,ImgReg5IN_340,ImgReg5IN_339,ImgReg5IN_338,
                    ImgReg5IN_337,ImgReg5IN_336}), .CLK (nx23960), .RST (RST), .EN (
                    nx23774), .Q ({OutputImg5[351],OutputImg5[350],
                    OutputImg5[349],OutputImg5[348],OutputImg5[347],
                    OutputImg5[346],OutputImg5[345],OutputImg5[344],
                    OutputImg5[343],OutputImg5[342],OutputImg5[341],
                    OutputImg5[340],OutputImg5[339],OutputImg5[338],
                    OutputImg5[337],OutputImg5[336]})) ;
    triStateBuffer_16 loop3_22_TriState0L (.D ({OutputImg0[383],OutputImg0[382],
                      OutputImg0[381],OutputImg0[380],OutputImg0[379],
                      OutputImg0[378],OutputImg0[377],OutputImg0[376],
                      OutputImg0[375],OutputImg0[374],OutputImg0[373],
                      OutputImg0[372],OutputImg0[371],OutputImg0[370],
                      OutputImg0[369],OutputImg0[368]}), .EN (nx23702), .F ({
                      ImgReg0IN_367,ImgReg0IN_366,ImgReg0IN_365,ImgReg0IN_364,
                      ImgReg0IN_363,ImgReg0IN_362,ImgReg0IN_361,ImgReg0IN_360,
                      ImgReg0IN_359,ImgReg0IN_358,ImgReg0IN_357,ImgReg0IN_356,
                      ImgReg0IN_355,ImgReg0IN_354,ImgReg0IN_353,ImgReg0IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState1L (.D ({OutputImg1[383],OutputImg1[382],
                      OutputImg1[381],OutputImg1[380],OutputImg1[379],
                      OutputImg1[378],OutputImg1[377],OutputImg1[376],
                      OutputImg1[375],OutputImg1[374],OutputImg1[373],
                      OutputImg1[372],OutputImg1[371],OutputImg1[370],
                      OutputImg1[369],OutputImg1[368]}), .EN (nx23704), .F ({
                      ImgReg1IN_367,ImgReg1IN_366,ImgReg1IN_365,ImgReg1IN_364,
                      ImgReg1IN_363,ImgReg1IN_362,ImgReg1IN_361,ImgReg1IN_360,
                      ImgReg1IN_359,ImgReg1IN_358,ImgReg1IN_357,ImgReg1IN_356,
                      ImgReg1IN_355,ImgReg1IN_354,ImgReg1IN_353,ImgReg1IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState2L (.D ({OutputImg2[383],OutputImg2[382],
                      OutputImg2[381],OutputImg2[380],OutputImg2[379],
                      OutputImg2[378],OutputImg2[377],OutputImg2[376],
                      OutputImg2[375],OutputImg2[374],OutputImg2[373],
                      OutputImg2[372],OutputImg2[371],OutputImg2[370],
                      OutputImg2[369],OutputImg2[368]}), .EN (nx23704), .F ({
                      ImgReg2IN_367,ImgReg2IN_366,ImgReg2IN_365,ImgReg2IN_364,
                      ImgReg2IN_363,ImgReg2IN_362,ImgReg2IN_361,ImgReg2IN_360,
                      ImgReg2IN_359,ImgReg2IN_358,ImgReg2IN_357,ImgReg2IN_356,
                      ImgReg2IN_355,ImgReg2IN_354,ImgReg2IN_353,ImgReg2IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState3L (.D ({OutputImg3[383],OutputImg3[382],
                      OutputImg3[381],OutputImg3[380],OutputImg3[379],
                      OutputImg3[378],OutputImg3[377],OutputImg3[376],
                      OutputImg3[375],OutputImg3[374],OutputImg3[373],
                      OutputImg3[372],OutputImg3[371],OutputImg3[370],
                      OutputImg3[369],OutputImg3[368]}), .EN (nx23704), .F ({
                      ImgReg3IN_367,ImgReg3IN_366,ImgReg3IN_365,ImgReg3IN_364,
                      ImgReg3IN_363,ImgReg3IN_362,ImgReg3IN_361,ImgReg3IN_360,
                      ImgReg3IN_359,ImgReg3IN_358,ImgReg3IN_357,ImgReg3IN_356,
                      ImgReg3IN_355,ImgReg3IN_354,ImgReg3IN_353,ImgReg3IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState4L (.D ({OutputImg4[383],OutputImg4[382],
                      OutputImg4[381],OutputImg4[380],OutputImg4[379],
                      OutputImg4[378],OutputImg4[377],OutputImg4[376],
                      OutputImg4[375],OutputImg4[374],OutputImg4[373],
                      OutputImg4[372],OutputImg4[371],OutputImg4[370],
                      OutputImg4[369],OutputImg4[368]}), .EN (nx23704), .F ({
                      ImgReg4IN_367,ImgReg4IN_366,ImgReg4IN_365,ImgReg4IN_364,
                      ImgReg4IN_363,ImgReg4IN_362,ImgReg4IN_361,ImgReg4IN_360,
                      ImgReg4IN_359,ImgReg4IN_358,ImgReg4IN_357,ImgReg4IN_356,
                      ImgReg4IN_355,ImgReg4IN_354,ImgReg4IN_353,ImgReg4IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState5L (.D ({OutputImg5[383],OutputImg5[382],
                      OutputImg5[381],OutputImg5[380],OutputImg5[379],
                      OutputImg5[378],OutputImg5[377],OutputImg5[376],
                      OutputImg5[375],OutputImg5[374],OutputImg5[373],
                      OutputImg5[372],OutputImg5[371],OutputImg5[370],
                      OutputImg5[369],OutputImg5[368]}), .EN (nx23704), .F ({
                      ImgReg5IN_367,ImgReg5IN_366,ImgReg5IN_365,ImgReg5IN_364,
                      ImgReg5IN_363,ImgReg5IN_362,ImgReg5IN_361,ImgReg5IN_360,
                      ImgReg5IN_359,ImgReg5IN_358,ImgReg5IN_357,ImgReg5IN_356,
                      ImgReg5IN_355,ImgReg5IN_354,ImgReg5IN_353,ImgReg5IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState0N (.D ({DATA[367],DATA[366],DATA[365],
                      DATA[364],DATA[363],DATA[362],DATA[361],DATA[360],
                      DATA[359],DATA[358],DATA[357],DATA[356],DATA[355],
                      DATA[354],DATA[353],DATA[352]}), .EN (nx23660), .F ({
                      ImgReg0IN_367,ImgReg0IN_366,ImgReg0IN_365,ImgReg0IN_364,
                      ImgReg0IN_363,ImgReg0IN_362,ImgReg0IN_361,ImgReg0IN_360,
                      ImgReg0IN_359,ImgReg0IN_358,ImgReg0IN_357,ImgReg0IN_356,
                      ImgReg0IN_355,ImgReg0IN_354,ImgReg0IN_353,ImgReg0IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState1N (.D ({DATA[367],DATA[366],DATA[365],
                      DATA[364],DATA[363],DATA[362],DATA[361],DATA[360],
                      DATA[359],DATA[358],DATA[357],DATA[356],DATA[355],
                      DATA[354],DATA[353],DATA[352]}), .EN (nx23648), .F ({
                      ImgReg1IN_367,ImgReg1IN_366,ImgReg1IN_365,ImgReg1IN_364,
                      ImgReg1IN_363,ImgReg1IN_362,ImgReg1IN_361,ImgReg1IN_360,
                      ImgReg1IN_359,ImgReg1IN_358,ImgReg1IN_357,ImgReg1IN_356,
                      ImgReg1IN_355,ImgReg1IN_354,ImgReg1IN_353,ImgReg1IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState2N (.D ({DATA[367],DATA[366],DATA[365],
                      DATA[364],DATA[363],DATA[362],DATA[361],DATA[360],
                      DATA[359],DATA[358],DATA[357],DATA[356],DATA[355],
                      DATA[354],DATA[353],DATA[352]}), .EN (nx23636), .F ({
                      ImgReg2IN_367,ImgReg2IN_366,ImgReg2IN_365,ImgReg2IN_364,
                      ImgReg2IN_363,ImgReg2IN_362,ImgReg2IN_361,ImgReg2IN_360,
                      ImgReg2IN_359,ImgReg2IN_358,ImgReg2IN_357,ImgReg2IN_356,
                      ImgReg2IN_355,ImgReg2IN_354,ImgReg2IN_353,ImgReg2IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState3N (.D ({DATA[367],DATA[366],DATA[365],
                      DATA[364],DATA[363],DATA[362],DATA[361],DATA[360],
                      DATA[359],DATA[358],DATA[357],DATA[356],DATA[355],
                      DATA[354],DATA[353],DATA[352]}), .EN (nx23624), .F ({
                      ImgReg3IN_367,ImgReg3IN_366,ImgReg3IN_365,ImgReg3IN_364,
                      ImgReg3IN_363,ImgReg3IN_362,ImgReg3IN_361,ImgReg3IN_360,
                      ImgReg3IN_359,ImgReg3IN_358,ImgReg3IN_357,ImgReg3IN_356,
                      ImgReg3IN_355,ImgReg3IN_354,ImgReg3IN_353,ImgReg3IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState4N (.D ({DATA[367],DATA[366],DATA[365],
                      DATA[364],DATA[363],DATA[362],DATA[361],DATA[360],
                      DATA[359],DATA[358],DATA[357],DATA[356],DATA[355],
                      DATA[354],DATA[353],DATA[352]}), .EN (nx23612), .F ({
                      ImgReg4IN_367,ImgReg4IN_366,ImgReg4IN_365,ImgReg4IN_364,
                      ImgReg4IN_363,ImgReg4IN_362,ImgReg4IN_361,ImgReg4IN_360,
                      ImgReg4IN_359,ImgReg4IN_358,ImgReg4IN_357,ImgReg4IN_356,
                      ImgReg4IN_355,ImgReg4IN_354,ImgReg4IN_353,ImgReg4IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState5N (.D ({DATA[367],DATA[366],DATA[365],
                      DATA[364],DATA[363],DATA[362],DATA[361],DATA[360],
                      DATA[359],DATA[358],DATA[357],DATA[356],DATA[355],
                      DATA[354],DATA[353],DATA[352]}), .EN (nx23600), .F ({
                      ImgReg5IN_367,ImgReg5IN_366,ImgReg5IN_365,ImgReg5IN_364,
                      ImgReg5IN_363,ImgReg5IN_362,ImgReg5IN_361,ImgReg5IN_360,
                      ImgReg5IN_359,ImgReg5IN_358,ImgReg5IN_357,ImgReg5IN_356,
                      ImgReg5IN_355,ImgReg5IN_354,ImgReg5IN_353,ImgReg5IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState0U (.D ({OutputImg1[367],OutputImg1[366],
                      OutputImg1[365],OutputImg1[364],OutputImg1[363],
                      OutputImg1[362],OutputImg1[361],OutputImg1[360],
                      OutputImg1[359],OutputImg1[358],OutputImg1[357],
                      OutputImg1[356],OutputImg1[355],OutputImg1[354],
                      OutputImg1[353],OutputImg1[352]}), .EN (nx23816), .F ({
                      ImgReg0IN_367,ImgReg0IN_366,ImgReg0IN_365,ImgReg0IN_364,
                      ImgReg0IN_363,ImgReg0IN_362,ImgReg0IN_361,ImgReg0IN_360,
                      ImgReg0IN_359,ImgReg0IN_358,ImgReg0IN_357,ImgReg0IN_356,
                      ImgReg0IN_355,ImgReg0IN_354,ImgReg0IN_353,ImgReg0IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState1U (.D ({OutputImg2[367],OutputImg2[366],
                      OutputImg2[365],OutputImg2[364],OutputImg2[363],
                      OutputImg2[362],OutputImg2[361],OutputImg2[360],
                      OutputImg2[359],OutputImg2[358],OutputImg2[357],
                      OutputImg2[356],OutputImg2[355],OutputImg2[354],
                      OutputImg2[353],OutputImg2[352]}), .EN (nx23816), .F ({
                      ImgReg1IN_367,ImgReg1IN_366,ImgReg1IN_365,ImgReg1IN_364,
                      ImgReg1IN_363,ImgReg1IN_362,ImgReg1IN_361,ImgReg1IN_360,
                      ImgReg1IN_359,ImgReg1IN_358,ImgReg1IN_357,ImgReg1IN_356,
                      ImgReg1IN_355,ImgReg1IN_354,ImgReg1IN_353,ImgReg1IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState2U (.D ({OutputImg3[367],OutputImg3[366],
                      OutputImg3[365],OutputImg3[364],OutputImg3[363],
                      OutputImg3[362],OutputImg3[361],OutputImg3[360],
                      OutputImg3[359],OutputImg3[358],OutputImg3[357],
                      OutputImg3[356],OutputImg3[355],OutputImg3[354],
                      OutputImg3[353],OutputImg3[352]}), .EN (nx23818), .F ({
                      ImgReg2IN_367,ImgReg2IN_366,ImgReg2IN_365,ImgReg2IN_364,
                      ImgReg2IN_363,ImgReg2IN_362,ImgReg2IN_361,ImgReg2IN_360,
                      ImgReg2IN_359,ImgReg2IN_358,ImgReg2IN_357,ImgReg2IN_356,
                      ImgReg2IN_355,ImgReg2IN_354,ImgReg2IN_353,ImgReg2IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState3U (.D ({OutputImg4[367],OutputImg4[366],
                      OutputImg4[365],OutputImg4[364],OutputImg4[363],
                      OutputImg4[362],OutputImg4[361],OutputImg4[360],
                      OutputImg4[359],OutputImg4[358],OutputImg4[357],
                      OutputImg4[356],OutputImg4[355],OutputImg4[354],
                      OutputImg4[353],OutputImg4[352]}), .EN (nx23818), .F ({
                      ImgReg3IN_367,ImgReg3IN_366,ImgReg3IN_365,ImgReg3IN_364,
                      ImgReg3IN_363,ImgReg3IN_362,ImgReg3IN_361,ImgReg3IN_360,
                      ImgReg3IN_359,ImgReg3IN_358,ImgReg3IN_357,ImgReg3IN_356,
                      ImgReg3IN_355,ImgReg3IN_354,ImgReg3IN_353,ImgReg3IN_352})
                      ) ;
    triStateBuffer_16 loop3_22_TriState4U (.D ({OutputImg5[367],OutputImg5[366],
                      OutputImg5[365],OutputImg5[364],OutputImg5[363],
                      OutputImg5[362],OutputImg5[361],OutputImg5[360],
                      OutputImg5[359],OutputImg5[358],OutputImg5[357],
                      OutputImg5[356],OutputImg5[355],OutputImg5[354],
                      OutputImg5[353],OutputImg5[352]}), .EN (nx23818), .F ({
                      ImgReg4IN_367,ImgReg4IN_366,ImgReg4IN_365,ImgReg4IN_364,
                      ImgReg4IN_363,ImgReg4IN_362,ImgReg4IN_361,ImgReg4IN_360,
                      ImgReg4IN_359,ImgReg4IN_358,ImgReg4IN_357,ImgReg4IN_356,
                      ImgReg4IN_355,ImgReg4IN_354,ImgReg4IN_353,ImgReg4IN_352})
                      ) ;
    nBitRegister_16 loop3_22_reg1 (.D ({ImgReg0IN_367,ImgReg0IN_366,
                    ImgReg0IN_365,ImgReg0IN_364,ImgReg0IN_363,ImgReg0IN_362,
                    ImgReg0IN_361,ImgReg0IN_360,ImgReg0IN_359,ImgReg0IN_358,
                    ImgReg0IN_357,ImgReg0IN_356,ImgReg0IN_355,ImgReg0IN_354,
                    ImgReg0IN_353,ImgReg0IN_352}), .CLK (nx23960), .RST (RST), .EN (
                    nx23724), .Q ({OutputImg0[367],OutputImg0[366],
                    OutputImg0[365],OutputImg0[364],OutputImg0[363],
                    OutputImg0[362],OutputImg0[361],OutputImg0[360],
                    OutputImg0[359],OutputImg0[358],OutputImg0[357],
                    OutputImg0[356],OutputImg0[355],OutputImg0[354],
                    OutputImg0[353],OutputImg0[352]})) ;
    nBitRegister_16 loop3_22_reg2 (.D ({ImgReg1IN_367,ImgReg1IN_366,
                    ImgReg1IN_365,ImgReg1IN_364,ImgReg1IN_363,ImgReg1IN_362,
                    ImgReg1IN_361,ImgReg1IN_360,ImgReg1IN_359,ImgReg1IN_358,
                    ImgReg1IN_357,ImgReg1IN_356,ImgReg1IN_355,ImgReg1IN_354,
                    ImgReg1IN_353,ImgReg1IN_352}), .CLK (nx23962), .RST (RST), .EN (
                    nx23734), .Q ({OutputImg1[367],OutputImg1[366],
                    OutputImg1[365],OutputImg1[364],OutputImg1[363],
                    OutputImg1[362],OutputImg1[361],OutputImg1[360],
                    OutputImg1[359],OutputImg1[358],OutputImg1[357],
                    OutputImg1[356],OutputImg1[355],OutputImg1[354],
                    OutputImg1[353],OutputImg1[352]})) ;
    nBitRegister_16 loop3_22_reg3 (.D ({ImgReg2IN_367,ImgReg2IN_366,
                    ImgReg2IN_365,ImgReg2IN_364,ImgReg2IN_363,ImgReg2IN_362,
                    ImgReg2IN_361,ImgReg2IN_360,ImgReg2IN_359,ImgReg2IN_358,
                    ImgReg2IN_357,ImgReg2IN_356,ImgReg2IN_355,ImgReg2IN_354,
                    ImgReg2IN_353,ImgReg2IN_352}), .CLK (nx23962), .RST (RST), .EN (
                    nx23744), .Q ({OutputImg2[367],OutputImg2[366],
                    OutputImg2[365],OutputImg2[364],OutputImg2[363],
                    OutputImg2[362],OutputImg2[361],OutputImg2[360],
                    OutputImg2[359],OutputImg2[358],OutputImg2[357],
                    OutputImg2[356],OutputImg2[355],OutputImg2[354],
                    OutputImg2[353],OutputImg2[352]})) ;
    nBitRegister_16 loop3_22_reg4 (.D ({ImgReg3IN_367,ImgReg3IN_366,
                    ImgReg3IN_365,ImgReg3IN_364,ImgReg3IN_363,ImgReg3IN_362,
                    ImgReg3IN_361,ImgReg3IN_360,ImgReg3IN_359,ImgReg3IN_358,
                    ImgReg3IN_357,ImgReg3IN_356,ImgReg3IN_355,ImgReg3IN_354,
                    ImgReg3IN_353,ImgReg3IN_352}), .CLK (nx23964), .RST (RST), .EN (
                    nx23754), .Q ({OutputImg3[367],OutputImg3[366],
                    OutputImg3[365],OutputImg3[364],OutputImg3[363],
                    OutputImg3[362],OutputImg3[361],OutputImg3[360],
                    OutputImg3[359],OutputImg3[358],OutputImg3[357],
                    OutputImg3[356],OutputImg3[355],OutputImg3[354],
                    OutputImg3[353],OutputImg3[352]})) ;
    nBitRegister_16 loop3_22_reg5 (.D ({ImgReg4IN_367,ImgReg4IN_366,
                    ImgReg4IN_365,ImgReg4IN_364,ImgReg4IN_363,ImgReg4IN_362,
                    ImgReg4IN_361,ImgReg4IN_360,ImgReg4IN_359,ImgReg4IN_358,
                    ImgReg4IN_357,ImgReg4IN_356,ImgReg4IN_355,ImgReg4IN_354,
                    ImgReg4IN_353,ImgReg4IN_352}), .CLK (nx23964), .RST (RST), .EN (
                    nx23764), .Q ({OutputImg4[367],OutputImg4[366],
                    OutputImg4[365],OutputImg4[364],OutputImg4[363],
                    OutputImg4[362],OutputImg4[361],OutputImg4[360],
                    OutputImg4[359],OutputImg4[358],OutputImg4[357],
                    OutputImg4[356],OutputImg4[355],OutputImg4[354],
                    OutputImg4[353],OutputImg4[352]})) ;
    nBitRegister_16 loop3_22_reg6 (.D ({ImgReg5IN_367,ImgReg5IN_366,
                    ImgReg5IN_365,ImgReg5IN_364,ImgReg5IN_363,ImgReg5IN_362,
                    ImgReg5IN_361,ImgReg5IN_360,ImgReg5IN_359,ImgReg5IN_358,
                    ImgReg5IN_357,ImgReg5IN_356,ImgReg5IN_355,ImgReg5IN_354,
                    ImgReg5IN_353,ImgReg5IN_352}), .CLK (nx23966), .RST (RST), .EN (
                    nx23774), .Q ({OutputImg5[367],OutputImg5[366],
                    OutputImg5[365],OutputImg5[364],OutputImg5[363],
                    OutputImg5[362],OutputImg5[361],OutputImg5[360],
                    OutputImg5[359],OutputImg5[358],OutputImg5[357],
                    OutputImg5[356],OutputImg5[355],OutputImg5[354],
                    OutputImg5[353],OutputImg5[352]})) ;
    triStateBuffer_16 loop3_23_TriState0L (.D ({OutputImg0[399],OutputImg0[398],
                      OutputImg0[397],OutputImg0[396],OutputImg0[395],
                      OutputImg0[394],OutputImg0[393],OutputImg0[392],
                      OutputImg0[391],OutputImg0[390],OutputImg0[389],
                      OutputImg0[388],OutputImg0[387],OutputImg0[386],
                      OutputImg0[385],OutputImg0[384]}), .EN (nx23704), .F ({
                      ImgReg0IN_383,ImgReg0IN_382,ImgReg0IN_381,ImgReg0IN_380,
                      ImgReg0IN_379,ImgReg0IN_378,ImgReg0IN_377,ImgReg0IN_376,
                      ImgReg0IN_375,ImgReg0IN_374,ImgReg0IN_373,ImgReg0IN_372,
                      ImgReg0IN_371,ImgReg0IN_370,ImgReg0IN_369,ImgReg0IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState1L (.D ({OutputImg1[399],OutputImg1[398],
                      OutputImg1[397],OutputImg1[396],OutputImg1[395],
                      OutputImg1[394],OutputImg1[393],OutputImg1[392],
                      OutputImg1[391],OutputImg1[390],OutputImg1[389],
                      OutputImg1[388],OutputImg1[387],OutputImg1[386],
                      OutputImg1[385],OutputImg1[384]}), .EN (nx23704), .F ({
                      ImgReg1IN_383,ImgReg1IN_382,ImgReg1IN_381,ImgReg1IN_380,
                      ImgReg1IN_379,ImgReg1IN_378,ImgReg1IN_377,ImgReg1IN_376,
                      ImgReg1IN_375,ImgReg1IN_374,ImgReg1IN_373,ImgReg1IN_372,
                      ImgReg1IN_371,ImgReg1IN_370,ImgReg1IN_369,ImgReg1IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState2L (.D ({OutputImg2[399],OutputImg2[398],
                      OutputImg2[397],OutputImg2[396],OutputImg2[395],
                      OutputImg2[394],OutputImg2[393],OutputImg2[392],
                      OutputImg2[391],OutputImg2[390],OutputImg2[389],
                      OutputImg2[388],OutputImg2[387],OutputImg2[386],
                      OutputImg2[385],OutputImg2[384]}), .EN (nx23706), .F ({
                      ImgReg2IN_383,ImgReg2IN_382,ImgReg2IN_381,ImgReg2IN_380,
                      ImgReg2IN_379,ImgReg2IN_378,ImgReg2IN_377,ImgReg2IN_376,
                      ImgReg2IN_375,ImgReg2IN_374,ImgReg2IN_373,ImgReg2IN_372,
                      ImgReg2IN_371,ImgReg2IN_370,ImgReg2IN_369,ImgReg2IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState3L (.D ({OutputImg3[399],OutputImg3[398],
                      OutputImg3[397],OutputImg3[396],OutputImg3[395],
                      OutputImg3[394],OutputImg3[393],OutputImg3[392],
                      OutputImg3[391],OutputImg3[390],OutputImg3[389],
                      OutputImg3[388],OutputImg3[387],OutputImg3[386],
                      OutputImg3[385],OutputImg3[384]}), .EN (nx23706), .F ({
                      ImgReg3IN_383,ImgReg3IN_382,ImgReg3IN_381,ImgReg3IN_380,
                      ImgReg3IN_379,ImgReg3IN_378,ImgReg3IN_377,ImgReg3IN_376,
                      ImgReg3IN_375,ImgReg3IN_374,ImgReg3IN_373,ImgReg3IN_372,
                      ImgReg3IN_371,ImgReg3IN_370,ImgReg3IN_369,ImgReg3IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState4L (.D ({OutputImg4[399],OutputImg4[398],
                      OutputImg4[397],OutputImg4[396],OutputImg4[395],
                      OutputImg4[394],OutputImg4[393],OutputImg4[392],
                      OutputImg4[391],OutputImg4[390],OutputImg4[389],
                      OutputImg4[388],OutputImg4[387],OutputImg4[386],
                      OutputImg4[385],OutputImg4[384]}), .EN (nx23706), .F ({
                      ImgReg4IN_383,ImgReg4IN_382,ImgReg4IN_381,ImgReg4IN_380,
                      ImgReg4IN_379,ImgReg4IN_378,ImgReg4IN_377,ImgReg4IN_376,
                      ImgReg4IN_375,ImgReg4IN_374,ImgReg4IN_373,ImgReg4IN_372,
                      ImgReg4IN_371,ImgReg4IN_370,ImgReg4IN_369,ImgReg4IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState5L (.D ({OutputImg5[399],OutputImg5[398],
                      OutputImg5[397],OutputImg5[396],OutputImg5[395],
                      OutputImg5[394],OutputImg5[393],OutputImg5[392],
                      OutputImg5[391],OutputImg5[390],OutputImg5[389],
                      OutputImg5[388],OutputImg5[387],OutputImg5[386],
                      OutputImg5[385],OutputImg5[384]}), .EN (nx23706), .F ({
                      ImgReg5IN_383,ImgReg5IN_382,ImgReg5IN_381,ImgReg5IN_380,
                      ImgReg5IN_379,ImgReg5IN_378,ImgReg5IN_377,ImgReg5IN_376,
                      ImgReg5IN_375,ImgReg5IN_374,ImgReg5IN_373,ImgReg5IN_372,
                      ImgReg5IN_371,ImgReg5IN_370,ImgReg5IN_369,ImgReg5IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState0N (.D ({DATA[383],DATA[382],DATA[381],
                      DATA[380],DATA[379],DATA[378],DATA[377],DATA[376],
                      DATA[375],DATA[374],DATA[373],DATA[372],DATA[371],
                      DATA[370],DATA[369],DATA[368]}), .EN (nx23660), .F ({
                      ImgReg0IN_383,ImgReg0IN_382,ImgReg0IN_381,ImgReg0IN_380,
                      ImgReg0IN_379,ImgReg0IN_378,ImgReg0IN_377,ImgReg0IN_376,
                      ImgReg0IN_375,ImgReg0IN_374,ImgReg0IN_373,ImgReg0IN_372,
                      ImgReg0IN_371,ImgReg0IN_370,ImgReg0IN_369,ImgReg0IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState1N (.D ({DATA[383],DATA[382],DATA[381],
                      DATA[380],DATA[379],DATA[378],DATA[377],DATA[376],
                      DATA[375],DATA[374],DATA[373],DATA[372],DATA[371],
                      DATA[370],DATA[369],DATA[368]}), .EN (nx23648), .F ({
                      ImgReg1IN_383,ImgReg1IN_382,ImgReg1IN_381,ImgReg1IN_380,
                      ImgReg1IN_379,ImgReg1IN_378,ImgReg1IN_377,ImgReg1IN_376,
                      ImgReg1IN_375,ImgReg1IN_374,ImgReg1IN_373,ImgReg1IN_372,
                      ImgReg1IN_371,ImgReg1IN_370,ImgReg1IN_369,ImgReg1IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState2N (.D ({DATA[383],DATA[382],DATA[381],
                      DATA[380],DATA[379],DATA[378],DATA[377],DATA[376],
                      DATA[375],DATA[374],DATA[373],DATA[372],DATA[371],
                      DATA[370],DATA[369],DATA[368]}), .EN (nx23636), .F ({
                      ImgReg2IN_383,ImgReg2IN_382,ImgReg2IN_381,ImgReg2IN_380,
                      ImgReg2IN_379,ImgReg2IN_378,ImgReg2IN_377,ImgReg2IN_376,
                      ImgReg2IN_375,ImgReg2IN_374,ImgReg2IN_373,ImgReg2IN_372,
                      ImgReg2IN_371,ImgReg2IN_370,ImgReg2IN_369,ImgReg2IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState3N (.D ({DATA[383],DATA[382],DATA[381],
                      DATA[380],DATA[379],DATA[378],DATA[377],DATA[376],
                      DATA[375],DATA[374],DATA[373],DATA[372],DATA[371],
                      DATA[370],DATA[369],DATA[368]}), .EN (nx23624), .F ({
                      ImgReg3IN_383,ImgReg3IN_382,ImgReg3IN_381,ImgReg3IN_380,
                      ImgReg3IN_379,ImgReg3IN_378,ImgReg3IN_377,ImgReg3IN_376,
                      ImgReg3IN_375,ImgReg3IN_374,ImgReg3IN_373,ImgReg3IN_372,
                      ImgReg3IN_371,ImgReg3IN_370,ImgReg3IN_369,ImgReg3IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState4N (.D ({DATA[383],DATA[382],DATA[381],
                      DATA[380],DATA[379],DATA[378],DATA[377],DATA[376],
                      DATA[375],DATA[374],DATA[373],DATA[372],DATA[371],
                      DATA[370],DATA[369],DATA[368]}), .EN (nx23612), .F ({
                      ImgReg4IN_383,ImgReg4IN_382,ImgReg4IN_381,ImgReg4IN_380,
                      ImgReg4IN_379,ImgReg4IN_378,ImgReg4IN_377,ImgReg4IN_376,
                      ImgReg4IN_375,ImgReg4IN_374,ImgReg4IN_373,ImgReg4IN_372,
                      ImgReg4IN_371,ImgReg4IN_370,ImgReg4IN_369,ImgReg4IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState5N (.D ({DATA[383],DATA[382],DATA[381],
                      DATA[380],DATA[379],DATA[378],DATA[377],DATA[376],
                      DATA[375],DATA[374],DATA[373],DATA[372],DATA[371],
                      DATA[370],DATA[369],DATA[368]}), .EN (nx23600), .F ({
                      ImgReg5IN_383,ImgReg5IN_382,ImgReg5IN_381,ImgReg5IN_380,
                      ImgReg5IN_379,ImgReg5IN_378,ImgReg5IN_377,ImgReg5IN_376,
                      ImgReg5IN_375,ImgReg5IN_374,ImgReg5IN_373,ImgReg5IN_372,
                      ImgReg5IN_371,ImgReg5IN_370,ImgReg5IN_369,ImgReg5IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState0U (.D ({OutputImg1[383],OutputImg1[382],
                      OutputImg1[381],OutputImg1[380],OutputImg1[379],
                      OutputImg1[378],OutputImg1[377],OutputImg1[376],
                      OutputImg1[375],OutputImg1[374],OutputImg1[373],
                      OutputImg1[372],OutputImg1[371],OutputImg1[370],
                      OutputImg1[369],OutputImg1[368]}), .EN (nx23818), .F ({
                      ImgReg0IN_383,ImgReg0IN_382,ImgReg0IN_381,ImgReg0IN_380,
                      ImgReg0IN_379,ImgReg0IN_378,ImgReg0IN_377,ImgReg0IN_376,
                      ImgReg0IN_375,ImgReg0IN_374,ImgReg0IN_373,ImgReg0IN_372,
                      ImgReg0IN_371,ImgReg0IN_370,ImgReg0IN_369,ImgReg0IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState1U (.D ({OutputImg2[383],OutputImg2[382],
                      OutputImg2[381],OutputImg2[380],OutputImg2[379],
                      OutputImg2[378],OutputImg2[377],OutputImg2[376],
                      OutputImg2[375],OutputImg2[374],OutputImg2[373],
                      OutputImg2[372],OutputImg2[371],OutputImg2[370],
                      OutputImg2[369],OutputImg2[368]}), .EN (nx23818), .F ({
                      ImgReg1IN_383,ImgReg1IN_382,ImgReg1IN_381,ImgReg1IN_380,
                      ImgReg1IN_379,ImgReg1IN_378,ImgReg1IN_377,ImgReg1IN_376,
                      ImgReg1IN_375,ImgReg1IN_374,ImgReg1IN_373,ImgReg1IN_372,
                      ImgReg1IN_371,ImgReg1IN_370,ImgReg1IN_369,ImgReg1IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState2U (.D ({OutputImg3[383],OutputImg3[382],
                      OutputImg3[381],OutputImg3[380],OutputImg3[379],
                      OutputImg3[378],OutputImg3[377],OutputImg3[376],
                      OutputImg3[375],OutputImg3[374],OutputImg3[373],
                      OutputImg3[372],OutputImg3[371],OutputImg3[370],
                      OutputImg3[369],OutputImg3[368]}), .EN (nx23818), .F ({
                      ImgReg2IN_383,ImgReg2IN_382,ImgReg2IN_381,ImgReg2IN_380,
                      ImgReg2IN_379,ImgReg2IN_378,ImgReg2IN_377,ImgReg2IN_376,
                      ImgReg2IN_375,ImgReg2IN_374,ImgReg2IN_373,ImgReg2IN_372,
                      ImgReg2IN_371,ImgReg2IN_370,ImgReg2IN_369,ImgReg2IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState3U (.D ({OutputImg4[383],OutputImg4[382],
                      OutputImg4[381],OutputImg4[380],OutputImg4[379],
                      OutputImg4[378],OutputImg4[377],OutputImg4[376],
                      OutputImg4[375],OutputImg4[374],OutputImg4[373],
                      OutputImg4[372],OutputImg4[371],OutputImg4[370],
                      OutputImg4[369],OutputImg4[368]}), .EN (nx23818), .F ({
                      ImgReg3IN_383,ImgReg3IN_382,ImgReg3IN_381,ImgReg3IN_380,
                      ImgReg3IN_379,ImgReg3IN_378,ImgReg3IN_377,ImgReg3IN_376,
                      ImgReg3IN_375,ImgReg3IN_374,ImgReg3IN_373,ImgReg3IN_372,
                      ImgReg3IN_371,ImgReg3IN_370,ImgReg3IN_369,ImgReg3IN_368})
                      ) ;
    triStateBuffer_16 loop3_23_TriState4U (.D ({OutputImg5[383],OutputImg5[382],
                      OutputImg5[381],OutputImg5[380],OutputImg5[379],
                      OutputImg5[378],OutputImg5[377],OutputImg5[376],
                      OutputImg5[375],OutputImg5[374],OutputImg5[373],
                      OutputImg5[372],OutputImg5[371],OutputImg5[370],
                      OutputImg5[369],OutputImg5[368]}), .EN (nx23820), .F ({
                      ImgReg4IN_383,ImgReg4IN_382,ImgReg4IN_381,ImgReg4IN_380,
                      ImgReg4IN_379,ImgReg4IN_378,ImgReg4IN_377,ImgReg4IN_376,
                      ImgReg4IN_375,ImgReg4IN_374,ImgReg4IN_373,ImgReg4IN_372,
                      ImgReg4IN_371,ImgReg4IN_370,ImgReg4IN_369,ImgReg4IN_368})
                      ) ;
    nBitRegister_16 loop3_23_reg1 (.D ({ImgReg0IN_383,ImgReg0IN_382,
                    ImgReg0IN_381,ImgReg0IN_380,ImgReg0IN_379,ImgReg0IN_378,
                    ImgReg0IN_377,ImgReg0IN_376,ImgReg0IN_375,ImgReg0IN_374,
                    ImgReg0IN_373,ImgReg0IN_372,ImgReg0IN_371,ImgReg0IN_370,
                    ImgReg0IN_369,ImgReg0IN_368}), .CLK (nx23966), .RST (RST), .EN (
                    nx23724), .Q ({OutputImg0[383],OutputImg0[382],
                    OutputImg0[381],OutputImg0[380],OutputImg0[379],
                    OutputImg0[378],OutputImg0[377],OutputImg0[376],
                    OutputImg0[375],OutputImg0[374],OutputImg0[373],
                    OutputImg0[372],OutputImg0[371],OutputImg0[370],
                    OutputImg0[369],OutputImg0[368]})) ;
    nBitRegister_16 loop3_23_reg2 (.D ({ImgReg1IN_383,ImgReg1IN_382,
                    ImgReg1IN_381,ImgReg1IN_380,ImgReg1IN_379,ImgReg1IN_378,
                    ImgReg1IN_377,ImgReg1IN_376,ImgReg1IN_375,ImgReg1IN_374,
                    ImgReg1IN_373,ImgReg1IN_372,ImgReg1IN_371,ImgReg1IN_370,
                    ImgReg1IN_369,ImgReg1IN_368}), .CLK (nx23968), .RST (RST), .EN (
                    nx23734), .Q ({OutputImg1[383],OutputImg1[382],
                    OutputImg1[381],OutputImg1[380],OutputImg1[379],
                    OutputImg1[378],OutputImg1[377],OutputImg1[376],
                    OutputImg1[375],OutputImg1[374],OutputImg1[373],
                    OutputImg1[372],OutputImg1[371],OutputImg1[370],
                    OutputImg1[369],OutputImg1[368]})) ;
    nBitRegister_16 loop3_23_reg3 (.D ({ImgReg2IN_383,ImgReg2IN_382,
                    ImgReg2IN_381,ImgReg2IN_380,ImgReg2IN_379,ImgReg2IN_378,
                    ImgReg2IN_377,ImgReg2IN_376,ImgReg2IN_375,ImgReg2IN_374,
                    ImgReg2IN_373,ImgReg2IN_372,ImgReg2IN_371,ImgReg2IN_370,
                    ImgReg2IN_369,ImgReg2IN_368}), .CLK (nx23968), .RST (RST), .EN (
                    nx23744), .Q ({OutputImg2[383],OutputImg2[382],
                    OutputImg2[381],OutputImg2[380],OutputImg2[379],
                    OutputImg2[378],OutputImg2[377],OutputImg2[376],
                    OutputImg2[375],OutputImg2[374],OutputImg2[373],
                    OutputImg2[372],OutputImg2[371],OutputImg2[370],
                    OutputImg2[369],OutputImg2[368]})) ;
    nBitRegister_16 loop3_23_reg4 (.D ({ImgReg3IN_383,ImgReg3IN_382,
                    ImgReg3IN_381,ImgReg3IN_380,ImgReg3IN_379,ImgReg3IN_378,
                    ImgReg3IN_377,ImgReg3IN_376,ImgReg3IN_375,ImgReg3IN_374,
                    ImgReg3IN_373,ImgReg3IN_372,ImgReg3IN_371,ImgReg3IN_370,
                    ImgReg3IN_369,ImgReg3IN_368}), .CLK (nx23970), .RST (RST), .EN (
                    nx23754), .Q ({OutputImg3[383],OutputImg3[382],
                    OutputImg3[381],OutputImg3[380],OutputImg3[379],
                    OutputImg3[378],OutputImg3[377],OutputImg3[376],
                    OutputImg3[375],OutputImg3[374],OutputImg3[373],
                    OutputImg3[372],OutputImg3[371],OutputImg3[370],
                    OutputImg3[369],OutputImg3[368]})) ;
    nBitRegister_16 loop3_23_reg5 (.D ({ImgReg4IN_383,ImgReg4IN_382,
                    ImgReg4IN_381,ImgReg4IN_380,ImgReg4IN_379,ImgReg4IN_378,
                    ImgReg4IN_377,ImgReg4IN_376,ImgReg4IN_375,ImgReg4IN_374,
                    ImgReg4IN_373,ImgReg4IN_372,ImgReg4IN_371,ImgReg4IN_370,
                    ImgReg4IN_369,ImgReg4IN_368}), .CLK (nx23970), .RST (RST), .EN (
                    nx23764), .Q ({OutputImg4[383],OutputImg4[382],
                    OutputImg4[381],OutputImg4[380],OutputImg4[379],
                    OutputImg4[378],OutputImg4[377],OutputImg4[376],
                    OutputImg4[375],OutputImg4[374],OutputImg4[373],
                    OutputImg4[372],OutputImg4[371],OutputImg4[370],
                    OutputImg4[369],OutputImg4[368]})) ;
    nBitRegister_16 loop3_23_reg6 (.D ({ImgReg5IN_383,ImgReg5IN_382,
                    ImgReg5IN_381,ImgReg5IN_380,ImgReg5IN_379,ImgReg5IN_378,
                    ImgReg5IN_377,ImgReg5IN_376,ImgReg5IN_375,ImgReg5IN_374,
                    ImgReg5IN_373,ImgReg5IN_372,ImgReg5IN_371,ImgReg5IN_370,
                    ImgReg5IN_369,ImgReg5IN_368}), .CLK (nx23972), .RST (RST), .EN (
                    nx23774), .Q ({OutputImg5[383],OutputImg5[382],
                    OutputImg5[381],OutputImg5[380],OutputImg5[379],
                    OutputImg5[378],OutputImg5[377],OutputImg5[376],
                    OutputImg5[375],OutputImg5[374],OutputImg5[373],
                    OutputImg5[372],OutputImg5[371],OutputImg5[370],
                    OutputImg5[369],OutputImg5[368]})) ;
    triStateBuffer_16 loop3_24_TriState0L (.D ({OutputImg0[415],OutputImg0[414],
                      OutputImg0[413],OutputImg0[412],OutputImg0[411],
                      OutputImg0[410],OutputImg0[409],OutputImg0[408],
                      OutputImg0[407],OutputImg0[406],OutputImg0[405],
                      OutputImg0[404],OutputImg0[403],OutputImg0[402],
                      OutputImg0[401],OutputImg0[400]}), .EN (nx23706), .F ({
                      ImgReg0IN_399,ImgReg0IN_398,ImgReg0IN_397,ImgReg0IN_396,
                      ImgReg0IN_395,ImgReg0IN_394,ImgReg0IN_393,ImgReg0IN_392,
                      ImgReg0IN_391,ImgReg0IN_390,ImgReg0IN_389,ImgReg0IN_388,
                      ImgReg0IN_387,ImgReg0IN_386,ImgReg0IN_385,ImgReg0IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState1L (.D ({OutputImg1[415],OutputImg1[414],
                      OutputImg1[413],OutputImg1[412],OutputImg1[411],
                      OutputImg1[410],OutputImg1[409],OutputImg1[408],
                      OutputImg1[407],OutputImg1[406],OutputImg1[405],
                      OutputImg1[404],OutputImg1[403],OutputImg1[402],
                      OutputImg1[401],OutputImg1[400]}), .EN (nx23706), .F ({
                      ImgReg1IN_399,ImgReg1IN_398,ImgReg1IN_397,ImgReg1IN_396,
                      ImgReg1IN_395,ImgReg1IN_394,ImgReg1IN_393,ImgReg1IN_392,
                      ImgReg1IN_391,ImgReg1IN_390,ImgReg1IN_389,ImgReg1IN_388,
                      ImgReg1IN_387,ImgReg1IN_386,ImgReg1IN_385,ImgReg1IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState2L (.D ({OutputImg2[415],OutputImg2[414],
                      OutputImg2[413],OutputImg2[412],OutputImg2[411],
                      OutputImg2[410],OutputImg2[409],OutputImg2[408],
                      OutputImg2[407],OutputImg2[406],OutputImg2[405],
                      OutputImg2[404],OutputImg2[403],OutputImg2[402],
                      OutputImg2[401],OutputImg2[400]}), .EN (nx23706), .F ({
                      ImgReg2IN_399,ImgReg2IN_398,ImgReg2IN_397,ImgReg2IN_396,
                      ImgReg2IN_395,ImgReg2IN_394,ImgReg2IN_393,ImgReg2IN_392,
                      ImgReg2IN_391,ImgReg2IN_390,ImgReg2IN_389,ImgReg2IN_388,
                      ImgReg2IN_387,ImgReg2IN_386,ImgReg2IN_385,ImgReg2IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState3L (.D ({OutputImg3[415],OutputImg3[414],
                      OutputImg3[413],OutputImg3[412],OutputImg3[411],
                      OutputImg3[410],OutputImg3[409],OutputImg3[408],
                      OutputImg3[407],OutputImg3[406],OutputImg3[405],
                      OutputImg3[404],OutputImg3[403],OutputImg3[402],
                      OutputImg3[401],OutputImg3[400]}), .EN (nx23708), .F ({
                      ImgReg3IN_399,ImgReg3IN_398,ImgReg3IN_397,ImgReg3IN_396,
                      ImgReg3IN_395,ImgReg3IN_394,ImgReg3IN_393,ImgReg3IN_392,
                      ImgReg3IN_391,ImgReg3IN_390,ImgReg3IN_389,ImgReg3IN_388,
                      ImgReg3IN_387,ImgReg3IN_386,ImgReg3IN_385,ImgReg3IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState4L (.D ({OutputImg4[415],OutputImg4[414],
                      OutputImg4[413],OutputImg4[412],OutputImg4[411],
                      OutputImg4[410],OutputImg4[409],OutputImg4[408],
                      OutputImg4[407],OutputImg4[406],OutputImg4[405],
                      OutputImg4[404],OutputImg4[403],OutputImg4[402],
                      OutputImg4[401],OutputImg4[400]}), .EN (nx23708), .F ({
                      ImgReg4IN_399,ImgReg4IN_398,ImgReg4IN_397,ImgReg4IN_396,
                      ImgReg4IN_395,ImgReg4IN_394,ImgReg4IN_393,ImgReg4IN_392,
                      ImgReg4IN_391,ImgReg4IN_390,ImgReg4IN_389,ImgReg4IN_388,
                      ImgReg4IN_387,ImgReg4IN_386,ImgReg4IN_385,ImgReg4IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState5L (.D ({OutputImg5[415],OutputImg5[414],
                      OutputImg5[413],OutputImg5[412],OutputImg5[411],
                      OutputImg5[410],OutputImg5[409],OutputImg5[408],
                      OutputImg5[407],OutputImg5[406],OutputImg5[405],
                      OutputImg5[404],OutputImg5[403],OutputImg5[402],
                      OutputImg5[401],OutputImg5[400]}), .EN (nx23708), .F ({
                      ImgReg5IN_399,ImgReg5IN_398,ImgReg5IN_397,ImgReg5IN_396,
                      ImgReg5IN_395,ImgReg5IN_394,ImgReg5IN_393,ImgReg5IN_392,
                      ImgReg5IN_391,ImgReg5IN_390,ImgReg5IN_389,ImgReg5IN_388,
                      ImgReg5IN_387,ImgReg5IN_386,ImgReg5IN_385,ImgReg5IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState0N (.D ({DATA[399],DATA[398],DATA[397],
                      DATA[396],DATA[395],DATA[394],DATA[393],DATA[392],
                      DATA[391],DATA[390],DATA[389],DATA[388],DATA[387],
                      DATA[386],DATA[385],DATA[384]}), .EN (nx23660), .F ({
                      ImgReg0IN_399,ImgReg0IN_398,ImgReg0IN_397,ImgReg0IN_396,
                      ImgReg0IN_395,ImgReg0IN_394,ImgReg0IN_393,ImgReg0IN_392,
                      ImgReg0IN_391,ImgReg0IN_390,ImgReg0IN_389,ImgReg0IN_388,
                      ImgReg0IN_387,ImgReg0IN_386,ImgReg0IN_385,ImgReg0IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState1N (.D ({DATA[399],DATA[398],DATA[397],
                      DATA[396],DATA[395],DATA[394],DATA[393],DATA[392],
                      DATA[391],DATA[390],DATA[389],DATA[388],DATA[387],
                      DATA[386],DATA[385],DATA[384]}), .EN (nx23648), .F ({
                      ImgReg1IN_399,ImgReg1IN_398,ImgReg1IN_397,ImgReg1IN_396,
                      ImgReg1IN_395,ImgReg1IN_394,ImgReg1IN_393,ImgReg1IN_392,
                      ImgReg1IN_391,ImgReg1IN_390,ImgReg1IN_389,ImgReg1IN_388,
                      ImgReg1IN_387,ImgReg1IN_386,ImgReg1IN_385,ImgReg1IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState2N (.D ({DATA[399],DATA[398],DATA[397],
                      DATA[396],DATA[395],DATA[394],DATA[393],DATA[392],
                      DATA[391],DATA[390],DATA[389],DATA[388],DATA[387],
                      DATA[386],DATA[385],DATA[384]}), .EN (nx23636), .F ({
                      ImgReg2IN_399,ImgReg2IN_398,ImgReg2IN_397,ImgReg2IN_396,
                      ImgReg2IN_395,ImgReg2IN_394,ImgReg2IN_393,ImgReg2IN_392,
                      ImgReg2IN_391,ImgReg2IN_390,ImgReg2IN_389,ImgReg2IN_388,
                      ImgReg2IN_387,ImgReg2IN_386,ImgReg2IN_385,ImgReg2IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState3N (.D ({DATA[399],DATA[398],DATA[397],
                      DATA[396],DATA[395],DATA[394],DATA[393],DATA[392],
                      DATA[391],DATA[390],DATA[389],DATA[388],DATA[387],
                      DATA[386],DATA[385],DATA[384]}), .EN (nx23624), .F ({
                      ImgReg3IN_399,ImgReg3IN_398,ImgReg3IN_397,ImgReg3IN_396,
                      ImgReg3IN_395,ImgReg3IN_394,ImgReg3IN_393,ImgReg3IN_392,
                      ImgReg3IN_391,ImgReg3IN_390,ImgReg3IN_389,ImgReg3IN_388,
                      ImgReg3IN_387,ImgReg3IN_386,ImgReg3IN_385,ImgReg3IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState4N (.D ({DATA[399],DATA[398],DATA[397],
                      DATA[396],DATA[395],DATA[394],DATA[393],DATA[392],
                      DATA[391],DATA[390],DATA[389],DATA[388],DATA[387],
                      DATA[386],DATA[385],DATA[384]}), .EN (nx23612), .F ({
                      ImgReg4IN_399,ImgReg4IN_398,ImgReg4IN_397,ImgReg4IN_396,
                      ImgReg4IN_395,ImgReg4IN_394,ImgReg4IN_393,ImgReg4IN_392,
                      ImgReg4IN_391,ImgReg4IN_390,ImgReg4IN_389,ImgReg4IN_388,
                      ImgReg4IN_387,ImgReg4IN_386,ImgReg4IN_385,ImgReg4IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState5N (.D ({DATA[399],DATA[398],DATA[397],
                      DATA[396],DATA[395],DATA[394],DATA[393],DATA[392],
                      DATA[391],DATA[390],DATA[389],DATA[388],DATA[387],
                      DATA[386],DATA[385],DATA[384]}), .EN (nx23600), .F ({
                      ImgReg5IN_399,ImgReg5IN_398,ImgReg5IN_397,ImgReg5IN_396,
                      ImgReg5IN_395,ImgReg5IN_394,ImgReg5IN_393,ImgReg5IN_392,
                      ImgReg5IN_391,ImgReg5IN_390,ImgReg5IN_389,ImgReg5IN_388,
                      ImgReg5IN_387,ImgReg5IN_386,ImgReg5IN_385,ImgReg5IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState0U (.D ({OutputImg1[399],OutputImg1[398],
                      OutputImg1[397],OutputImg1[396],OutputImg1[395],
                      OutputImg1[394],OutputImg1[393],OutputImg1[392],
                      OutputImg1[391],OutputImg1[390],OutputImg1[389],
                      OutputImg1[388],OutputImg1[387],OutputImg1[386],
                      OutputImg1[385],OutputImg1[384]}), .EN (nx23820), .F ({
                      ImgReg0IN_399,ImgReg0IN_398,ImgReg0IN_397,ImgReg0IN_396,
                      ImgReg0IN_395,ImgReg0IN_394,ImgReg0IN_393,ImgReg0IN_392,
                      ImgReg0IN_391,ImgReg0IN_390,ImgReg0IN_389,ImgReg0IN_388,
                      ImgReg0IN_387,ImgReg0IN_386,ImgReg0IN_385,ImgReg0IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState1U (.D ({OutputImg2[399],OutputImg2[398],
                      OutputImg2[397],OutputImg2[396],OutputImg2[395],
                      OutputImg2[394],OutputImg2[393],OutputImg2[392],
                      OutputImg2[391],OutputImg2[390],OutputImg2[389],
                      OutputImg2[388],OutputImg2[387],OutputImg2[386],
                      OutputImg2[385],OutputImg2[384]}), .EN (nx23820), .F ({
                      ImgReg1IN_399,ImgReg1IN_398,ImgReg1IN_397,ImgReg1IN_396,
                      ImgReg1IN_395,ImgReg1IN_394,ImgReg1IN_393,ImgReg1IN_392,
                      ImgReg1IN_391,ImgReg1IN_390,ImgReg1IN_389,ImgReg1IN_388,
                      ImgReg1IN_387,ImgReg1IN_386,ImgReg1IN_385,ImgReg1IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState2U (.D ({OutputImg3[399],OutputImg3[398],
                      OutputImg3[397],OutputImg3[396],OutputImg3[395],
                      OutputImg3[394],OutputImg3[393],OutputImg3[392],
                      OutputImg3[391],OutputImg3[390],OutputImg3[389],
                      OutputImg3[388],OutputImg3[387],OutputImg3[386],
                      OutputImg3[385],OutputImg3[384]}), .EN (nx23820), .F ({
                      ImgReg2IN_399,ImgReg2IN_398,ImgReg2IN_397,ImgReg2IN_396,
                      ImgReg2IN_395,ImgReg2IN_394,ImgReg2IN_393,ImgReg2IN_392,
                      ImgReg2IN_391,ImgReg2IN_390,ImgReg2IN_389,ImgReg2IN_388,
                      ImgReg2IN_387,ImgReg2IN_386,ImgReg2IN_385,ImgReg2IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState3U (.D ({OutputImg4[399],OutputImg4[398],
                      OutputImg4[397],OutputImg4[396],OutputImg4[395],
                      OutputImg4[394],OutputImg4[393],OutputImg4[392],
                      OutputImg4[391],OutputImg4[390],OutputImg4[389],
                      OutputImg4[388],OutputImg4[387],OutputImg4[386],
                      OutputImg4[385],OutputImg4[384]}), .EN (nx23820), .F ({
                      ImgReg3IN_399,ImgReg3IN_398,ImgReg3IN_397,ImgReg3IN_396,
                      ImgReg3IN_395,ImgReg3IN_394,ImgReg3IN_393,ImgReg3IN_392,
                      ImgReg3IN_391,ImgReg3IN_390,ImgReg3IN_389,ImgReg3IN_388,
                      ImgReg3IN_387,ImgReg3IN_386,ImgReg3IN_385,ImgReg3IN_384})
                      ) ;
    triStateBuffer_16 loop3_24_TriState4U (.D ({OutputImg5[399],OutputImg5[398],
                      OutputImg5[397],OutputImg5[396],OutputImg5[395],
                      OutputImg5[394],OutputImg5[393],OutputImg5[392],
                      OutputImg5[391],OutputImg5[390],OutputImg5[389],
                      OutputImg5[388],OutputImg5[387],OutputImg5[386],
                      OutputImg5[385],OutputImg5[384]}), .EN (nx23820), .F ({
                      ImgReg4IN_399,ImgReg4IN_398,ImgReg4IN_397,ImgReg4IN_396,
                      ImgReg4IN_395,ImgReg4IN_394,ImgReg4IN_393,ImgReg4IN_392,
                      ImgReg4IN_391,ImgReg4IN_390,ImgReg4IN_389,ImgReg4IN_388,
                      ImgReg4IN_387,ImgReg4IN_386,ImgReg4IN_385,ImgReg4IN_384})
                      ) ;
    nBitRegister_16 loop3_24_reg1 (.D ({ImgReg0IN_399,ImgReg0IN_398,
                    ImgReg0IN_397,ImgReg0IN_396,ImgReg0IN_395,ImgReg0IN_394,
                    ImgReg0IN_393,ImgReg0IN_392,ImgReg0IN_391,ImgReg0IN_390,
                    ImgReg0IN_389,ImgReg0IN_388,ImgReg0IN_387,ImgReg0IN_386,
                    ImgReg0IN_385,ImgReg0IN_384}), .CLK (nx23972), .RST (RST), .EN (
                    nx23724), .Q ({OutputImg0[399],OutputImg0[398],
                    OutputImg0[397],OutputImg0[396],OutputImg0[395],
                    OutputImg0[394],OutputImg0[393],OutputImg0[392],
                    OutputImg0[391],OutputImg0[390],OutputImg0[389],
                    OutputImg0[388],OutputImg0[387],OutputImg0[386],
                    OutputImg0[385],OutputImg0[384]})) ;
    nBitRegister_16 loop3_24_reg2 (.D ({ImgReg1IN_399,ImgReg1IN_398,
                    ImgReg1IN_397,ImgReg1IN_396,ImgReg1IN_395,ImgReg1IN_394,
                    ImgReg1IN_393,ImgReg1IN_392,ImgReg1IN_391,ImgReg1IN_390,
                    ImgReg1IN_389,ImgReg1IN_388,ImgReg1IN_387,ImgReg1IN_386,
                    ImgReg1IN_385,ImgReg1IN_384}), .CLK (nx23974), .RST (RST), .EN (
                    nx23734), .Q ({OutputImg1[399],OutputImg1[398],
                    OutputImg1[397],OutputImg1[396],OutputImg1[395],
                    OutputImg1[394],OutputImg1[393],OutputImg1[392],
                    OutputImg1[391],OutputImg1[390],OutputImg1[389],
                    OutputImg1[388],OutputImg1[387],OutputImg1[386],
                    OutputImg1[385],OutputImg1[384]})) ;
    nBitRegister_16 loop3_24_reg3 (.D ({ImgReg2IN_399,ImgReg2IN_398,
                    ImgReg2IN_397,ImgReg2IN_396,ImgReg2IN_395,ImgReg2IN_394,
                    ImgReg2IN_393,ImgReg2IN_392,ImgReg2IN_391,ImgReg2IN_390,
                    ImgReg2IN_389,ImgReg2IN_388,ImgReg2IN_387,ImgReg2IN_386,
                    ImgReg2IN_385,ImgReg2IN_384}), .CLK (nx23974), .RST (RST), .EN (
                    nx23744), .Q ({OutputImg2[399],OutputImg2[398],
                    OutputImg2[397],OutputImg2[396],OutputImg2[395],
                    OutputImg2[394],OutputImg2[393],OutputImg2[392],
                    OutputImg2[391],OutputImg2[390],OutputImg2[389],
                    OutputImg2[388],OutputImg2[387],OutputImg2[386],
                    OutputImg2[385],OutputImg2[384]})) ;
    nBitRegister_16 loop3_24_reg4 (.D ({ImgReg3IN_399,ImgReg3IN_398,
                    ImgReg3IN_397,ImgReg3IN_396,ImgReg3IN_395,ImgReg3IN_394,
                    ImgReg3IN_393,ImgReg3IN_392,ImgReg3IN_391,ImgReg3IN_390,
                    ImgReg3IN_389,ImgReg3IN_388,ImgReg3IN_387,ImgReg3IN_386,
                    ImgReg3IN_385,ImgReg3IN_384}), .CLK (nx23976), .RST (RST), .EN (
                    nx23754), .Q ({OutputImg3[399],OutputImg3[398],
                    OutputImg3[397],OutputImg3[396],OutputImg3[395],
                    OutputImg3[394],OutputImg3[393],OutputImg3[392],
                    OutputImg3[391],OutputImg3[390],OutputImg3[389],
                    OutputImg3[388],OutputImg3[387],OutputImg3[386],
                    OutputImg3[385],OutputImg3[384]})) ;
    nBitRegister_16 loop3_24_reg5 (.D ({ImgReg4IN_399,ImgReg4IN_398,
                    ImgReg4IN_397,ImgReg4IN_396,ImgReg4IN_395,ImgReg4IN_394,
                    ImgReg4IN_393,ImgReg4IN_392,ImgReg4IN_391,ImgReg4IN_390,
                    ImgReg4IN_389,ImgReg4IN_388,ImgReg4IN_387,ImgReg4IN_386,
                    ImgReg4IN_385,ImgReg4IN_384}), .CLK (nx23976), .RST (RST), .EN (
                    nx23764), .Q ({OutputImg4[399],OutputImg4[398],
                    OutputImg4[397],OutputImg4[396],OutputImg4[395],
                    OutputImg4[394],OutputImg4[393],OutputImg4[392],
                    OutputImg4[391],OutputImg4[390],OutputImg4[389],
                    OutputImg4[388],OutputImg4[387],OutputImg4[386],
                    OutputImg4[385],OutputImg4[384]})) ;
    nBitRegister_16 loop3_24_reg6 (.D ({ImgReg5IN_399,ImgReg5IN_398,
                    ImgReg5IN_397,ImgReg5IN_396,ImgReg5IN_395,ImgReg5IN_394,
                    ImgReg5IN_393,ImgReg5IN_392,ImgReg5IN_391,ImgReg5IN_390,
                    ImgReg5IN_389,ImgReg5IN_388,ImgReg5IN_387,ImgReg5IN_386,
                    ImgReg5IN_385,ImgReg5IN_384}), .CLK (nx23978), .RST (RST), .EN (
                    nx23774), .Q ({OutputImg5[399],OutputImg5[398],
                    OutputImg5[397],OutputImg5[396],OutputImg5[395],
                    OutputImg5[394],OutputImg5[393],OutputImg5[392],
                    OutputImg5[391],OutputImg5[390],OutputImg5[389],
                    OutputImg5[388],OutputImg5[387],OutputImg5[386],
                    OutputImg5[385],OutputImg5[384]})) ;
    triStateBuffer_16 loop3_25_TriState0L (.D ({OutputImg0[431],OutputImg0[430],
                      OutputImg0[429],OutputImg0[428],OutputImg0[427],
                      OutputImg0[426],OutputImg0[425],OutputImg0[424],
                      OutputImg0[423],OutputImg0[422],OutputImg0[421],
                      OutputImg0[420],OutputImg0[419],OutputImg0[418],
                      OutputImg0[417],OutputImg0[416]}), .EN (nx23708), .F ({
                      ImgReg0IN_415,ImgReg0IN_414,ImgReg0IN_413,ImgReg0IN_412,
                      ImgReg0IN_411,ImgReg0IN_410,ImgReg0IN_409,ImgReg0IN_408,
                      ImgReg0IN_407,ImgReg0IN_406,ImgReg0IN_405,ImgReg0IN_404,
                      ImgReg0IN_403,ImgReg0IN_402,ImgReg0IN_401,ImgReg0IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState1L (.D ({OutputImg1[431],OutputImg1[430],
                      OutputImg1[429],OutputImg1[428],OutputImg1[427],
                      OutputImg1[426],OutputImg1[425],OutputImg1[424],
                      OutputImg1[423],OutputImg1[422],OutputImg1[421],
                      OutputImg1[420],OutputImg1[419],OutputImg1[418],
                      OutputImg1[417],OutputImg1[416]}), .EN (nx23708), .F ({
                      ImgReg1IN_415,ImgReg1IN_414,ImgReg1IN_413,ImgReg1IN_412,
                      ImgReg1IN_411,ImgReg1IN_410,ImgReg1IN_409,ImgReg1IN_408,
                      ImgReg1IN_407,ImgReg1IN_406,ImgReg1IN_405,ImgReg1IN_404,
                      ImgReg1IN_403,ImgReg1IN_402,ImgReg1IN_401,ImgReg1IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState2L (.D ({OutputImg2[431],OutputImg2[430],
                      OutputImg2[429],OutputImg2[428],OutputImg2[427],
                      OutputImg2[426],OutputImg2[425],OutputImg2[424],
                      OutputImg2[423],OutputImg2[422],OutputImg2[421],
                      OutputImg2[420],OutputImg2[419],OutputImg2[418],
                      OutputImg2[417],OutputImg2[416]}), .EN (nx23708), .F ({
                      ImgReg2IN_415,ImgReg2IN_414,ImgReg2IN_413,ImgReg2IN_412,
                      ImgReg2IN_411,ImgReg2IN_410,ImgReg2IN_409,ImgReg2IN_408,
                      ImgReg2IN_407,ImgReg2IN_406,ImgReg2IN_405,ImgReg2IN_404,
                      ImgReg2IN_403,ImgReg2IN_402,ImgReg2IN_401,ImgReg2IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState3L (.D ({OutputImg3[431],OutputImg3[430],
                      OutputImg3[429],OutputImg3[428],OutputImg3[427],
                      OutputImg3[426],OutputImg3[425],OutputImg3[424],
                      OutputImg3[423],OutputImg3[422],OutputImg3[421],
                      OutputImg3[420],OutputImg3[419],OutputImg3[418],
                      OutputImg3[417],OutputImg3[416]}), .EN (nx23708), .F ({
                      ImgReg3IN_415,ImgReg3IN_414,ImgReg3IN_413,ImgReg3IN_412,
                      ImgReg3IN_411,ImgReg3IN_410,ImgReg3IN_409,ImgReg3IN_408,
                      ImgReg3IN_407,ImgReg3IN_406,ImgReg3IN_405,ImgReg3IN_404,
                      ImgReg3IN_403,ImgReg3IN_402,ImgReg3IN_401,ImgReg3IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState4L (.D ({OutputImg4[431],OutputImg4[430],
                      OutputImg4[429],OutputImg4[428],OutputImg4[427],
                      OutputImg4[426],OutputImg4[425],OutputImg4[424],
                      OutputImg4[423],OutputImg4[422],OutputImg4[421],
                      OutputImg4[420],OutputImg4[419],OutputImg4[418],
                      OutputImg4[417],OutputImg4[416]}), .EN (nx23710), .F ({
                      ImgReg4IN_415,ImgReg4IN_414,ImgReg4IN_413,ImgReg4IN_412,
                      ImgReg4IN_411,ImgReg4IN_410,ImgReg4IN_409,ImgReg4IN_408,
                      ImgReg4IN_407,ImgReg4IN_406,ImgReg4IN_405,ImgReg4IN_404,
                      ImgReg4IN_403,ImgReg4IN_402,ImgReg4IN_401,ImgReg4IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState5L (.D ({OutputImg5[431],OutputImg5[430],
                      OutputImg5[429],OutputImg5[428],OutputImg5[427],
                      OutputImg5[426],OutputImg5[425],OutputImg5[424],
                      OutputImg5[423],OutputImg5[422],OutputImg5[421],
                      OutputImg5[420],OutputImg5[419],OutputImg5[418],
                      OutputImg5[417],OutputImg5[416]}), .EN (nx23710), .F ({
                      ImgReg5IN_415,ImgReg5IN_414,ImgReg5IN_413,ImgReg5IN_412,
                      ImgReg5IN_411,ImgReg5IN_410,ImgReg5IN_409,ImgReg5IN_408,
                      ImgReg5IN_407,ImgReg5IN_406,ImgReg5IN_405,ImgReg5IN_404,
                      ImgReg5IN_403,ImgReg5IN_402,ImgReg5IN_401,ImgReg5IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState0N (.D ({DATA[415],DATA[414],DATA[413],
                      DATA[412],DATA[411],DATA[410],DATA[409],DATA[408],
                      DATA[407],DATA[406],DATA[405],DATA[404],DATA[403],
                      DATA[402],DATA[401],DATA[400]}), .EN (nx23660), .F ({
                      ImgReg0IN_415,ImgReg0IN_414,ImgReg0IN_413,ImgReg0IN_412,
                      ImgReg0IN_411,ImgReg0IN_410,ImgReg0IN_409,ImgReg0IN_408,
                      ImgReg0IN_407,ImgReg0IN_406,ImgReg0IN_405,ImgReg0IN_404,
                      ImgReg0IN_403,ImgReg0IN_402,ImgReg0IN_401,ImgReg0IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState1N (.D ({DATA[415],DATA[414],DATA[413],
                      DATA[412],DATA[411],DATA[410],DATA[409],DATA[408],
                      DATA[407],DATA[406],DATA[405],DATA[404],DATA[403],
                      DATA[402],DATA[401],DATA[400]}), .EN (nx23648), .F ({
                      ImgReg1IN_415,ImgReg1IN_414,ImgReg1IN_413,ImgReg1IN_412,
                      ImgReg1IN_411,ImgReg1IN_410,ImgReg1IN_409,ImgReg1IN_408,
                      ImgReg1IN_407,ImgReg1IN_406,ImgReg1IN_405,ImgReg1IN_404,
                      ImgReg1IN_403,ImgReg1IN_402,ImgReg1IN_401,ImgReg1IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState2N (.D ({DATA[415],DATA[414],DATA[413],
                      DATA[412],DATA[411],DATA[410],DATA[409],DATA[408],
                      DATA[407],DATA[406],DATA[405],DATA[404],DATA[403],
                      DATA[402],DATA[401],DATA[400]}), .EN (nx23636), .F ({
                      ImgReg2IN_415,ImgReg2IN_414,ImgReg2IN_413,ImgReg2IN_412,
                      ImgReg2IN_411,ImgReg2IN_410,ImgReg2IN_409,ImgReg2IN_408,
                      ImgReg2IN_407,ImgReg2IN_406,ImgReg2IN_405,ImgReg2IN_404,
                      ImgReg2IN_403,ImgReg2IN_402,ImgReg2IN_401,ImgReg2IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState3N (.D ({DATA[415],DATA[414],DATA[413],
                      DATA[412],DATA[411],DATA[410],DATA[409],DATA[408],
                      DATA[407],DATA[406],DATA[405],DATA[404],DATA[403],
                      DATA[402],DATA[401],DATA[400]}), .EN (nx23624), .F ({
                      ImgReg3IN_415,ImgReg3IN_414,ImgReg3IN_413,ImgReg3IN_412,
                      ImgReg3IN_411,ImgReg3IN_410,ImgReg3IN_409,ImgReg3IN_408,
                      ImgReg3IN_407,ImgReg3IN_406,ImgReg3IN_405,ImgReg3IN_404,
                      ImgReg3IN_403,ImgReg3IN_402,ImgReg3IN_401,ImgReg3IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState4N (.D ({DATA[415],DATA[414],DATA[413],
                      DATA[412],DATA[411],DATA[410],DATA[409],DATA[408],
                      DATA[407],DATA[406],DATA[405],DATA[404],DATA[403],
                      DATA[402],DATA[401],DATA[400]}), .EN (nx23612), .F ({
                      ImgReg4IN_415,ImgReg4IN_414,ImgReg4IN_413,ImgReg4IN_412,
                      ImgReg4IN_411,ImgReg4IN_410,ImgReg4IN_409,ImgReg4IN_408,
                      ImgReg4IN_407,ImgReg4IN_406,ImgReg4IN_405,ImgReg4IN_404,
                      ImgReg4IN_403,ImgReg4IN_402,ImgReg4IN_401,ImgReg4IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState5N (.D ({DATA[415],DATA[414],DATA[413],
                      DATA[412],DATA[411],DATA[410],DATA[409],DATA[408],
                      DATA[407],DATA[406],DATA[405],DATA[404],DATA[403],
                      DATA[402],DATA[401],DATA[400]}), .EN (nx23600), .F ({
                      ImgReg5IN_415,ImgReg5IN_414,ImgReg5IN_413,ImgReg5IN_412,
                      ImgReg5IN_411,ImgReg5IN_410,ImgReg5IN_409,ImgReg5IN_408,
                      ImgReg5IN_407,ImgReg5IN_406,ImgReg5IN_405,ImgReg5IN_404,
                      ImgReg5IN_403,ImgReg5IN_402,ImgReg5IN_401,ImgReg5IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState0U (.D ({OutputImg1[415],OutputImg1[414],
                      OutputImg1[413],OutputImg1[412],OutputImg1[411],
                      OutputImg1[410],OutputImg1[409],OutputImg1[408],
                      OutputImg1[407],OutputImg1[406],OutputImg1[405],
                      OutputImg1[404],OutputImg1[403],OutputImg1[402],
                      OutputImg1[401],OutputImg1[400]}), .EN (nx23820), .F ({
                      ImgReg0IN_415,ImgReg0IN_414,ImgReg0IN_413,ImgReg0IN_412,
                      ImgReg0IN_411,ImgReg0IN_410,ImgReg0IN_409,ImgReg0IN_408,
                      ImgReg0IN_407,ImgReg0IN_406,ImgReg0IN_405,ImgReg0IN_404,
                      ImgReg0IN_403,ImgReg0IN_402,ImgReg0IN_401,ImgReg0IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState1U (.D ({OutputImg2[415],OutputImg2[414],
                      OutputImg2[413],OutputImg2[412],OutputImg2[411],
                      OutputImg2[410],OutputImg2[409],OutputImg2[408],
                      OutputImg2[407],OutputImg2[406],OutputImg2[405],
                      OutputImg2[404],OutputImg2[403],OutputImg2[402],
                      OutputImg2[401],OutputImg2[400]}), .EN (nx23822), .F ({
                      ImgReg1IN_415,ImgReg1IN_414,ImgReg1IN_413,ImgReg1IN_412,
                      ImgReg1IN_411,ImgReg1IN_410,ImgReg1IN_409,ImgReg1IN_408,
                      ImgReg1IN_407,ImgReg1IN_406,ImgReg1IN_405,ImgReg1IN_404,
                      ImgReg1IN_403,ImgReg1IN_402,ImgReg1IN_401,ImgReg1IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState2U (.D ({OutputImg3[415],OutputImg3[414],
                      OutputImg3[413],OutputImg3[412],OutputImg3[411],
                      OutputImg3[410],OutputImg3[409],OutputImg3[408],
                      OutputImg3[407],OutputImg3[406],OutputImg3[405],
                      OutputImg3[404],OutputImg3[403],OutputImg3[402],
                      OutputImg3[401],OutputImg3[400]}), .EN (nx23822), .F ({
                      ImgReg2IN_415,ImgReg2IN_414,ImgReg2IN_413,ImgReg2IN_412,
                      ImgReg2IN_411,ImgReg2IN_410,ImgReg2IN_409,ImgReg2IN_408,
                      ImgReg2IN_407,ImgReg2IN_406,ImgReg2IN_405,ImgReg2IN_404,
                      ImgReg2IN_403,ImgReg2IN_402,ImgReg2IN_401,ImgReg2IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState3U (.D ({OutputImg4[415],OutputImg4[414],
                      OutputImg4[413],OutputImg4[412],OutputImg4[411],
                      OutputImg4[410],OutputImg4[409],OutputImg4[408],
                      OutputImg4[407],OutputImg4[406],OutputImg4[405],
                      OutputImg4[404],OutputImg4[403],OutputImg4[402],
                      OutputImg4[401],OutputImg4[400]}), .EN (nx23822), .F ({
                      ImgReg3IN_415,ImgReg3IN_414,ImgReg3IN_413,ImgReg3IN_412,
                      ImgReg3IN_411,ImgReg3IN_410,ImgReg3IN_409,ImgReg3IN_408,
                      ImgReg3IN_407,ImgReg3IN_406,ImgReg3IN_405,ImgReg3IN_404,
                      ImgReg3IN_403,ImgReg3IN_402,ImgReg3IN_401,ImgReg3IN_400})
                      ) ;
    triStateBuffer_16 loop3_25_TriState4U (.D ({OutputImg5[415],OutputImg5[414],
                      OutputImg5[413],OutputImg5[412],OutputImg5[411],
                      OutputImg5[410],OutputImg5[409],OutputImg5[408],
                      OutputImg5[407],OutputImg5[406],OutputImg5[405],
                      OutputImg5[404],OutputImg5[403],OutputImg5[402],
                      OutputImg5[401],OutputImg5[400]}), .EN (nx23822), .F ({
                      ImgReg4IN_415,ImgReg4IN_414,ImgReg4IN_413,ImgReg4IN_412,
                      ImgReg4IN_411,ImgReg4IN_410,ImgReg4IN_409,ImgReg4IN_408,
                      ImgReg4IN_407,ImgReg4IN_406,ImgReg4IN_405,ImgReg4IN_404,
                      ImgReg4IN_403,ImgReg4IN_402,ImgReg4IN_401,ImgReg4IN_400})
                      ) ;
    nBitRegister_16 loop3_25_reg1 (.D ({ImgReg0IN_415,ImgReg0IN_414,
                    ImgReg0IN_413,ImgReg0IN_412,ImgReg0IN_411,ImgReg0IN_410,
                    ImgReg0IN_409,ImgReg0IN_408,ImgReg0IN_407,ImgReg0IN_406,
                    ImgReg0IN_405,ImgReg0IN_404,ImgReg0IN_403,ImgReg0IN_402,
                    ImgReg0IN_401,ImgReg0IN_400}), .CLK (nx23978), .RST (RST), .EN (
                    nx23724), .Q ({OutputImg0[415],OutputImg0[414],
                    OutputImg0[413],OutputImg0[412],OutputImg0[411],
                    OutputImg0[410],OutputImg0[409],OutputImg0[408],
                    OutputImg0[407],OutputImg0[406],OutputImg0[405],
                    OutputImg0[404],OutputImg0[403],OutputImg0[402],
                    OutputImg0[401],OutputImg0[400]})) ;
    nBitRegister_16 loop3_25_reg2 (.D ({ImgReg1IN_415,ImgReg1IN_414,
                    ImgReg1IN_413,ImgReg1IN_412,ImgReg1IN_411,ImgReg1IN_410,
                    ImgReg1IN_409,ImgReg1IN_408,ImgReg1IN_407,ImgReg1IN_406,
                    ImgReg1IN_405,ImgReg1IN_404,ImgReg1IN_403,ImgReg1IN_402,
                    ImgReg1IN_401,ImgReg1IN_400}), .CLK (nx23980), .RST (RST), .EN (
                    nx23734), .Q ({OutputImg1[415],OutputImg1[414],
                    OutputImg1[413],OutputImg1[412],OutputImg1[411],
                    OutputImg1[410],OutputImg1[409],OutputImg1[408],
                    OutputImg1[407],OutputImg1[406],OutputImg1[405],
                    OutputImg1[404],OutputImg1[403],OutputImg1[402],
                    OutputImg1[401],OutputImg1[400]})) ;
    nBitRegister_16 loop3_25_reg3 (.D ({ImgReg2IN_415,ImgReg2IN_414,
                    ImgReg2IN_413,ImgReg2IN_412,ImgReg2IN_411,ImgReg2IN_410,
                    ImgReg2IN_409,ImgReg2IN_408,ImgReg2IN_407,ImgReg2IN_406,
                    ImgReg2IN_405,ImgReg2IN_404,ImgReg2IN_403,ImgReg2IN_402,
                    ImgReg2IN_401,ImgReg2IN_400}), .CLK (nx23980), .RST (RST), .EN (
                    nx23744), .Q ({OutputImg2[415],OutputImg2[414],
                    OutputImg2[413],OutputImg2[412],OutputImg2[411],
                    OutputImg2[410],OutputImg2[409],OutputImg2[408],
                    OutputImg2[407],OutputImg2[406],OutputImg2[405],
                    OutputImg2[404],OutputImg2[403],OutputImg2[402],
                    OutputImg2[401],OutputImg2[400]})) ;
    nBitRegister_16 loop3_25_reg4 (.D ({ImgReg3IN_415,ImgReg3IN_414,
                    ImgReg3IN_413,ImgReg3IN_412,ImgReg3IN_411,ImgReg3IN_410,
                    ImgReg3IN_409,ImgReg3IN_408,ImgReg3IN_407,ImgReg3IN_406,
                    ImgReg3IN_405,ImgReg3IN_404,ImgReg3IN_403,ImgReg3IN_402,
                    ImgReg3IN_401,ImgReg3IN_400}), .CLK (nx23982), .RST (RST), .EN (
                    nx23754), .Q ({OutputImg3[415],OutputImg3[414],
                    OutputImg3[413],OutputImg3[412],OutputImg3[411],
                    OutputImg3[410],OutputImg3[409],OutputImg3[408],
                    OutputImg3[407],OutputImg3[406],OutputImg3[405],
                    OutputImg3[404],OutputImg3[403],OutputImg3[402],
                    OutputImg3[401],OutputImg3[400]})) ;
    nBitRegister_16 loop3_25_reg5 (.D ({ImgReg4IN_415,ImgReg4IN_414,
                    ImgReg4IN_413,ImgReg4IN_412,ImgReg4IN_411,ImgReg4IN_410,
                    ImgReg4IN_409,ImgReg4IN_408,ImgReg4IN_407,ImgReg4IN_406,
                    ImgReg4IN_405,ImgReg4IN_404,ImgReg4IN_403,ImgReg4IN_402,
                    ImgReg4IN_401,ImgReg4IN_400}), .CLK (nx23982), .RST (RST), .EN (
                    nx23764), .Q ({OutputImg4[415],OutputImg4[414],
                    OutputImg4[413],OutputImg4[412],OutputImg4[411],
                    OutputImg4[410],OutputImg4[409],OutputImg4[408],
                    OutputImg4[407],OutputImg4[406],OutputImg4[405],
                    OutputImg4[404],OutputImg4[403],OutputImg4[402],
                    OutputImg4[401],OutputImg4[400]})) ;
    nBitRegister_16 loop3_25_reg6 (.D ({ImgReg5IN_415,ImgReg5IN_414,
                    ImgReg5IN_413,ImgReg5IN_412,ImgReg5IN_411,ImgReg5IN_410,
                    ImgReg5IN_409,ImgReg5IN_408,ImgReg5IN_407,ImgReg5IN_406,
                    ImgReg5IN_405,ImgReg5IN_404,ImgReg5IN_403,ImgReg5IN_402,
                    ImgReg5IN_401,ImgReg5IN_400}), .CLK (nx23984), .RST (RST), .EN (
                    nx23774), .Q ({OutputImg5[415],OutputImg5[414],
                    OutputImg5[413],OutputImg5[412],OutputImg5[411],
                    OutputImg5[410],OutputImg5[409],OutputImg5[408],
                    OutputImg5[407],OutputImg5[406],OutputImg5[405],
                    OutputImg5[404],OutputImg5[403],OutputImg5[402],
                    OutputImg5[401],OutputImg5[400]})) ;
    triStateBuffer_16 loop3_26_TriState0L (.D ({OutputImg0[447],OutputImg0[446],
                      OutputImg0[445],OutputImg0[444],OutputImg0[443],
                      OutputImg0[442],OutputImg0[441],OutputImg0[440],
                      OutputImg0[439],OutputImg0[438],OutputImg0[437],
                      OutputImg0[436],OutputImg0[435],OutputImg0[434],
                      OutputImg0[433],OutputImg0[432]}), .EN (nx23710), .F ({
                      ImgReg0IN_431,ImgReg0IN_430,ImgReg0IN_429,ImgReg0IN_428,
                      ImgReg0IN_427,ImgReg0IN_426,ImgReg0IN_425,ImgReg0IN_424,
                      ImgReg0IN_423,ImgReg0IN_422,ImgReg0IN_421,ImgReg0IN_420,
                      ImgReg0IN_419,ImgReg0IN_418,ImgReg0IN_417,ImgReg0IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState1L (.D ({OutputImg1[447],OutputImg1[446],
                      OutputImg1[445],OutputImg1[444],OutputImg1[443],
                      OutputImg1[442],OutputImg1[441],OutputImg1[440],
                      OutputImg1[439],OutputImg1[438],OutputImg1[437],
                      OutputImg1[436],OutputImg1[435],OutputImg1[434],
                      OutputImg1[433],OutputImg1[432]}), .EN (nx23710), .F ({
                      ImgReg1IN_431,ImgReg1IN_430,ImgReg1IN_429,ImgReg1IN_428,
                      ImgReg1IN_427,ImgReg1IN_426,ImgReg1IN_425,ImgReg1IN_424,
                      ImgReg1IN_423,ImgReg1IN_422,ImgReg1IN_421,ImgReg1IN_420,
                      ImgReg1IN_419,ImgReg1IN_418,ImgReg1IN_417,ImgReg1IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState2L (.D ({OutputImg2[447],OutputImg2[446],
                      OutputImg2[445],OutputImg2[444],OutputImg2[443],
                      OutputImg2[442],OutputImg2[441],OutputImg2[440],
                      OutputImg2[439],OutputImg2[438],OutputImg2[437],
                      OutputImg2[436],OutputImg2[435],OutputImg2[434],
                      OutputImg2[433],OutputImg2[432]}), .EN (nx23710), .F ({
                      ImgReg2IN_431,ImgReg2IN_430,ImgReg2IN_429,ImgReg2IN_428,
                      ImgReg2IN_427,ImgReg2IN_426,ImgReg2IN_425,ImgReg2IN_424,
                      ImgReg2IN_423,ImgReg2IN_422,ImgReg2IN_421,ImgReg2IN_420,
                      ImgReg2IN_419,ImgReg2IN_418,ImgReg2IN_417,ImgReg2IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState3L (.D ({OutputImg3[447],OutputImg3[446],
                      OutputImg3[445],OutputImg3[444],OutputImg3[443],
                      OutputImg3[442],OutputImg3[441],OutputImg3[440],
                      OutputImg3[439],OutputImg3[438],OutputImg3[437],
                      OutputImg3[436],OutputImg3[435],OutputImg3[434],
                      OutputImg3[433],OutputImg3[432]}), .EN (nx23710), .F ({
                      ImgReg3IN_431,ImgReg3IN_430,ImgReg3IN_429,ImgReg3IN_428,
                      ImgReg3IN_427,ImgReg3IN_426,ImgReg3IN_425,ImgReg3IN_424,
                      ImgReg3IN_423,ImgReg3IN_422,ImgReg3IN_421,ImgReg3IN_420,
                      ImgReg3IN_419,ImgReg3IN_418,ImgReg3IN_417,ImgReg3IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState4L (.D ({OutputImg4[447],OutputImg4[446],
                      OutputImg4[445],OutputImg4[444],OutputImg4[443],
                      OutputImg4[442],OutputImg4[441],OutputImg4[440],
                      OutputImg4[439],OutputImg4[438],OutputImg4[437],
                      OutputImg4[436],OutputImg4[435],OutputImg4[434],
                      OutputImg4[433],OutputImg4[432]}), .EN (nx23710), .F ({
                      ImgReg4IN_431,ImgReg4IN_430,ImgReg4IN_429,ImgReg4IN_428,
                      ImgReg4IN_427,ImgReg4IN_426,ImgReg4IN_425,ImgReg4IN_424,
                      ImgReg4IN_423,ImgReg4IN_422,ImgReg4IN_421,ImgReg4IN_420,
                      ImgReg4IN_419,ImgReg4IN_418,ImgReg4IN_417,ImgReg4IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState5L (.D ({OutputImg5[447],OutputImg5[446],
                      OutputImg5[445],OutputImg5[444],OutputImg5[443],
                      OutputImg5[442],OutputImg5[441],OutputImg5[440],
                      OutputImg5[439],OutputImg5[438],OutputImg5[437],
                      OutputImg5[436],OutputImg5[435],OutputImg5[434],
                      OutputImg5[433],OutputImg5[432]}), .EN (nx23712), .F ({
                      ImgReg5IN_431,ImgReg5IN_430,ImgReg5IN_429,ImgReg5IN_428,
                      ImgReg5IN_427,ImgReg5IN_426,ImgReg5IN_425,ImgReg5IN_424,
                      ImgReg5IN_423,ImgReg5IN_422,ImgReg5IN_421,ImgReg5IN_420,
                      ImgReg5IN_419,ImgReg5IN_418,ImgReg5IN_417,ImgReg5IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState0N (.D ({DATA[431],DATA[430],DATA[429],
                      DATA[428],DATA[427],DATA[426],DATA[425],DATA[424],
                      DATA[423],DATA[422],DATA[421],DATA[420],DATA[419],
                      DATA[418],DATA[417],DATA[416]}), .EN (nx23660), .F ({
                      ImgReg0IN_431,ImgReg0IN_430,ImgReg0IN_429,ImgReg0IN_428,
                      ImgReg0IN_427,ImgReg0IN_426,ImgReg0IN_425,ImgReg0IN_424,
                      ImgReg0IN_423,ImgReg0IN_422,ImgReg0IN_421,ImgReg0IN_420,
                      ImgReg0IN_419,ImgReg0IN_418,ImgReg0IN_417,ImgReg0IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState1N (.D ({DATA[431],DATA[430],DATA[429],
                      DATA[428],DATA[427],DATA[426],DATA[425],DATA[424],
                      DATA[423],DATA[422],DATA[421],DATA[420],DATA[419],
                      DATA[418],DATA[417],DATA[416]}), .EN (nx23648), .F ({
                      ImgReg1IN_431,ImgReg1IN_430,ImgReg1IN_429,ImgReg1IN_428,
                      ImgReg1IN_427,ImgReg1IN_426,ImgReg1IN_425,ImgReg1IN_424,
                      ImgReg1IN_423,ImgReg1IN_422,ImgReg1IN_421,ImgReg1IN_420,
                      ImgReg1IN_419,ImgReg1IN_418,ImgReg1IN_417,ImgReg1IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState2N (.D ({DATA[431],DATA[430],DATA[429],
                      DATA[428],DATA[427],DATA[426],DATA[425],DATA[424],
                      DATA[423],DATA[422],DATA[421],DATA[420],DATA[419],
                      DATA[418],DATA[417],DATA[416]}), .EN (nx23636), .F ({
                      ImgReg2IN_431,ImgReg2IN_430,ImgReg2IN_429,ImgReg2IN_428,
                      ImgReg2IN_427,ImgReg2IN_426,ImgReg2IN_425,ImgReg2IN_424,
                      ImgReg2IN_423,ImgReg2IN_422,ImgReg2IN_421,ImgReg2IN_420,
                      ImgReg2IN_419,ImgReg2IN_418,ImgReg2IN_417,ImgReg2IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState3N (.D ({DATA[431],DATA[430],DATA[429],
                      DATA[428],DATA[427],DATA[426],DATA[425],DATA[424],
                      DATA[423],DATA[422],DATA[421],DATA[420],DATA[419],
                      DATA[418],DATA[417],DATA[416]}), .EN (nx23624), .F ({
                      ImgReg3IN_431,ImgReg3IN_430,ImgReg3IN_429,ImgReg3IN_428,
                      ImgReg3IN_427,ImgReg3IN_426,ImgReg3IN_425,ImgReg3IN_424,
                      ImgReg3IN_423,ImgReg3IN_422,ImgReg3IN_421,ImgReg3IN_420,
                      ImgReg3IN_419,ImgReg3IN_418,ImgReg3IN_417,ImgReg3IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState4N (.D ({DATA[431],DATA[430],DATA[429],
                      DATA[428],DATA[427],DATA[426],DATA[425],DATA[424],
                      DATA[423],DATA[422],DATA[421],DATA[420],DATA[419],
                      DATA[418],DATA[417],DATA[416]}), .EN (nx23612), .F ({
                      ImgReg4IN_431,ImgReg4IN_430,ImgReg4IN_429,ImgReg4IN_428,
                      ImgReg4IN_427,ImgReg4IN_426,ImgReg4IN_425,ImgReg4IN_424,
                      ImgReg4IN_423,ImgReg4IN_422,ImgReg4IN_421,ImgReg4IN_420,
                      ImgReg4IN_419,ImgReg4IN_418,ImgReg4IN_417,ImgReg4IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState5N (.D ({DATA[431],DATA[430],DATA[429],
                      DATA[428],DATA[427],DATA[426],DATA[425],DATA[424],
                      DATA[423],DATA[422],DATA[421],DATA[420],DATA[419],
                      DATA[418],DATA[417],DATA[416]}), .EN (nx23600), .F ({
                      ImgReg5IN_431,ImgReg5IN_430,ImgReg5IN_429,ImgReg5IN_428,
                      ImgReg5IN_427,ImgReg5IN_426,ImgReg5IN_425,ImgReg5IN_424,
                      ImgReg5IN_423,ImgReg5IN_422,ImgReg5IN_421,ImgReg5IN_420,
                      ImgReg5IN_419,ImgReg5IN_418,ImgReg5IN_417,ImgReg5IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState0U (.D ({OutputImg1[431],OutputImg1[430],
                      OutputImg1[429],OutputImg1[428],OutputImg1[427],
                      OutputImg1[426],OutputImg1[425],OutputImg1[424],
                      OutputImg1[423],OutputImg1[422],OutputImg1[421],
                      OutputImg1[420],OutputImg1[419],OutputImg1[418],
                      OutputImg1[417],OutputImg1[416]}), .EN (nx23822), .F ({
                      ImgReg0IN_431,ImgReg0IN_430,ImgReg0IN_429,ImgReg0IN_428,
                      ImgReg0IN_427,ImgReg0IN_426,ImgReg0IN_425,ImgReg0IN_424,
                      ImgReg0IN_423,ImgReg0IN_422,ImgReg0IN_421,ImgReg0IN_420,
                      ImgReg0IN_419,ImgReg0IN_418,ImgReg0IN_417,ImgReg0IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState1U (.D ({OutputImg2[431],OutputImg2[430],
                      OutputImg2[429],OutputImg2[428],OutputImg2[427],
                      OutputImg2[426],OutputImg2[425],OutputImg2[424],
                      OutputImg2[423],OutputImg2[422],OutputImg2[421],
                      OutputImg2[420],OutputImg2[419],OutputImg2[418],
                      OutputImg2[417],OutputImg2[416]}), .EN (nx23822), .F ({
                      ImgReg1IN_431,ImgReg1IN_430,ImgReg1IN_429,ImgReg1IN_428,
                      ImgReg1IN_427,ImgReg1IN_426,ImgReg1IN_425,ImgReg1IN_424,
                      ImgReg1IN_423,ImgReg1IN_422,ImgReg1IN_421,ImgReg1IN_420,
                      ImgReg1IN_419,ImgReg1IN_418,ImgReg1IN_417,ImgReg1IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState2U (.D ({OutputImg3[431],OutputImg3[430],
                      OutputImg3[429],OutputImg3[428],OutputImg3[427],
                      OutputImg3[426],OutputImg3[425],OutputImg3[424],
                      OutputImg3[423],OutputImg3[422],OutputImg3[421],
                      OutputImg3[420],OutputImg3[419],OutputImg3[418],
                      OutputImg3[417],OutputImg3[416]}), .EN (nx23822), .F ({
                      ImgReg2IN_431,ImgReg2IN_430,ImgReg2IN_429,ImgReg2IN_428,
                      ImgReg2IN_427,ImgReg2IN_426,ImgReg2IN_425,ImgReg2IN_424,
                      ImgReg2IN_423,ImgReg2IN_422,ImgReg2IN_421,ImgReg2IN_420,
                      ImgReg2IN_419,ImgReg2IN_418,ImgReg2IN_417,ImgReg2IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState3U (.D ({OutputImg4[431],OutputImg4[430],
                      OutputImg4[429],OutputImg4[428],OutputImg4[427],
                      OutputImg4[426],OutputImg4[425],OutputImg4[424],
                      OutputImg4[423],OutputImg4[422],OutputImg4[421],
                      OutputImg4[420],OutputImg4[419],OutputImg4[418],
                      OutputImg4[417],OutputImg4[416]}), .EN (nx23824), .F ({
                      ImgReg3IN_431,ImgReg3IN_430,ImgReg3IN_429,ImgReg3IN_428,
                      ImgReg3IN_427,ImgReg3IN_426,ImgReg3IN_425,ImgReg3IN_424,
                      ImgReg3IN_423,ImgReg3IN_422,ImgReg3IN_421,ImgReg3IN_420,
                      ImgReg3IN_419,ImgReg3IN_418,ImgReg3IN_417,ImgReg3IN_416})
                      ) ;
    triStateBuffer_16 loop3_26_TriState4U (.D ({OutputImg5[431],OutputImg5[430],
                      OutputImg5[429],OutputImg5[428],OutputImg5[427],
                      OutputImg5[426],OutputImg5[425],OutputImg5[424],
                      OutputImg5[423],OutputImg5[422],OutputImg5[421],
                      OutputImg5[420],OutputImg5[419],OutputImg5[418],
                      OutputImg5[417],OutputImg5[416]}), .EN (nx23824), .F ({
                      ImgReg4IN_431,ImgReg4IN_430,ImgReg4IN_429,ImgReg4IN_428,
                      ImgReg4IN_427,ImgReg4IN_426,ImgReg4IN_425,ImgReg4IN_424,
                      ImgReg4IN_423,ImgReg4IN_422,ImgReg4IN_421,ImgReg4IN_420,
                      ImgReg4IN_419,ImgReg4IN_418,ImgReg4IN_417,ImgReg4IN_416})
                      ) ;
    nBitRegister_16 loop3_26_reg1 (.D ({ImgReg0IN_431,ImgReg0IN_430,
                    ImgReg0IN_429,ImgReg0IN_428,ImgReg0IN_427,ImgReg0IN_426,
                    ImgReg0IN_425,ImgReg0IN_424,ImgReg0IN_423,ImgReg0IN_422,
                    ImgReg0IN_421,ImgReg0IN_420,ImgReg0IN_419,ImgReg0IN_418,
                    ImgReg0IN_417,ImgReg0IN_416}), .CLK (nx23984), .RST (RST), .EN (
                    nx23724), .Q ({OutputImg0[431],OutputImg0[430],
                    OutputImg0[429],OutputImg0[428],OutputImg0[427],
                    OutputImg0[426],OutputImg0[425],OutputImg0[424],
                    OutputImg0[423],OutputImg0[422],OutputImg0[421],
                    OutputImg0[420],OutputImg0[419],OutputImg0[418],
                    OutputImg0[417],OutputImg0[416]})) ;
    nBitRegister_16 loop3_26_reg2 (.D ({ImgReg1IN_431,ImgReg1IN_430,
                    ImgReg1IN_429,ImgReg1IN_428,ImgReg1IN_427,ImgReg1IN_426,
                    ImgReg1IN_425,ImgReg1IN_424,ImgReg1IN_423,ImgReg1IN_422,
                    ImgReg1IN_421,ImgReg1IN_420,ImgReg1IN_419,ImgReg1IN_418,
                    ImgReg1IN_417,ImgReg1IN_416}), .CLK (nx23986), .RST (RST), .EN (
                    nx23734), .Q ({OutputImg1[431],OutputImg1[430],
                    OutputImg1[429],OutputImg1[428],OutputImg1[427],
                    OutputImg1[426],OutputImg1[425],OutputImg1[424],
                    OutputImg1[423],OutputImg1[422],OutputImg1[421],
                    OutputImg1[420],OutputImg1[419],OutputImg1[418],
                    OutputImg1[417],OutputImg1[416]})) ;
    nBitRegister_16 loop3_26_reg3 (.D ({ImgReg2IN_431,ImgReg2IN_430,
                    ImgReg2IN_429,ImgReg2IN_428,ImgReg2IN_427,ImgReg2IN_426,
                    ImgReg2IN_425,ImgReg2IN_424,ImgReg2IN_423,ImgReg2IN_422,
                    ImgReg2IN_421,ImgReg2IN_420,ImgReg2IN_419,ImgReg2IN_418,
                    ImgReg2IN_417,ImgReg2IN_416}), .CLK (nx23986), .RST (RST), .EN (
                    nx23744), .Q ({OutputImg2[431],OutputImg2[430],
                    OutputImg2[429],OutputImg2[428],OutputImg2[427],
                    OutputImg2[426],OutputImg2[425],OutputImg2[424],
                    OutputImg2[423],OutputImg2[422],OutputImg2[421],
                    OutputImg2[420],OutputImg2[419],OutputImg2[418],
                    OutputImg2[417],OutputImg2[416]})) ;
    nBitRegister_16 loop3_26_reg4 (.D ({ImgReg3IN_431,ImgReg3IN_430,
                    ImgReg3IN_429,ImgReg3IN_428,ImgReg3IN_427,ImgReg3IN_426,
                    ImgReg3IN_425,ImgReg3IN_424,ImgReg3IN_423,ImgReg3IN_422,
                    ImgReg3IN_421,ImgReg3IN_420,ImgReg3IN_419,ImgReg3IN_418,
                    ImgReg3IN_417,ImgReg3IN_416}), .CLK (nx23988), .RST (RST), .EN (
                    nx23754), .Q ({OutputImg3[431],OutputImg3[430],
                    OutputImg3[429],OutputImg3[428],OutputImg3[427],
                    OutputImg3[426],OutputImg3[425],OutputImg3[424],
                    OutputImg3[423],OutputImg3[422],OutputImg3[421],
                    OutputImg3[420],OutputImg3[419],OutputImg3[418],
                    OutputImg3[417],OutputImg3[416]})) ;
    nBitRegister_16 loop3_26_reg5 (.D ({ImgReg4IN_431,ImgReg4IN_430,
                    ImgReg4IN_429,ImgReg4IN_428,ImgReg4IN_427,ImgReg4IN_426,
                    ImgReg4IN_425,ImgReg4IN_424,ImgReg4IN_423,ImgReg4IN_422,
                    ImgReg4IN_421,ImgReg4IN_420,ImgReg4IN_419,ImgReg4IN_418,
                    ImgReg4IN_417,ImgReg4IN_416}), .CLK (nx23988), .RST (RST), .EN (
                    nx23764), .Q ({OutputImg4[431],OutputImg4[430],
                    OutputImg4[429],OutputImg4[428],OutputImg4[427],
                    OutputImg4[426],OutputImg4[425],OutputImg4[424],
                    OutputImg4[423],OutputImg4[422],OutputImg4[421],
                    OutputImg4[420],OutputImg4[419],OutputImg4[418],
                    OutputImg4[417],OutputImg4[416]})) ;
    nBitRegister_16 loop3_26_reg6 (.D ({ImgReg5IN_431,ImgReg5IN_430,
                    ImgReg5IN_429,ImgReg5IN_428,ImgReg5IN_427,ImgReg5IN_426,
                    ImgReg5IN_425,ImgReg5IN_424,ImgReg5IN_423,ImgReg5IN_422,
                    ImgReg5IN_421,ImgReg5IN_420,ImgReg5IN_419,ImgReg5IN_418,
                    ImgReg5IN_417,ImgReg5IN_416}), .CLK (nx23990), .RST (RST), .EN (
                    nx23774), .Q ({OutputImg5[431],OutputImg5[430],
                    OutputImg5[429],OutputImg5[428],OutputImg5[427],
                    OutputImg5[426],OutputImg5[425],OutputImg5[424],
                    OutputImg5[423],OutputImg5[422],OutputImg5[421],
                    OutputImg5[420],OutputImg5[419],OutputImg5[418],
                    OutputImg5[417],OutputImg5[416]})) ;
    triStateBuffer_16 TriState00L (.D ({OutputImg0[15],OutputImg0[14],
                      OutputImg0[13],OutputImg0[12],OutputImg0[11],
                      OutputImg0[10],OutputImg0[9],OutputImg0[8],OutputImg0[7],
                      OutputImg0[6],OutputImg0[5],OutputImg0[4],OutputImg0[3],
                      OutputImg0[2],OutputImg0[1],OutputImg0[0]}), .EN (nx23712)
                      , .F ({ImgReg0IN_447,ImgReg0IN_446,ImgReg0IN_445,
                      ImgReg0IN_444,ImgReg0IN_443,ImgReg0IN_442,ImgReg0IN_441,
                      ImgReg0IN_440,ImgReg0IN_439,ImgReg0IN_438,ImgReg0IN_437,
                      ImgReg0IN_436,ImgReg0IN_435,ImgReg0IN_434,ImgReg0IN_433,
                      ImgReg0IN_432})) ;
    triStateBuffer_16 TriState11L (.D ({OutputImg1[15],OutputImg1[14],
                      OutputImg1[13],OutputImg1[12],OutputImg1[11],
                      OutputImg1[10],OutputImg1[9],OutputImg1[8],OutputImg1[7],
                      OutputImg1[6],OutputImg1[5],OutputImg1[4],OutputImg1[3],
                      OutputImg1[2],OutputImg1[1],OutputImg1[0]}), .EN (nx23712)
                      , .F ({ImgReg1IN_447,ImgReg1IN_446,ImgReg1IN_445,
                      ImgReg1IN_444,ImgReg1IN_443,ImgReg1IN_442,ImgReg1IN_441,
                      ImgReg1IN_440,ImgReg1IN_439,ImgReg1IN_438,ImgReg1IN_437,
                      ImgReg1IN_436,ImgReg1IN_435,ImgReg1IN_434,ImgReg1IN_433,
                      ImgReg1IN_432})) ;
    triStateBuffer_16 TriState22L (.D ({OutputImg2[15],OutputImg2[14],
                      OutputImg2[13],OutputImg2[12],OutputImg2[11],
                      OutputImg2[10],OutputImg2[9],OutputImg2[8],OutputImg2[7],
                      OutputImg2[6],OutputImg2[5],OutputImg2[4],OutputImg2[3],
                      OutputImg2[2],OutputImg2[1],OutputImg2[0]}), .EN (nx23712)
                      , .F ({ImgReg2IN_447,ImgReg2IN_446,ImgReg2IN_445,
                      ImgReg2IN_444,ImgReg2IN_443,ImgReg2IN_442,ImgReg2IN_441,
                      ImgReg2IN_440,ImgReg2IN_439,ImgReg2IN_438,ImgReg2IN_437,
                      ImgReg2IN_436,ImgReg2IN_435,ImgReg2IN_434,ImgReg2IN_433,
                      ImgReg2IN_432})) ;
    triStateBuffer_16 TriState33L (.D ({OutputImg3[15],OutputImg3[14],
                      OutputImg3[13],OutputImg3[12],OutputImg3[11],
                      OutputImg3[10],OutputImg3[9],OutputImg3[8],OutputImg3[7],
                      OutputImg3[6],OutputImg3[5],OutputImg3[4],OutputImg3[3],
                      OutputImg3[2],OutputImg3[1],OutputImg3[0]}), .EN (nx23712)
                      , .F ({ImgReg3IN_447,ImgReg3IN_446,ImgReg3IN_445,
                      ImgReg3IN_444,ImgReg3IN_443,ImgReg3IN_442,ImgReg3IN_441,
                      ImgReg3IN_440,ImgReg3IN_439,ImgReg3IN_438,ImgReg3IN_437,
                      ImgReg3IN_436,ImgReg3IN_435,ImgReg3IN_434,ImgReg3IN_433,
                      ImgReg3IN_432})) ;
    triStateBuffer_16 TriState44L (.D ({OutputImg4[15],OutputImg4[14],
                      OutputImg4[13],OutputImg4[12],OutputImg4[11],
                      OutputImg4[10],OutputImg4[9],OutputImg4[8],OutputImg4[7],
                      OutputImg4[6],OutputImg4[5],OutputImg4[4],OutputImg4[3],
                      OutputImg4[2],OutputImg4[1],OutputImg4[0]}), .EN (nx23712)
                      , .F ({ImgReg4IN_447,ImgReg4IN_446,ImgReg4IN_445,
                      ImgReg4IN_444,ImgReg4IN_443,ImgReg4IN_442,ImgReg4IN_441,
                      ImgReg4IN_440,ImgReg4IN_439,ImgReg4IN_438,ImgReg4IN_437,
                      ImgReg4IN_436,ImgReg4IN_435,ImgReg4IN_434,ImgReg4IN_433,
                      ImgReg4IN_432})) ;
    triStateBuffer_16 TriState55L (.D ({OutputImg5[15],OutputImg5[14],
                      OutputImg5[13],OutputImg5[12],OutputImg5[11],
                      OutputImg5[10],OutputImg5[9],OutputImg5[8],OutputImg5[7],
                      OutputImg5[6],OutputImg5[5],OutputImg5[4],OutputImg5[3],
                      OutputImg5[2],OutputImg5[1],OutputImg5[0]}), .EN (nx23712)
                      , .F ({ImgReg5IN_447,ImgReg5IN_446,ImgReg5IN_445,
                      ImgReg5IN_444,ImgReg5IN_443,ImgReg5IN_442,ImgReg5IN_441,
                      ImgReg5IN_440,ImgReg5IN_439,ImgReg5IN_438,ImgReg5IN_437,
                      ImgReg5IN_436,ImgReg5IN_435,ImgReg5IN_434,ImgReg5IN_433,
                      ImgReg5IN_432})) ;
    triStateBuffer_16 TriState00N (.D ({DATA[447],DATA[446],DATA[445],DATA[444],
                      DATA[443],DATA[442],DATA[441],DATA[440],DATA[439],
                      DATA[438],DATA[437],DATA[436],DATA[435],DATA[434],
                      DATA[433],DATA[432]}), .EN (nx23660), .F ({ImgReg0IN_447,
                      ImgReg0IN_446,ImgReg0IN_445,ImgReg0IN_444,ImgReg0IN_443,
                      ImgReg0IN_442,ImgReg0IN_441,ImgReg0IN_440,ImgReg0IN_439,
                      ImgReg0IN_438,ImgReg0IN_437,ImgReg0IN_436,ImgReg0IN_435,
                      ImgReg0IN_434,ImgReg0IN_433,ImgReg0IN_432})) ;
    triStateBuffer_16 TriState11N (.D ({DATA[447],DATA[446],DATA[445],DATA[444],
                      DATA[443],DATA[442],DATA[441],DATA[440],DATA[439],
                      DATA[438],DATA[437],DATA[436],DATA[435],DATA[434],
                      DATA[433],DATA[432]}), .EN (nx23648), .F ({ImgReg1IN_447,
                      ImgReg1IN_446,ImgReg1IN_445,ImgReg1IN_444,ImgReg1IN_443,
                      ImgReg1IN_442,ImgReg1IN_441,ImgReg1IN_440,ImgReg1IN_439,
                      ImgReg1IN_438,ImgReg1IN_437,ImgReg1IN_436,ImgReg1IN_435,
                      ImgReg1IN_434,ImgReg1IN_433,ImgReg1IN_432})) ;
    triStateBuffer_16 TriState22N (.D ({DATA[447],DATA[446],DATA[445],DATA[444],
                      DATA[443],DATA[442],DATA[441],DATA[440],DATA[439],
                      DATA[438],DATA[437],DATA[436],DATA[435],DATA[434],
                      DATA[433],DATA[432]}), .EN (nx23636), .F ({ImgReg2IN_447,
                      ImgReg2IN_446,ImgReg2IN_445,ImgReg2IN_444,ImgReg2IN_443,
                      ImgReg2IN_442,ImgReg2IN_441,ImgReg2IN_440,ImgReg2IN_439,
                      ImgReg2IN_438,ImgReg2IN_437,ImgReg2IN_436,ImgReg2IN_435,
                      ImgReg2IN_434,ImgReg2IN_433,ImgReg2IN_432})) ;
    triStateBuffer_16 TriState33N (.D ({DATA[447],DATA[446],DATA[445],DATA[444],
                      DATA[443],DATA[442],DATA[441],DATA[440],DATA[439],
                      DATA[438],DATA[437],DATA[436],DATA[435],DATA[434],
                      DATA[433],DATA[432]}), .EN (nx23624), .F ({ImgReg3IN_447,
                      ImgReg3IN_446,ImgReg3IN_445,ImgReg3IN_444,ImgReg3IN_443,
                      ImgReg3IN_442,ImgReg3IN_441,ImgReg3IN_440,ImgReg3IN_439,
                      ImgReg3IN_438,ImgReg3IN_437,ImgReg3IN_436,ImgReg3IN_435,
                      ImgReg3IN_434,ImgReg3IN_433,ImgReg3IN_432})) ;
    triStateBuffer_16 TriState44N (.D ({DATA[447],DATA[446],DATA[445],DATA[444],
                      DATA[443],DATA[442],DATA[441],DATA[440],DATA[439],
                      DATA[438],DATA[437],DATA[436],DATA[435],DATA[434],
                      DATA[433],DATA[432]}), .EN (nx23612), .F ({ImgReg4IN_447,
                      ImgReg4IN_446,ImgReg4IN_445,ImgReg4IN_444,ImgReg4IN_443,
                      ImgReg4IN_442,ImgReg4IN_441,ImgReg4IN_440,ImgReg4IN_439,
                      ImgReg4IN_438,ImgReg4IN_437,ImgReg4IN_436,ImgReg4IN_435,
                      ImgReg4IN_434,ImgReg4IN_433,ImgReg4IN_432})) ;
    triStateBuffer_16 TriState55N (.D ({DATA[447],DATA[446],DATA[445],DATA[444],
                      DATA[443],DATA[442],DATA[441],DATA[440],DATA[439],
                      DATA[438],DATA[437],DATA[436],DATA[435],DATA[434],
                      DATA[433],DATA[432]}), .EN (nx23600), .F ({ImgReg5IN_447,
                      ImgReg5IN_446,ImgReg5IN_445,ImgReg5IN_444,ImgReg5IN_443,
                      ImgReg5IN_442,ImgReg5IN_441,ImgReg5IN_440,ImgReg5IN_439,
                      ImgReg5IN_438,ImgReg5IN_437,ImgReg5IN_436,ImgReg5IN_435,
                      ImgReg5IN_434,ImgReg5IN_433,ImgReg5IN_432})) ;
    triStateBuffer_16 TriState00U (.D ({OutputImg1[447],OutputImg1[446],
                      OutputImg1[445],OutputImg1[444],OutputImg1[443],
                      OutputImg1[442],OutputImg1[441],OutputImg1[440],
                      OutputImg1[439],OutputImg1[438],OutputImg1[437],
                      OutputImg1[436],OutputImg1[435],OutputImg1[434],
                      OutputImg1[433],OutputImg1[432]}), .EN (nx23824), .F ({
                      ImgReg0IN_447,ImgReg0IN_446,ImgReg0IN_445,ImgReg0IN_444,
                      ImgReg0IN_443,ImgReg0IN_442,ImgReg0IN_441,ImgReg0IN_440,
                      ImgReg0IN_439,ImgReg0IN_438,ImgReg0IN_437,ImgReg0IN_436,
                      ImgReg0IN_435,ImgReg0IN_434,ImgReg0IN_433,ImgReg0IN_432})
                      ) ;
    triStateBuffer_16 TriState11U (.D ({OutputImg2[447],OutputImg2[446],
                      OutputImg2[445],OutputImg2[444],OutputImg2[443],
                      OutputImg2[442],OutputImg2[441],OutputImg2[440],
                      OutputImg2[439],OutputImg2[438],OutputImg2[437],
                      OutputImg2[436],OutputImg2[435],OutputImg2[434],
                      OutputImg2[433],OutputImg2[432]}), .EN (nx23824), .F ({
                      ImgReg1IN_447,ImgReg1IN_446,ImgReg1IN_445,ImgReg1IN_444,
                      ImgReg1IN_443,ImgReg1IN_442,ImgReg1IN_441,ImgReg1IN_440,
                      ImgReg1IN_439,ImgReg1IN_438,ImgReg1IN_437,ImgReg1IN_436,
                      ImgReg1IN_435,ImgReg1IN_434,ImgReg1IN_433,ImgReg1IN_432})
                      ) ;
    triStateBuffer_16 TriState22U (.D ({OutputImg3[447],OutputImg3[446],
                      OutputImg3[445],OutputImg3[444],OutputImg3[443],
                      OutputImg3[442],OutputImg3[441],OutputImg3[440],
                      OutputImg3[439],OutputImg3[438],OutputImg3[437],
                      OutputImg3[436],OutputImg3[435],OutputImg3[434],
                      OutputImg3[433],OutputImg3[432]}), .EN (nx23824), .F ({
                      ImgReg2IN_447,ImgReg2IN_446,ImgReg2IN_445,ImgReg2IN_444,
                      ImgReg2IN_443,ImgReg2IN_442,ImgReg2IN_441,ImgReg2IN_440,
                      ImgReg2IN_439,ImgReg2IN_438,ImgReg2IN_437,ImgReg2IN_436,
                      ImgReg2IN_435,ImgReg2IN_434,ImgReg2IN_433,ImgReg2IN_432})
                      ) ;
    triStateBuffer_16 TriState33U (.D ({OutputImg4[447],OutputImg4[446],
                      OutputImg4[445],OutputImg4[444],OutputImg4[443],
                      OutputImg4[442],OutputImg4[441],OutputImg4[440],
                      OutputImg4[439],OutputImg4[438],OutputImg4[437],
                      OutputImg4[436],OutputImg4[435],OutputImg4[434],
                      OutputImg4[433],OutputImg4[432]}), .EN (nx23824), .F ({
                      ImgReg3IN_447,ImgReg3IN_446,ImgReg3IN_445,ImgReg3IN_444,
                      ImgReg3IN_443,ImgReg3IN_442,ImgReg3IN_441,ImgReg3IN_440,
                      ImgReg3IN_439,ImgReg3IN_438,ImgReg3IN_437,ImgReg3IN_436,
                      ImgReg3IN_435,ImgReg3IN_434,ImgReg3IN_433,ImgReg3IN_432})
                      ) ;
    triStateBuffer_16 TriState44U (.D ({OutputImg5[447],OutputImg5[446],
                      OutputImg5[445],OutputImg5[444],OutputImg5[443],
                      OutputImg5[442],OutputImg5[441],OutputImg5[440],
                      OutputImg5[439],OutputImg5[438],OutputImg5[437],
                      OutputImg5[436],OutputImg5[435],OutputImg5[434],
                      OutputImg5[433],OutputImg5[432]}), .EN (nx23824), .F ({
                      ImgReg4IN_447,ImgReg4IN_446,ImgReg4IN_445,ImgReg4IN_444,
                      ImgReg4IN_443,ImgReg4IN_442,ImgReg4IN_441,ImgReg4IN_440,
                      ImgReg4IN_439,ImgReg4IN_438,ImgReg4IN_437,ImgReg4IN_436,
                      ImgReg4IN_435,ImgReg4IN_434,ImgReg4IN_433,ImgReg4IN_432})
                      ) ;
    nBitRegister_16 reg11 (.D ({ImgReg0IN_447,ImgReg0IN_446,ImgReg0IN_445,
                    ImgReg0IN_444,ImgReg0IN_443,ImgReg0IN_442,ImgReg0IN_441,
                    ImgReg0IN_440,ImgReg0IN_439,ImgReg0IN_438,ImgReg0IN_437,
                    ImgReg0IN_436,ImgReg0IN_435,ImgReg0IN_434,ImgReg0IN_433,
                    ImgReg0IN_432}), .CLK (nx23990), .RST (RST), .EN (nx23724), 
                    .Q ({OutputImg0[447],OutputImg0[446],OutputImg0[445],
                    OutputImg0[444],OutputImg0[443],OutputImg0[442],
                    OutputImg0[441],OutputImg0[440],OutputImg0[439],
                    OutputImg0[438],OutputImg0[437],OutputImg0[436],
                    OutputImg0[435],OutputImg0[434],OutputImg0[433],
                    OutputImg0[432]})) ;
    nBitRegister_16 reg22 (.D ({ImgReg1IN_447,ImgReg1IN_446,ImgReg1IN_445,
                    ImgReg1IN_444,ImgReg1IN_443,ImgReg1IN_442,ImgReg1IN_441,
                    ImgReg1IN_440,ImgReg1IN_439,ImgReg1IN_438,ImgReg1IN_437,
                    ImgReg1IN_436,ImgReg1IN_435,ImgReg1IN_434,ImgReg1IN_433,
                    ImgReg1IN_432}), .CLK (nx23992), .RST (RST), .EN (nx23734), 
                    .Q ({OutputImg1[447],OutputImg1[446],OutputImg1[445],
                    OutputImg1[444],OutputImg1[443],OutputImg1[442],
                    OutputImg1[441],OutputImg1[440],OutputImg1[439],
                    OutputImg1[438],OutputImg1[437],OutputImg1[436],
                    OutputImg1[435],OutputImg1[434],OutputImg1[433],
                    OutputImg1[432]})) ;
    nBitRegister_16 reg33 (.D ({ImgReg2IN_447,ImgReg2IN_446,ImgReg2IN_445,
                    ImgReg2IN_444,ImgReg2IN_443,ImgReg2IN_442,ImgReg2IN_441,
                    ImgReg2IN_440,ImgReg2IN_439,ImgReg2IN_438,ImgReg2IN_437,
                    ImgReg2IN_436,ImgReg2IN_435,ImgReg2IN_434,ImgReg2IN_433,
                    ImgReg2IN_432}), .CLK (nx23992), .RST (RST), .EN (nx23744), 
                    .Q ({OutputImg2[447],OutputImg2[446],OutputImg2[445],
                    OutputImg2[444],OutputImg2[443],OutputImg2[442],
                    OutputImg2[441],OutputImg2[440],OutputImg2[439],
                    OutputImg2[438],OutputImg2[437],OutputImg2[436],
                    OutputImg2[435],OutputImg2[434],OutputImg2[433],
                    OutputImg2[432]})) ;
    nBitRegister_16 reg44 (.D ({ImgReg3IN_447,ImgReg3IN_446,ImgReg3IN_445,
                    ImgReg3IN_444,ImgReg3IN_443,ImgReg3IN_442,ImgReg3IN_441,
                    ImgReg3IN_440,ImgReg3IN_439,ImgReg3IN_438,ImgReg3IN_437,
                    ImgReg3IN_436,ImgReg3IN_435,ImgReg3IN_434,ImgReg3IN_433,
                    ImgReg3IN_432}), .CLK (nx23994), .RST (RST), .EN (nx23754), 
                    .Q ({OutputImg3[447],OutputImg3[446],OutputImg3[445],
                    OutputImg3[444],OutputImg3[443],OutputImg3[442],
                    OutputImg3[441],OutputImg3[440],OutputImg3[439],
                    OutputImg3[438],OutputImg3[437],OutputImg3[436],
                    OutputImg3[435],OutputImg3[434],OutputImg3[433],
                    OutputImg3[432]})) ;
    nBitRegister_16 reg55 (.D ({ImgReg4IN_447,ImgReg4IN_446,ImgReg4IN_445,
                    ImgReg4IN_444,ImgReg4IN_443,ImgReg4IN_442,ImgReg4IN_441,
                    ImgReg4IN_440,ImgReg4IN_439,ImgReg4IN_438,ImgReg4IN_437,
                    ImgReg4IN_436,ImgReg4IN_435,ImgReg4IN_434,ImgReg4IN_433,
                    ImgReg4IN_432}), .CLK (nx23994), .RST (RST), .EN (nx23764), 
                    .Q ({OutputImg4[447],OutputImg4[446],OutputImg4[445],
                    OutputImg4[444],OutputImg4[443],OutputImg4[442],
                    OutputImg4[441],OutputImg4[440],OutputImg4[439],
                    OutputImg4[438],OutputImg4[437],OutputImg4[436],
                    OutputImg4[435],OutputImg4[434],OutputImg4[433],
                    OutputImg4[432]})) ;
    nBitRegister_16 reg66 (.D ({ImgReg5IN_447,ImgReg5IN_446,ImgReg5IN_445,
                    ImgReg5IN_444,ImgReg5IN_443,ImgReg5IN_442,ImgReg5IN_441,
                    ImgReg5IN_440,ImgReg5IN_439,ImgReg5IN_438,ImgReg5IN_437,
                    ImgReg5IN_436,ImgReg5IN_435,ImgReg5IN_434,ImgReg5IN_433,
                    ImgReg5IN_432}), .CLK (nx23996), .RST (RST), .EN (nx23774), 
                    .Q ({OutputImg5[447],OutputImg5[446],OutputImg5[445],
                    OutputImg5[444],OutputImg5[443],OutputImg5[442],
                    OutputImg5[441],OutputImg5[440],OutputImg5[439],
                    OutputImg5[438],OutputImg5[437],OutputImg5[436],
                    OutputImg5[435],OutputImg5[434],OutputImg5[433],
                    OutputImg5[432]})) ;
    inv01 ix23555 (.Y (NOT_ImgIndic_0), .A (ImgIndic[0])) ;
    fake_gnd ix23530 (.Y (firstOperand_15)) ;
    fake_vcc ix23528 (.Y (PWR)) ;
    or02 ix5 (.Y (TriImgLeftEn), .A0 (nx2), .A1 (current_state[10])) ;
    and03 ix3 (.Y (nx2), .A0 (ACK), .A1 (WI), .A2 (current_state[8])) ;
    oai21 ix43 (.Y (TriImgRegEn), .A0 (ImgIndic[0]), .A1 (nx34), .B0 (nx23568)
          ) ;
    nand02 ix35 (.Y (nx34), .A0 (current_state[7]), .A1 (ACK)) ;
    nor02ii ix29 (.Y (cEnable), .A0 (nx23573), .A1 (ACK)) ;
    nor04 ix23574 (.Y (nx23573), .A0 (current_state[2]), .A1 (current_state[3])
          , .A2 (nx20), .A3 (current_state[4])) ;
    or02 ix21 (.Y (nx20), .A0 (current_state[5]), .A1 (current_state[6])) ;
    or02 ix45 (.Y (cReset), .A0 (RST), .A1 (current_state[12])) ;
    oai21 ix51 (.Y (IndRst), .A0 (nx23998), .A1 (dontTrust), .B0 (nx23580)) ;
    inv01 ix23581 (.Y (nx23580), .A (RST)) ;
    oai21 ix63 (.Y (TriAddEn), .A0 (nx23583), .A1 (ImgIndic[0]), .B0 (nx23573)
          ) ;
    inv01 ix23584 (.Y (nx23583), .A (current_state[7])) ;
    dffr reg_DFFCLK_dup_0 (.Q (DFFCLK), .QB (\$dummy [4]), .D (PWR), .CLK (
         nx23830), .R (nx34)) ;
    inv01 ix23569 (.Y (nx23568), .A (cEnable)) ;
    inv01 ix23591 (.Y (nx23592), .A (ImgEn[5])) ;
    inv01 ix23593 (.Y (nx23594), .A (nx23592)) ;
    inv01 ix23595 (.Y (nx23596), .A (nx23592)) ;
    inv01 ix23597 (.Y (nx23598), .A (nx23592)) ;
    inv01 ix23599 (.Y (nx23600), .A (nx23592)) ;
    inv01 ix23603 (.Y (nx23604), .A (ImgEn[4])) ;
    inv01 ix23605 (.Y (nx23606), .A (nx23604)) ;
    inv01 ix23607 (.Y (nx23608), .A (nx23604)) ;
    inv01 ix23609 (.Y (nx23610), .A (nx23604)) ;
    inv01 ix23611 (.Y (nx23612), .A (nx23604)) ;
    inv01 ix23615 (.Y (nx23616), .A (ImgEn[3])) ;
    inv01 ix23617 (.Y (nx23618), .A (nx23616)) ;
    inv01 ix23619 (.Y (nx23620), .A (nx23616)) ;
    inv01 ix23621 (.Y (nx23622), .A (nx23616)) ;
    inv01 ix23623 (.Y (nx23624), .A (nx23616)) ;
    inv01 ix23627 (.Y (nx23628), .A (ImgEn[2])) ;
    inv01 ix23629 (.Y (nx23630), .A (nx23628)) ;
    inv01 ix23631 (.Y (nx23632), .A (nx23628)) ;
    inv01 ix23633 (.Y (nx23634), .A (nx23628)) ;
    inv01 ix23635 (.Y (nx23636), .A (nx23628)) ;
    inv01 ix23639 (.Y (nx23640), .A (ImgEn[1])) ;
    inv01 ix23641 (.Y (nx23642), .A (nx23640)) ;
    inv01 ix23643 (.Y (nx23644), .A (nx23640)) ;
    inv01 ix23645 (.Y (nx23646), .A (nx23640)) ;
    inv01 ix23647 (.Y (nx23648), .A (nx23640)) ;
    inv01 ix23651 (.Y (nx23652), .A (ImgEn[0])) ;
    inv01 ix23653 (.Y (nx23654), .A (nx23652)) ;
    inv01 ix23655 (.Y (nx23656), .A (nx23652)) ;
    inv01 ix23657 (.Y (nx23658), .A (nx23652)) ;
    inv01 ix23659 (.Y (nx23660), .A (nx23652)) ;
    inv01 ix23663 (.Y (nx23664), .A (TriImgLeftEn)) ;
    inv01 ix23665 (.Y (nx23666), .A (nx23776)) ;
    inv01 ix23667 (.Y (nx23668), .A (nx23776)) ;
    inv01 ix23669 (.Y (nx23670), .A (nx23776)) ;
    inv01 ix23671 (.Y (nx23672), .A (nx23776)) ;
    inv01 ix23673 (.Y (nx23674), .A (nx23776)) ;
    inv01 ix23675 (.Y (nx23676), .A (nx23776)) ;
    inv01 ix23677 (.Y (nx23678), .A (nx23776)) ;
    inv01 ix23679 (.Y (nx23680), .A (nx23778)) ;
    inv01 ix23681 (.Y (nx23682), .A (nx23778)) ;
    inv01 ix23683 (.Y (nx23684), .A (nx23778)) ;
    inv01 ix23685 (.Y (nx23686), .A (nx23778)) ;
    inv01 ix23687 (.Y (nx23688), .A (nx23778)) ;
    inv01 ix23689 (.Y (nx23690), .A (nx23778)) ;
    inv01 ix23691 (.Y (nx23692), .A (nx23778)) ;
    inv01 ix23693 (.Y (nx23694), .A (nx23780)) ;
    inv01 ix23695 (.Y (nx23696), .A (nx23780)) ;
    inv01 ix23697 (.Y (nx23698), .A (nx23780)) ;
    inv01 ix23699 (.Y (nx23700), .A (nx23780)) ;
    inv01 ix23701 (.Y (nx23702), .A (nx23780)) ;
    inv01 ix23703 (.Y (nx23704), .A (nx23780)) ;
    inv01 ix23705 (.Y (nx23706), .A (nx23780)) ;
    inv01 ix23707 (.Y (nx23708), .A (nx24006)) ;
    inv01 ix23709 (.Y (nx23710), .A (nx24006)) ;
    inv01 ix23711 (.Y (nx23712), .A (nx24006)) ;
    inv01 ix23717 (.Y (nx23718), .A (nx23716)) ;
    inv01 ix23719 (.Y (nx23720), .A (nx23716)) ;
    inv01 ix23721 (.Y (nx23722), .A (nx23716)) ;
    inv01 ix23723 (.Y (nx23724), .A (nx23716)) ;
    inv01 ix23727 (.Y (nx23728), .A (nx23726)) ;
    inv01 ix23729 (.Y (nx23730), .A (nx23726)) ;
    inv01 ix23731 (.Y (nx23732), .A (nx23726)) ;
    inv01 ix23733 (.Y (nx23734), .A (nx23726)) ;
    inv01 ix23737 (.Y (nx23738), .A (nx23736)) ;
    inv01 ix23739 (.Y (nx23740), .A (nx23736)) ;
    inv01 ix23741 (.Y (nx23742), .A (nx23736)) ;
    inv01 ix23743 (.Y (nx23744), .A (nx23736)) ;
    inv01 ix23747 (.Y (nx23748), .A (nx23746)) ;
    inv01 ix23749 (.Y (nx23750), .A (nx23746)) ;
    inv01 ix23751 (.Y (nx23752), .A (nx23746)) ;
    inv01 ix23753 (.Y (nx23754), .A (nx23746)) ;
    inv01 ix23757 (.Y (nx23758), .A (nx23756)) ;
    inv01 ix23759 (.Y (nx23760), .A (nx23756)) ;
    inv01 ix23761 (.Y (nx23762), .A (nx23756)) ;
    inv01 ix23763 (.Y (nx23764), .A (nx23756)) ;
    inv01 ix23767 (.Y (nx23768), .A (nx23766)) ;
    inv01 ix23769 (.Y (nx23770), .A (nx23766)) ;
    inv01 ix23771 (.Y (nx23772), .A (nx23766)) ;
    inv01 ix23773 (.Y (nx23774), .A (nx23766)) ;
    inv01 ix23775 (.Y (nx23776), .A (TriImgLeftEn)) ;
    inv01 ix23777 (.Y (nx23778), .A (TriImgLeftEn)) ;
    inv01 ix23779 (.Y (nx23780), .A (TriImgLeftEn)) ;
    and02 ix7 (.Y (nx23766), .A0 (nx24006), .A1 (nx23592)) ;
    and03 ix11 (.Y (nx23756), .A0 (nx24006), .A1 (nx23998), .A2 (nx23604)) ;
    and03 ix13 (.Y (nx23746), .A0 (nx24006), .A1 (nx23998), .A2 (nx23616)) ;
    and03 ix15 (.Y (nx23736), .A0 (nx24006), .A1 (nx23998), .A2 (nx23628)) ;
    and03 ix17 (.Y (nx23726), .A0 (nx23664), .A1 (nx23998), .A2 (nx23640)) ;
    and03 ix19 (.Y (nx23716), .A0 (nx23664), .A1 (nx23998), .A2 (nx23652)) ;
    inv01 ix23785 (.Y (nx23786), .A (nx23998)) ;
    inv01 ix23787 (.Y (nx23788), .A (nx24000)) ;
    inv01 ix23789 (.Y (nx23790), .A (nx24000)) ;
    inv01 ix23791 (.Y (nx23792), .A (nx24000)) ;
    inv01 ix23793 (.Y (nx23794), .A (nx24000)) ;
    inv01 ix23795 (.Y (nx23796), .A (nx24000)) ;
    inv01 ix23797 (.Y (nx23798), .A (nx24000)) ;
    inv01 ix23799 (.Y (nx23800), .A (nx24000)) ;
    inv01 ix23801 (.Y (nx23802), .A (nx24002)) ;
    inv01 ix23803 (.Y (nx23804), .A (nx24002)) ;
    inv01 ix23805 (.Y (nx23806), .A (nx24002)) ;
    inv01 ix23807 (.Y (nx23808), .A (nx24002)) ;
    inv01 ix23809 (.Y (nx23810), .A (nx24002)) ;
    inv01 ix23811 (.Y (nx23812), .A (nx24002)) ;
    inv01 ix23813 (.Y (nx23814), .A (nx24002)) ;
    inv01 ix23815 (.Y (nx23816), .A (nx24004)) ;
    inv01 ix23817 (.Y (nx23818), .A (nx24004)) ;
    inv01 ix23819 (.Y (nx23820), .A (nx24004)) ;
    inv01 ix23821 (.Y (nx23822), .A (nx24004)) ;
    inv01 ix23823 (.Y (nx23824), .A (nx24004)) ;
    inv02 ix23827 (.Y (nx23828), .A (nx24008)) ;
    inv02 ix23829 (.Y (nx23830), .A (nx24008)) ;
    inv02 ix23831 (.Y (nx23832), .A (nx24008)) ;
    inv02 ix23833 (.Y (nx23834), .A (nx24008)) ;
    inv02 ix23835 (.Y (nx23836), .A (nx24008)) ;
    inv02 ix23837 (.Y (nx23838), .A (nx24008)) ;
    inv02 ix23839 (.Y (nx23840), .A (nx24008)) ;
    inv02 ix23841 (.Y (nx23842), .A (nx24010)) ;
    inv02 ix23843 (.Y (nx23844), .A (nx24010)) ;
    inv02 ix23845 (.Y (nx23846), .A (nx24010)) ;
    inv02 ix23847 (.Y (nx23848), .A (nx24010)) ;
    inv02 ix23849 (.Y (nx23850), .A (nx24010)) ;
    inv02 ix23851 (.Y (nx23852), .A (nx24010)) ;
    inv02 ix23853 (.Y (nx23854), .A (nx24010)) ;
    inv02 ix23855 (.Y (nx23856), .A (nx24012)) ;
    inv02 ix23857 (.Y (nx23858), .A (nx24012)) ;
    inv02 ix23859 (.Y (nx23860), .A (nx24012)) ;
    inv02 ix23861 (.Y (nx23862), .A (nx24012)) ;
    inv02 ix23863 (.Y (nx23864), .A (nx24012)) ;
    inv02 ix23865 (.Y (nx23866), .A (nx24012)) ;
    inv02 ix23867 (.Y (nx23868), .A (nx24012)) ;
    inv02 ix23869 (.Y (nx23870), .A (nx24014)) ;
    inv02 ix23871 (.Y (nx23872), .A (nx24014)) ;
    inv02 ix23873 (.Y (nx23874), .A (nx24014)) ;
    inv02 ix23875 (.Y (nx23876), .A (nx24014)) ;
    inv02 ix23877 (.Y (nx23878), .A (nx24014)) ;
    inv02 ix23879 (.Y (nx23880), .A (nx24014)) ;
    inv02 ix23881 (.Y (nx23882), .A (nx24014)) ;
    inv02 ix23883 (.Y (nx23884), .A (nx24016)) ;
    inv02 ix23885 (.Y (nx23886), .A (nx24016)) ;
    inv02 ix23887 (.Y (nx23888), .A (nx24016)) ;
    inv02 ix23889 (.Y (nx23890), .A (nx24016)) ;
    inv02 ix23891 (.Y (nx23892), .A (nx24016)) ;
    inv02 ix23893 (.Y (nx23894), .A (nx24016)) ;
    inv02 ix23895 (.Y (nx23896), .A (nx24016)) ;
    inv02 ix23897 (.Y (nx23898), .A (nx24018)) ;
    inv02 ix23899 (.Y (nx23900), .A (nx24018)) ;
    inv02 ix23901 (.Y (nx23902), .A (nx24018)) ;
    inv02 ix23903 (.Y (nx23904), .A (nx24018)) ;
    inv02 ix23905 (.Y (nx23906), .A (nx24018)) ;
    inv02 ix23907 (.Y (nx23908), .A (nx24018)) ;
    inv02 ix23909 (.Y (nx23910), .A (nx24018)) ;
    inv02 ix23911 (.Y (nx23912), .A (nx24020)) ;
    inv02 ix23913 (.Y (nx23914), .A (nx24020)) ;
    inv02 ix23915 (.Y (nx23916), .A (nx24020)) ;
    inv02 ix23917 (.Y (nx23918), .A (nx24020)) ;
    inv02 ix23919 (.Y (nx23920), .A (nx24020)) ;
    inv02 ix23921 (.Y (nx23922), .A (nx24020)) ;
    inv02 ix23923 (.Y (nx23924), .A (nx24020)) ;
    inv02 ix23925 (.Y (nx23926), .A (nx24022)) ;
    inv02 ix23927 (.Y (nx23928), .A (nx24022)) ;
    inv02 ix23929 (.Y (nx23930), .A (nx24022)) ;
    inv02 ix23931 (.Y (nx23932), .A (nx24022)) ;
    inv02 ix23933 (.Y (nx23934), .A (nx24022)) ;
    inv02 ix23935 (.Y (nx23936), .A (nx24022)) ;
    inv02 ix23937 (.Y (nx23938), .A (nx24022)) ;
    inv02 ix23939 (.Y (nx23940), .A (nx24024)) ;
    inv02 ix23941 (.Y (nx23942), .A (nx24024)) ;
    inv02 ix23943 (.Y (nx23944), .A (nx24024)) ;
    inv02 ix23945 (.Y (nx23946), .A (nx24024)) ;
    inv02 ix23947 (.Y (nx23948), .A (nx24024)) ;
    inv02 ix23949 (.Y (nx23950), .A (nx24024)) ;
    inv02 ix23951 (.Y (nx23952), .A (nx24024)) ;
    inv02 ix23953 (.Y (nx23954), .A (nx24026)) ;
    inv02 ix23955 (.Y (nx23956), .A (nx24026)) ;
    inv02 ix23957 (.Y (nx23958), .A (nx24026)) ;
    inv02 ix23959 (.Y (nx23960), .A (nx24026)) ;
    inv02 ix23961 (.Y (nx23962), .A (nx24026)) ;
    inv02 ix23963 (.Y (nx23964), .A (nx24026)) ;
    inv02 ix23965 (.Y (nx23966), .A (nx24026)) ;
    inv02 ix23967 (.Y (nx23968), .A (nx24028)) ;
    inv02 ix23969 (.Y (nx23970), .A (nx24028)) ;
    inv02 ix23971 (.Y (nx23972), .A (nx24028)) ;
    inv02 ix23973 (.Y (nx23974), .A (nx24028)) ;
    inv02 ix23975 (.Y (nx23976), .A (nx24028)) ;
    inv02 ix23977 (.Y (nx23978), .A (nx24028)) ;
    inv02 ix23979 (.Y (nx23980), .A (nx24028)) ;
    inv02 ix23981 (.Y (nx23982), .A (nx24030)) ;
    inv02 ix23983 (.Y (nx23984), .A (nx24030)) ;
    inv02 ix23985 (.Y (nx23986), .A (nx24030)) ;
    inv02 ix23987 (.Y (nx23988), .A (nx24030)) ;
    inv02 ix23989 (.Y (nx23990), .A (nx24030)) ;
    inv02 ix23991 (.Y (nx23992), .A (nx24030)) ;
    inv02 ix23993 (.Y (nx23994), .A (nx24030)) ;
    inv02 ix23995 (.Y (nx23996), .A (nx24032)) ;
    inv02 ix23997 (.Y (nx23998), .A (current_state[11])) ;
    inv02 ix23999 (.Y (nx24000), .A (current_state[11])) ;
    inv02 ix24001 (.Y (nx24002), .A (current_state[11])) ;
    inv02 ix24003 (.Y (nx24004), .A (current_state[11])) ;
    inv01 ix24005 (.Y (nx24006), .A (TriImgLeftEn)) ;
    inv02 ix24007 (.Y (nx24008), .A (CLK)) ;
    inv02 ix24009 (.Y (nx24010), .A (nx24038)) ;
    inv02 ix24011 (.Y (nx24012), .A (nx24038)) ;
    inv02 ix24013 (.Y (nx24014), .A (nx24038)) ;
    inv02 ix24015 (.Y (nx24016), .A (nx24038)) ;
    inv02 ix24017 (.Y (nx24018), .A (nx24038)) ;
    inv02 ix24019 (.Y (nx24020), .A (nx24038)) ;
    inv02 ix24021 (.Y (nx24022), .A (nx24038)) ;
    inv02 ix24023 (.Y (nx24024), .A (nx24040)) ;
    inv02 ix24025 (.Y (nx24026), .A (nx24040)) ;
    inv02 ix24027 (.Y (nx24028), .A (nx24040)) ;
    inv02 ix24029 (.Y (nx24030), .A (nx24040)) ;
    inv02 ix24031 (.Y (nx24032), .A (nx24040)) ;
    inv02 ix24037 (.Y (nx24038), .A (nx24008)) ;
    inv02 ix24039 (.Y (nx24040), .A (nx24008)) ;
endmodule


module triStateBuffer_6 ( D, EN, F ) ;

    input [5:0]D ;
    input EN ;
    output [5:0]F ;

    wire nx115, nx118, nx121, nx124, nx127, nx130;



    tri01 tri_F_0 (.Y (F[0]), .A (nx115), .E (EN)) ;
    inv01 ix116 (.Y (nx115), .A (D[0])) ;
    tri01 tri_F_1 (.Y (F[1]), .A (nx118), .E (EN)) ;
    inv01 ix119 (.Y (nx118), .A (D[1])) ;
    tri01 tri_F_2 (.Y (F[2]), .A (nx121), .E (EN)) ;
    inv01 ix122 (.Y (nx121), .A (D[2])) ;
    tri01 tri_F_3 (.Y (F[3]), .A (nx124), .E (EN)) ;
    inv01 ix125 (.Y (nx124), .A (D[3])) ;
    tri01 tri_F_4 (.Y (F[4]), .A (nx127), .E (EN)) ;
    inv01 ix128 (.Y (nx127), .A (D[4])) ;
    tri01 tri_F_5 (.Y (F[5]), .A (nx130), .E (EN)) ;
    inv01 ix131 (.Y (nx130), .A (D[5])) ;
endmodule


module Decoder ( \input , \output  ) ;

    input [2:0]\input  ;
    output [5:0]\output  ;

    wire nx4, nx14, nx28, nx42, nx54, nx68, nx80, nx145, nx149, nx155, nx164, 
         nx166;



    latch lat_output_0 (.Q (\output [0]), .D (nx14), .CLK (nx4)) ;
    nor03_2x ix15 (.Y (nx14), .A0 (nx164), .A1 (nx166), .A2 (\input [0])) ;
    nand02 ix5 (.Y (nx4), .A0 (nx164), .A1 (nx166)) ;
    latch lat_output_1 (.Q (\output [1]), .D (nx28), .CLK (nx4)) ;
    nor03_2x ix29 (.Y (nx28), .A0 (nx164), .A1 (nx166), .A2 (nx145)) ;
    inv01 ix146 (.Y (nx145), .A (\input [0])) ;
    latch lat_output_2 (.Q (\output [2]), .D (nx42), .CLK (nx4)) ;
    nor03_2x ix43 (.Y (nx42), .A0 (nx164), .A1 (nx149), .A2 (\input [0])) ;
    inv01 ix150 (.Y (nx149), .A (\input [1])) ;
    latch lat_output_3 (.Q (\output [3]), .D (nx54), .CLK (nx4)) ;
    nor03_2x ix55 (.Y (nx54), .A0 (nx164), .A1 (nx149), .A2 (nx145)) ;
    latch lat_output_4 (.Q (\output [4]), .D (nx68), .CLK (nx4)) ;
    nor03_2x ix69 (.Y (nx68), .A0 (nx155), .A1 (nx166), .A2 (\input [0])) ;
    inv01 ix156 (.Y (nx155), .A (\input [2])) ;
    latch lat_output_5 (.Q (\output [5]), .D (nx80), .CLK (nx4)) ;
    nor03_2x ix81 (.Y (nx80), .A0 (nx155), .A1 (nx166), .A2 (nx145)) ;
    inv02 ix163 (.Y (nx164), .A (nx155)) ;
    inv02 ix165 (.Y (nx166), .A (nx149)) ;
endmodule


module Counter_3 ( enable, reset, clk, load, \output , \input  ) ;

    input enable ;
    input reset ;
    input clk ;
    input load ;
    output [2:0]\output  ;
    input [2:0]\input  ;

    wire addResult_2, addResult_1, addResult_0, one_0, one_2, nx40, NOT_clk, nx8, 
         nx12, nx34, nx20, nx24, nx28, nx33, nx37, nx114, nx124, nx134, nx143;
    wire [6:0] \$dummy ;




    my_nadder_3 A1 (.a ({\output [2],\output [1],\output [0]}), .b ({one_2,one_2
                ,one_0}), .cin (one_2), .s ({addResult_2,addResult_1,addResult_0
                }), .cout (\$dummy [0])) ;
    fake_gnd ix94 (.Y (one_2)) ;
    fake_vcc ix92 (.Y (one_0)) ;
    dffsr_ni reg_toOutput_0__dup_1 (.Q (\output [0]), .QB (\$dummy [1]), .D (
             nx114), .CLK (clk), .S (nx8), .R (nx12)) ;
    mux21_ni ix115 (.Y (nx114), .A0 (\output [0]), .A1 (addResult_0), .S0 (
             enable)) ;
    nor02ii ix9 (.Y (nx8), .A0 (nx143), .A1 (nx40)) ;
    nor02_2x ix144 (.Y (nx143), .A0 (reset), .A1 (load)) ;
    dffr ix41 (.Q (nx40), .QB (\$dummy [2]), .D (\input [0]), .CLK (NOT_clk), .R (
         reset)) ;
    inv01 ix147 (.Y (NOT_clk), .A (clk)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (nx40), .A1 (nx143)) ;
    dffsr_ni reg_toOutput_1__dup_1 (.Q (\output [1]), .QB (\$dummy [3]), .D (
             nx124), .CLK (clk), .S (nx20), .R (nx24)) ;
    mux21_ni ix125 (.Y (nx124), .A0 (\output [1]), .A1 (addResult_1), .S0 (
             enable)) ;
    nor02ii ix21 (.Y (nx20), .A0 (nx143), .A1 (nx34)) ;
    dffr ix35 (.Q (nx34), .QB (\$dummy [4]), .D (\input [1]), .CLK (NOT_clk), .R (
         reset)) ;
    nor02_2x ix25 (.Y (nx24), .A0 (nx34), .A1 (nx143)) ;
    dffsr_ni reg_toOutput_2__dup_1 (.Q (\output [2]), .QB (\$dummy [5]), .D (
             nx134), .CLK (clk), .S (nx33), .R (nx37)) ;
    mux21_ni ix135 (.Y (nx134), .A0 (\output [2]), .A1 (addResult_2), .S0 (
             enable)) ;
    nor02ii ix34 (.Y (nx33), .A0 (nx143), .A1 (nx28)) ;
    dffr ix29 (.Q (nx28), .QB (\$dummy [6]), .D (\input [2]), .CLK (NOT_clk), .R (
         reset)) ;
    nor02_2x ix38 (.Y (nx37), .A0 (nx28), .A1 (nx143)) ;
endmodule


module my_nadder_3 ( a, b, cin, s, cout ) ;

    input [2:0]a ;
    input [2:0]b ;
    input cin ;
    output [2:0]s ;
    output cout ;

    wire temp_1, temp_0;



    my_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (s[0]), .cout (temp_0)) ;
    my_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (s[1]), .cout (
             temp_1)) ;
    my_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (s[2]), .cout (
             cout)) ;
endmodule


module my_nadder_16 ( a, b, cin, s, cout ) ;

    input [15:0]a ;
    input [15:0]b ;
    input cin ;
    output [15:0]s ;
    output cout ;

    wire temp_14, temp_13, temp_12, temp_11, temp_10, temp_9, temp_8, temp_7, 
         temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0;



    my_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (s[0]), .cout (temp_0)) ;
    my_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (s[1]), .cout (
             temp_1)) ;
    my_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (s[2]), .cout (
             temp_2)) ;
    my_adder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (s[3]), .cout (
             temp_3)) ;
    my_adder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (s[4]), .cout (
             temp_4)) ;
    my_adder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (s[5]), .cout (
             temp_5)) ;
    my_adder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (s[6]), .cout (
             temp_6)) ;
    my_adder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (s[7]), .cout (
             temp_7)) ;
    my_adder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (s[8]), .cout (
             temp_8)) ;
    my_adder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (s[9]), .cout (
             temp_9)) ;
    my_adder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (s[10]), .cout (
             temp_10)) ;
    my_adder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (s[11]), .cout (
             temp_11)) ;
    my_adder loop1_12_fx (.a (a[12]), .b (b[12]), .cin (temp_11), .s (s[12]), .cout (
             temp_12)) ;
    my_adder loop1_13_fx (.a (a[13]), .b (b[13]), .cin (temp_12), .s (s[13]), .cout (
             temp_13)) ;
    my_adder loop1_14_fx (.a (a[14]), .b (b[14]), .cin (temp_13), .s (s[14]), .cout (
             temp_14)) ;
    my_adder loop1_15_fx (.a (a[15]), .b (b[15]), .cin (temp_14), .s (s[15]), .cout (
             cout)) ;
endmodule


module ReadFilter ( current_state, LayerInfo, depthcounter, FilterCounter, 
                    Heightcounter, FILTER, FilterAddress, msbNoOfFilters, CLK, 
                    RST, QImgStat, ACKF, IndicatorFilter, DMAAddress, 
                    UpdatedAddress, outFilter0, outFilter1, donttrust, 
                    LastFilterIND, LastHeightOut, lastDepthOut ) ;

    input [14:0]current_state ;
    input [15:0]LayerInfo ;
    input [3:0]depthcounter ;
    input [3:0]FilterCounter ;
    input [4:0]Heightcounter ;
    input [399:0]FILTER ;
    input [12:0]FilterAddress ;
    input msbNoOfFilters ;
    input CLK ;
    input RST ;
    input QImgStat ;
    input ACKF ;
    output [0:0]IndicatorFilter ;
    output [12:0]DMAAddress ;
    output [12:0]UpdatedAddress ;
    output [399:0]outFilter0 ;
    output [399:0]outFilter1 ;
    output donttrust ;
    output LastFilterIND ;
    output LastHeightOut ;
    output lastDepthOut ;

    wire DFFCLK, newAddress_12, newAddress_11, newAddress_10, newAddress_9, 
         newAddress_8, newAddress_7, newAddress_6, newAddress_5, newAddress_4, 
         newAddress_3, newAddress_2, newAddress_1, newAddress_0, depthminus_3, 
         depthminus_2, depthminus_1, depthminus_0, FilterMinus_3, FilterMinus_2, 
         FilterMinus_1, FilterMinus_0, Heightminus_4, Heightminus_3, 
         Heightminus_2, Heightminus_1, Heightminus_0, filter1EN, filter2EN, 
         IndRst, tristateAddEn, secOperand_12, secOperand_3, 
         NOT_IndicatorFilter_0, nx2, nx22, nx24, nx96, nx108, nx120, nx130, 
         nx1466, nx1469, nx1471, nx1473, nx1475, nx1477, nx1479, nx1482, nx1484, 
         nx1486, nx1488, nx1491, nx1493, nx1495, nx1497;
    wire [4:0] \$dummy ;




    assign LastHeightOut = donttrust ;
    my_nadder_4 adder2 (.a ({LayerInfo[12],LayerInfo[11],LayerInfo[10],
                LayerInfo[9]}), .b ({secOperand_3,secOperand_3,secOperand_3,
                secOperand_3}), .cin (secOperand_12), .s ({depthminus_3,
                depthminus_2,depthminus_1,depthminus_0}), .cout (\$dummy [0])) ;
    my_nadder_5 adder3 (.a ({LayerInfo[8],LayerInfo[7],LayerInfo[6],LayerInfo[5]
                ,LayerInfo[4]}), .b ({secOperand_3,secOperand_3,secOperand_3,
                secOperand_3,secOperand_3}), .cin (secOperand_12), .s ({
                Heightminus_4,Heightminus_3,Heightminus_2,Heightminus_1,
                Heightminus_0}), .cout (\$dummy [1])) ;
    my_nadder_4 adder4 (.a ({LayerInfo[3],LayerInfo[2],LayerInfo[1],LayerInfo[0]
                }), .b ({secOperand_3,secOperand_3,secOperand_3,secOperand_3}), 
                .cin (secOperand_12), .s ({FilterMinus_3,FilterMinus_2,
                FilterMinus_1,FilterMinus_0}), .cout (\$dummy [2])) ;
    nBitRegister_400 F0 (.D ({FILTER[399],FILTER[398],FILTER[397],FILTER[396],
                     FILTER[395],FILTER[394],FILTER[393],FILTER[392],FILTER[391]
                     ,FILTER[390],FILTER[389],FILTER[388],FILTER[387],
                     FILTER[386],FILTER[385],FILTER[384],FILTER[383],FILTER[382]
                     ,FILTER[381],FILTER[380],FILTER[379],FILTER[378],
                     FILTER[377],FILTER[376],FILTER[375],FILTER[374],FILTER[373]
                     ,FILTER[372],FILTER[371],FILTER[370],FILTER[369],
                     FILTER[368],FILTER[367],FILTER[366],FILTER[365],FILTER[364]
                     ,FILTER[363],FILTER[362],FILTER[361],FILTER[360],
                     FILTER[359],FILTER[358],FILTER[357],FILTER[356],FILTER[355]
                     ,FILTER[354],FILTER[353],FILTER[352],FILTER[351],
                     FILTER[350],FILTER[349],FILTER[348],FILTER[347],FILTER[346]
                     ,FILTER[345],FILTER[344],FILTER[343],FILTER[342],
                     FILTER[341],FILTER[340],FILTER[339],FILTER[338],FILTER[337]
                     ,FILTER[336],FILTER[335],FILTER[334],FILTER[333],
                     FILTER[332],FILTER[331],FILTER[330],FILTER[329],FILTER[328]
                     ,FILTER[327],FILTER[326],FILTER[325],FILTER[324],
                     FILTER[323],FILTER[322],FILTER[321],FILTER[320],FILTER[319]
                     ,FILTER[318],FILTER[317],FILTER[316],FILTER[315],
                     FILTER[314],FILTER[313],FILTER[312],FILTER[311],FILTER[310]
                     ,FILTER[309],FILTER[308],FILTER[307],FILTER[306],
                     FILTER[305],FILTER[304],FILTER[303],FILTER[302],FILTER[301]
                     ,FILTER[300],FILTER[299],FILTER[298],FILTER[297],
                     FILTER[296],FILTER[295],FILTER[294],FILTER[293],FILTER[292]
                     ,FILTER[291],FILTER[290],FILTER[289],FILTER[288],
                     FILTER[287],FILTER[286],FILTER[285],FILTER[284],FILTER[283]
                     ,FILTER[282],FILTER[281],FILTER[280],FILTER[279],
                     FILTER[278],FILTER[277],FILTER[276],FILTER[275],FILTER[274]
                     ,FILTER[273],FILTER[272],FILTER[271],FILTER[270],
                     FILTER[269],FILTER[268],FILTER[267],FILTER[266],FILTER[265]
                     ,FILTER[264],FILTER[263],FILTER[262],FILTER[261],
                     FILTER[260],FILTER[259],FILTER[258],FILTER[257],FILTER[256]
                     ,FILTER[255],FILTER[254],FILTER[253],FILTER[252],
                     FILTER[251],FILTER[250],FILTER[249],FILTER[248],FILTER[247]
                     ,FILTER[246],FILTER[245],FILTER[244],FILTER[243],
                     FILTER[242],FILTER[241],FILTER[240],FILTER[239],FILTER[238]
                     ,FILTER[237],FILTER[236],FILTER[235],FILTER[234],
                     FILTER[233],FILTER[232],FILTER[231],FILTER[230],FILTER[229]
                     ,FILTER[228],FILTER[227],FILTER[226],FILTER[225],
                     FILTER[224],FILTER[223],FILTER[222],FILTER[221],FILTER[220]
                     ,FILTER[219],FILTER[218],FILTER[217],FILTER[216],
                     FILTER[215],FILTER[214],FILTER[213],FILTER[212],FILTER[211]
                     ,FILTER[210],FILTER[209],FILTER[208],FILTER[207],
                     FILTER[206],FILTER[205],FILTER[204],FILTER[203],FILTER[202]
                     ,FILTER[201],FILTER[200],FILTER[199],FILTER[198],
                     FILTER[197],FILTER[196],FILTER[195],FILTER[194],FILTER[193]
                     ,FILTER[192],FILTER[191],FILTER[190],FILTER[189],
                     FILTER[188],FILTER[187],FILTER[186],FILTER[185],FILTER[184]
                     ,FILTER[183],FILTER[182],FILTER[181],FILTER[180],
                     FILTER[179],FILTER[178],FILTER[177],FILTER[176],FILTER[175]
                     ,FILTER[174],FILTER[173],FILTER[172],FILTER[171],
                     FILTER[170],FILTER[169],FILTER[168],FILTER[167],FILTER[166]
                     ,FILTER[165],FILTER[164],FILTER[163],FILTER[162],
                     FILTER[161],FILTER[160],FILTER[159],FILTER[158],FILTER[157]
                     ,FILTER[156],FILTER[155],FILTER[154],FILTER[153],
                     FILTER[152],FILTER[151],FILTER[150],FILTER[149],FILTER[148]
                     ,FILTER[147],FILTER[146],FILTER[145],FILTER[144],
                     FILTER[143],FILTER[142],FILTER[141],FILTER[140],FILTER[139]
                     ,FILTER[138],FILTER[137],FILTER[136],FILTER[135],
                     FILTER[134],FILTER[133],FILTER[132],FILTER[131],FILTER[130]
                     ,FILTER[129],FILTER[128],FILTER[127],FILTER[126],
                     FILTER[125],FILTER[124],FILTER[123],FILTER[122],FILTER[121]
                     ,FILTER[120],FILTER[119],FILTER[118],FILTER[117],
                     FILTER[116],FILTER[115],FILTER[114],FILTER[113],FILTER[112]
                     ,FILTER[111],FILTER[110],FILTER[109],FILTER[108],
                     FILTER[107],FILTER[106],FILTER[105],FILTER[104],FILTER[103]
                     ,FILTER[102],FILTER[101],FILTER[100],FILTER[99],FILTER[98],
                     FILTER[97],FILTER[96],FILTER[95],FILTER[94],FILTER[93],
                     FILTER[92],FILTER[91],FILTER[90],FILTER[89],FILTER[88],
                     FILTER[87],FILTER[86],FILTER[85],FILTER[84],FILTER[83],
                     FILTER[82],FILTER[81],FILTER[80],FILTER[79],FILTER[78],
                     FILTER[77],FILTER[76],FILTER[75],FILTER[74],FILTER[73],
                     FILTER[72],FILTER[71],FILTER[70],FILTER[69],FILTER[68],
                     FILTER[67],FILTER[66],FILTER[65],FILTER[64],FILTER[63],
                     FILTER[62],FILTER[61],FILTER[60],FILTER[59],FILTER[58],
                     FILTER[57],FILTER[56],FILTER[55],FILTER[54],FILTER[53],
                     FILTER[52],FILTER[51],FILTER[50],FILTER[49],FILTER[48],
                     FILTER[47],FILTER[46],FILTER[45],FILTER[44],FILTER[43],
                     FILTER[42],FILTER[41],FILTER[40],FILTER[39],FILTER[38],
                     FILTER[37],FILTER[36],FILTER[35],FILTER[34],FILTER[33],
                     FILTER[32],FILTER[31],FILTER[30],FILTER[29],FILTER[28],
                     FILTER[27],FILTER[26],FILTER[25],FILTER[24],FILTER[23],
                     FILTER[22],FILTER[21],FILTER[20],FILTER[19],FILTER[18],
                     FILTER[17],FILTER[16],FILTER[15],FILTER[14],FILTER[13],
                     FILTER[12],FILTER[11],FILTER[10],FILTER[9],FILTER[8],
                     FILTER[7],FILTER[6],FILTER[5],FILTER[4],FILTER[3],FILTER[2]
                     ,FILTER[1],FILTER[0]}), .CLK (CLK), .RST (RST), .EN (
                     filter1EN), .Q ({outFilter0[399],outFilter0[398],
                     outFilter0[397],outFilter0[396],outFilter0[395],
                     outFilter0[394],outFilter0[393],outFilter0[392],
                     outFilter0[391],outFilter0[390],outFilter0[389],
                     outFilter0[388],outFilter0[387],outFilter0[386],
                     outFilter0[385],outFilter0[384],outFilter0[383],
                     outFilter0[382],outFilter0[381],outFilter0[380],
                     outFilter0[379],outFilter0[378],outFilter0[377],
                     outFilter0[376],outFilter0[375],outFilter0[374],
                     outFilter0[373],outFilter0[372],outFilter0[371],
                     outFilter0[370],outFilter0[369],outFilter0[368],
                     outFilter0[367],outFilter0[366],outFilter0[365],
                     outFilter0[364],outFilter0[363],outFilter0[362],
                     outFilter0[361],outFilter0[360],outFilter0[359],
                     outFilter0[358],outFilter0[357],outFilter0[356],
                     outFilter0[355],outFilter0[354],outFilter0[353],
                     outFilter0[352],outFilter0[351],outFilter0[350],
                     outFilter0[349],outFilter0[348],outFilter0[347],
                     outFilter0[346],outFilter0[345],outFilter0[344],
                     outFilter0[343],outFilter0[342],outFilter0[341],
                     outFilter0[340],outFilter0[339],outFilter0[338],
                     outFilter0[337],outFilter0[336],outFilter0[335],
                     outFilter0[334],outFilter0[333],outFilter0[332],
                     outFilter0[331],outFilter0[330],outFilter0[329],
                     outFilter0[328],outFilter0[327],outFilter0[326],
                     outFilter0[325],outFilter0[324],outFilter0[323],
                     outFilter0[322],outFilter0[321],outFilter0[320],
                     outFilter0[319],outFilter0[318],outFilter0[317],
                     outFilter0[316],outFilter0[315],outFilter0[314],
                     outFilter0[313],outFilter0[312],outFilter0[311],
                     outFilter0[310],outFilter0[309],outFilter0[308],
                     outFilter0[307],outFilter0[306],outFilter0[305],
                     outFilter0[304],outFilter0[303],outFilter0[302],
                     outFilter0[301],outFilter0[300],outFilter0[299],
                     outFilter0[298],outFilter0[297],outFilter0[296],
                     outFilter0[295],outFilter0[294],outFilter0[293],
                     outFilter0[292],outFilter0[291],outFilter0[290],
                     outFilter0[289],outFilter0[288],outFilter0[287],
                     outFilter0[286],outFilter0[285],outFilter0[284],
                     outFilter0[283],outFilter0[282],outFilter0[281],
                     outFilter0[280],outFilter0[279],outFilter0[278],
                     outFilter0[277],outFilter0[276],outFilter0[275],
                     outFilter0[274],outFilter0[273],outFilter0[272],
                     outFilter0[271],outFilter0[270],outFilter0[269],
                     outFilter0[268],outFilter0[267],outFilter0[266],
                     outFilter0[265],outFilter0[264],outFilter0[263],
                     outFilter0[262],outFilter0[261],outFilter0[260],
                     outFilter0[259],outFilter0[258],outFilter0[257],
                     outFilter0[256],outFilter0[255],outFilter0[254],
                     outFilter0[253],outFilter0[252],outFilter0[251],
                     outFilter0[250],outFilter0[249],outFilter0[248],
                     outFilter0[247],outFilter0[246],outFilter0[245],
                     outFilter0[244],outFilter0[243],outFilter0[242],
                     outFilter0[241],outFilter0[240],outFilter0[239],
                     outFilter0[238],outFilter0[237],outFilter0[236],
                     outFilter0[235],outFilter0[234],outFilter0[233],
                     outFilter0[232],outFilter0[231],outFilter0[230],
                     outFilter0[229],outFilter0[228],outFilter0[227],
                     outFilter0[226],outFilter0[225],outFilter0[224],
                     outFilter0[223],outFilter0[222],outFilter0[221],
                     outFilter0[220],outFilter0[219],outFilter0[218],
                     outFilter0[217],outFilter0[216],outFilter0[215],
                     outFilter0[214],outFilter0[213],outFilter0[212],
                     outFilter0[211],outFilter0[210],outFilter0[209],
                     outFilter0[208],outFilter0[207],outFilter0[206],
                     outFilter0[205],outFilter0[204],outFilter0[203],
                     outFilter0[202],outFilter0[201],outFilter0[200],
                     outFilter0[199],outFilter0[198],outFilter0[197],
                     outFilter0[196],outFilter0[195],outFilter0[194],
                     outFilter0[193],outFilter0[192],outFilter0[191],
                     outFilter0[190],outFilter0[189],outFilter0[188],
                     outFilter0[187],outFilter0[186],outFilter0[185],
                     outFilter0[184],outFilter0[183],outFilter0[182],
                     outFilter0[181],outFilter0[180],outFilter0[179],
                     outFilter0[178],outFilter0[177],outFilter0[176],
                     outFilter0[175],outFilter0[174],outFilter0[173],
                     outFilter0[172],outFilter0[171],outFilter0[170],
                     outFilter0[169],outFilter0[168],outFilter0[167],
                     outFilter0[166],outFilter0[165],outFilter0[164],
                     outFilter0[163],outFilter0[162],outFilter0[161],
                     outFilter0[160],outFilter0[159],outFilter0[158],
                     outFilter0[157],outFilter0[156],outFilter0[155],
                     outFilter0[154],outFilter0[153],outFilter0[152],
                     outFilter0[151],outFilter0[150],outFilter0[149],
                     outFilter0[148],outFilter0[147],outFilter0[146],
                     outFilter0[145],outFilter0[144],outFilter0[143],
                     outFilter0[142],outFilter0[141],outFilter0[140],
                     outFilter0[139],outFilter0[138],outFilter0[137],
                     outFilter0[136],outFilter0[135],outFilter0[134],
                     outFilter0[133],outFilter0[132],outFilter0[131],
                     outFilter0[130],outFilter0[129],outFilter0[128],
                     outFilter0[127],outFilter0[126],outFilter0[125],
                     outFilter0[124],outFilter0[123],outFilter0[122],
                     outFilter0[121],outFilter0[120],outFilter0[119],
                     outFilter0[118],outFilter0[117],outFilter0[116],
                     outFilter0[115],outFilter0[114],outFilter0[113],
                     outFilter0[112],outFilter0[111],outFilter0[110],
                     outFilter0[109],outFilter0[108],outFilter0[107],
                     outFilter0[106],outFilter0[105],outFilter0[104],
                     outFilter0[103],outFilter0[102],outFilter0[101],
                     outFilter0[100],outFilter0[99],outFilter0[98],
                     outFilter0[97],outFilter0[96],outFilter0[95],outFilter0[94]
                     ,outFilter0[93],outFilter0[92],outFilter0[91],
                     outFilter0[90],outFilter0[89],outFilter0[88],outFilter0[87]
                     ,outFilter0[86],outFilter0[85],outFilter0[84],
                     outFilter0[83],outFilter0[82],outFilter0[81],outFilter0[80]
                     ,outFilter0[79],outFilter0[78],outFilter0[77],
                     outFilter0[76],outFilter0[75],outFilter0[74],outFilter0[73]
                     ,outFilter0[72],outFilter0[71],outFilter0[70],
                     outFilter0[69],outFilter0[68],outFilter0[67],outFilter0[66]
                     ,outFilter0[65],outFilter0[64],outFilter0[63],
                     outFilter0[62],outFilter0[61],outFilter0[60],outFilter0[59]
                     ,outFilter0[58],outFilter0[57],outFilter0[56],
                     outFilter0[55],outFilter0[54],outFilter0[53],outFilter0[52]
                     ,outFilter0[51],outFilter0[50],outFilter0[49],
                     outFilter0[48],outFilter0[47],outFilter0[46],outFilter0[45]
                     ,outFilter0[44],outFilter0[43],outFilter0[42],
                     outFilter0[41],outFilter0[40],outFilter0[39],outFilter0[38]
                     ,outFilter0[37],outFilter0[36],outFilter0[35],
                     outFilter0[34],outFilter0[33],outFilter0[32],outFilter0[31]
                     ,outFilter0[30],outFilter0[29],outFilter0[28],
                     outFilter0[27],outFilter0[26],outFilter0[25],outFilter0[24]
                     ,outFilter0[23],outFilter0[22],outFilter0[21],
                     outFilter0[20],outFilter0[19],outFilter0[18],outFilter0[17]
                     ,outFilter0[16],outFilter0[15],outFilter0[14],
                     outFilter0[13],outFilter0[12],outFilter0[11],outFilter0[10]
                     ,outFilter0[9],outFilter0[8],outFilter0[7],outFilter0[6],
                     outFilter0[5],outFilter0[4],outFilter0[3],outFilter0[2],
                     outFilter0[1],outFilter0[0]})) ;
    nBitRegister_400 F1 (.D ({FILTER[399],FILTER[398],FILTER[397],FILTER[396],
                     FILTER[395],FILTER[394],FILTER[393],FILTER[392],FILTER[391]
                     ,FILTER[390],FILTER[389],FILTER[388],FILTER[387],
                     FILTER[386],FILTER[385],FILTER[384],FILTER[383],FILTER[382]
                     ,FILTER[381],FILTER[380],FILTER[379],FILTER[378],
                     FILTER[377],FILTER[376],FILTER[375],FILTER[374],FILTER[373]
                     ,FILTER[372],FILTER[371],FILTER[370],FILTER[369],
                     FILTER[368],FILTER[367],FILTER[366],FILTER[365],FILTER[364]
                     ,FILTER[363],FILTER[362],FILTER[361],FILTER[360],
                     FILTER[359],FILTER[358],FILTER[357],FILTER[356],FILTER[355]
                     ,FILTER[354],FILTER[353],FILTER[352],FILTER[351],
                     FILTER[350],FILTER[349],FILTER[348],FILTER[347],FILTER[346]
                     ,FILTER[345],FILTER[344],FILTER[343],FILTER[342],
                     FILTER[341],FILTER[340],FILTER[339],FILTER[338],FILTER[337]
                     ,FILTER[336],FILTER[335],FILTER[334],FILTER[333],
                     FILTER[332],FILTER[331],FILTER[330],FILTER[329],FILTER[328]
                     ,FILTER[327],FILTER[326],FILTER[325],FILTER[324],
                     FILTER[323],FILTER[322],FILTER[321],FILTER[320],FILTER[319]
                     ,FILTER[318],FILTER[317],FILTER[316],FILTER[315],
                     FILTER[314],FILTER[313],FILTER[312],FILTER[311],FILTER[310]
                     ,FILTER[309],FILTER[308],FILTER[307],FILTER[306],
                     FILTER[305],FILTER[304],FILTER[303],FILTER[302],FILTER[301]
                     ,FILTER[300],FILTER[299],FILTER[298],FILTER[297],
                     FILTER[296],FILTER[295],FILTER[294],FILTER[293],FILTER[292]
                     ,FILTER[291],FILTER[290],FILTER[289],FILTER[288],
                     FILTER[287],FILTER[286],FILTER[285],FILTER[284],FILTER[283]
                     ,FILTER[282],FILTER[281],FILTER[280],FILTER[279],
                     FILTER[278],FILTER[277],FILTER[276],FILTER[275],FILTER[274]
                     ,FILTER[273],FILTER[272],FILTER[271],FILTER[270],
                     FILTER[269],FILTER[268],FILTER[267],FILTER[266],FILTER[265]
                     ,FILTER[264],FILTER[263],FILTER[262],FILTER[261],
                     FILTER[260],FILTER[259],FILTER[258],FILTER[257],FILTER[256]
                     ,FILTER[255],FILTER[254],FILTER[253],FILTER[252],
                     FILTER[251],FILTER[250],FILTER[249],FILTER[248],FILTER[247]
                     ,FILTER[246],FILTER[245],FILTER[244],FILTER[243],
                     FILTER[242],FILTER[241],FILTER[240],FILTER[239],FILTER[238]
                     ,FILTER[237],FILTER[236],FILTER[235],FILTER[234],
                     FILTER[233],FILTER[232],FILTER[231],FILTER[230],FILTER[229]
                     ,FILTER[228],FILTER[227],FILTER[226],FILTER[225],
                     FILTER[224],FILTER[223],FILTER[222],FILTER[221],FILTER[220]
                     ,FILTER[219],FILTER[218],FILTER[217],FILTER[216],
                     FILTER[215],FILTER[214],FILTER[213],FILTER[212],FILTER[211]
                     ,FILTER[210],FILTER[209],FILTER[208],FILTER[207],
                     FILTER[206],FILTER[205],FILTER[204],FILTER[203],FILTER[202]
                     ,FILTER[201],FILTER[200],FILTER[199],FILTER[198],
                     FILTER[197],FILTER[196],FILTER[195],FILTER[194],FILTER[193]
                     ,FILTER[192],FILTER[191],FILTER[190],FILTER[189],
                     FILTER[188],FILTER[187],FILTER[186],FILTER[185],FILTER[184]
                     ,FILTER[183],FILTER[182],FILTER[181],FILTER[180],
                     FILTER[179],FILTER[178],FILTER[177],FILTER[176],FILTER[175]
                     ,FILTER[174],FILTER[173],FILTER[172],FILTER[171],
                     FILTER[170],FILTER[169],FILTER[168],FILTER[167],FILTER[166]
                     ,FILTER[165],FILTER[164],FILTER[163],FILTER[162],
                     FILTER[161],FILTER[160],FILTER[159],FILTER[158],FILTER[157]
                     ,FILTER[156],FILTER[155],FILTER[154],FILTER[153],
                     FILTER[152],FILTER[151],FILTER[150],FILTER[149],FILTER[148]
                     ,FILTER[147],FILTER[146],FILTER[145],FILTER[144],
                     FILTER[143],FILTER[142],FILTER[141],FILTER[140],FILTER[139]
                     ,FILTER[138],FILTER[137],FILTER[136],FILTER[135],
                     FILTER[134],FILTER[133],FILTER[132],FILTER[131],FILTER[130]
                     ,FILTER[129],FILTER[128],FILTER[127],FILTER[126],
                     FILTER[125],FILTER[124],FILTER[123],FILTER[122],FILTER[121]
                     ,FILTER[120],FILTER[119],FILTER[118],FILTER[117],
                     FILTER[116],FILTER[115],FILTER[114],FILTER[113],FILTER[112]
                     ,FILTER[111],FILTER[110],FILTER[109],FILTER[108],
                     FILTER[107],FILTER[106],FILTER[105],FILTER[104],FILTER[103]
                     ,FILTER[102],FILTER[101],FILTER[100],FILTER[99],FILTER[98],
                     FILTER[97],FILTER[96],FILTER[95],FILTER[94],FILTER[93],
                     FILTER[92],FILTER[91],FILTER[90],FILTER[89],FILTER[88],
                     FILTER[87],FILTER[86],FILTER[85],FILTER[84],FILTER[83],
                     FILTER[82],FILTER[81],FILTER[80],FILTER[79],FILTER[78],
                     FILTER[77],FILTER[76],FILTER[75],FILTER[74],FILTER[73],
                     FILTER[72],FILTER[71],FILTER[70],FILTER[69],FILTER[68],
                     FILTER[67],FILTER[66],FILTER[65],FILTER[64],FILTER[63],
                     FILTER[62],FILTER[61],FILTER[60],FILTER[59],FILTER[58],
                     FILTER[57],FILTER[56],FILTER[55],FILTER[54],FILTER[53],
                     FILTER[52],FILTER[51],FILTER[50],FILTER[49],FILTER[48],
                     FILTER[47],FILTER[46],FILTER[45],FILTER[44],FILTER[43],
                     FILTER[42],FILTER[41],FILTER[40],FILTER[39],FILTER[38],
                     FILTER[37],FILTER[36],FILTER[35],FILTER[34],FILTER[33],
                     FILTER[32],FILTER[31],FILTER[30],FILTER[29],FILTER[28],
                     FILTER[27],FILTER[26],FILTER[25],FILTER[24],FILTER[23],
                     FILTER[22],FILTER[21],FILTER[20],FILTER[19],FILTER[18],
                     FILTER[17],FILTER[16],FILTER[15],FILTER[14],FILTER[13],
                     FILTER[12],FILTER[11],FILTER[10],FILTER[9],FILTER[8],
                     FILTER[7],FILTER[6],FILTER[5],FILTER[4],FILTER[3],FILTER[2]
                     ,FILTER[1],FILTER[0]}), .CLK (CLK), .RST (RST), .EN (
                     filter2EN), .Q ({outFilter1[399],outFilter1[398],
                     outFilter1[397],outFilter1[396],outFilter1[395],
                     outFilter1[394],outFilter1[393],outFilter1[392],
                     outFilter1[391],outFilter1[390],outFilter1[389],
                     outFilter1[388],outFilter1[387],outFilter1[386],
                     outFilter1[385],outFilter1[384],outFilter1[383],
                     outFilter1[382],outFilter1[381],outFilter1[380],
                     outFilter1[379],outFilter1[378],outFilter1[377],
                     outFilter1[376],outFilter1[375],outFilter1[374],
                     outFilter1[373],outFilter1[372],outFilter1[371],
                     outFilter1[370],outFilter1[369],outFilter1[368],
                     outFilter1[367],outFilter1[366],outFilter1[365],
                     outFilter1[364],outFilter1[363],outFilter1[362],
                     outFilter1[361],outFilter1[360],outFilter1[359],
                     outFilter1[358],outFilter1[357],outFilter1[356],
                     outFilter1[355],outFilter1[354],outFilter1[353],
                     outFilter1[352],outFilter1[351],outFilter1[350],
                     outFilter1[349],outFilter1[348],outFilter1[347],
                     outFilter1[346],outFilter1[345],outFilter1[344],
                     outFilter1[343],outFilter1[342],outFilter1[341],
                     outFilter1[340],outFilter1[339],outFilter1[338],
                     outFilter1[337],outFilter1[336],outFilter1[335],
                     outFilter1[334],outFilter1[333],outFilter1[332],
                     outFilter1[331],outFilter1[330],outFilter1[329],
                     outFilter1[328],outFilter1[327],outFilter1[326],
                     outFilter1[325],outFilter1[324],outFilter1[323],
                     outFilter1[322],outFilter1[321],outFilter1[320],
                     outFilter1[319],outFilter1[318],outFilter1[317],
                     outFilter1[316],outFilter1[315],outFilter1[314],
                     outFilter1[313],outFilter1[312],outFilter1[311],
                     outFilter1[310],outFilter1[309],outFilter1[308],
                     outFilter1[307],outFilter1[306],outFilter1[305],
                     outFilter1[304],outFilter1[303],outFilter1[302],
                     outFilter1[301],outFilter1[300],outFilter1[299],
                     outFilter1[298],outFilter1[297],outFilter1[296],
                     outFilter1[295],outFilter1[294],outFilter1[293],
                     outFilter1[292],outFilter1[291],outFilter1[290],
                     outFilter1[289],outFilter1[288],outFilter1[287],
                     outFilter1[286],outFilter1[285],outFilter1[284],
                     outFilter1[283],outFilter1[282],outFilter1[281],
                     outFilter1[280],outFilter1[279],outFilter1[278],
                     outFilter1[277],outFilter1[276],outFilter1[275],
                     outFilter1[274],outFilter1[273],outFilter1[272],
                     outFilter1[271],outFilter1[270],outFilter1[269],
                     outFilter1[268],outFilter1[267],outFilter1[266],
                     outFilter1[265],outFilter1[264],outFilter1[263],
                     outFilter1[262],outFilter1[261],outFilter1[260],
                     outFilter1[259],outFilter1[258],outFilter1[257],
                     outFilter1[256],outFilter1[255],outFilter1[254],
                     outFilter1[253],outFilter1[252],outFilter1[251],
                     outFilter1[250],outFilter1[249],outFilter1[248],
                     outFilter1[247],outFilter1[246],outFilter1[245],
                     outFilter1[244],outFilter1[243],outFilter1[242],
                     outFilter1[241],outFilter1[240],outFilter1[239],
                     outFilter1[238],outFilter1[237],outFilter1[236],
                     outFilter1[235],outFilter1[234],outFilter1[233],
                     outFilter1[232],outFilter1[231],outFilter1[230],
                     outFilter1[229],outFilter1[228],outFilter1[227],
                     outFilter1[226],outFilter1[225],outFilter1[224],
                     outFilter1[223],outFilter1[222],outFilter1[221],
                     outFilter1[220],outFilter1[219],outFilter1[218],
                     outFilter1[217],outFilter1[216],outFilter1[215],
                     outFilter1[214],outFilter1[213],outFilter1[212],
                     outFilter1[211],outFilter1[210],outFilter1[209],
                     outFilter1[208],outFilter1[207],outFilter1[206],
                     outFilter1[205],outFilter1[204],outFilter1[203],
                     outFilter1[202],outFilter1[201],outFilter1[200],
                     outFilter1[199],outFilter1[198],outFilter1[197],
                     outFilter1[196],outFilter1[195],outFilter1[194],
                     outFilter1[193],outFilter1[192],outFilter1[191],
                     outFilter1[190],outFilter1[189],outFilter1[188],
                     outFilter1[187],outFilter1[186],outFilter1[185],
                     outFilter1[184],outFilter1[183],outFilter1[182],
                     outFilter1[181],outFilter1[180],outFilter1[179],
                     outFilter1[178],outFilter1[177],outFilter1[176],
                     outFilter1[175],outFilter1[174],outFilter1[173],
                     outFilter1[172],outFilter1[171],outFilter1[170],
                     outFilter1[169],outFilter1[168],outFilter1[167],
                     outFilter1[166],outFilter1[165],outFilter1[164],
                     outFilter1[163],outFilter1[162],outFilter1[161],
                     outFilter1[160],outFilter1[159],outFilter1[158],
                     outFilter1[157],outFilter1[156],outFilter1[155],
                     outFilter1[154],outFilter1[153],outFilter1[152],
                     outFilter1[151],outFilter1[150],outFilter1[149],
                     outFilter1[148],outFilter1[147],outFilter1[146],
                     outFilter1[145],outFilter1[144],outFilter1[143],
                     outFilter1[142],outFilter1[141],outFilter1[140],
                     outFilter1[139],outFilter1[138],outFilter1[137],
                     outFilter1[136],outFilter1[135],outFilter1[134],
                     outFilter1[133],outFilter1[132],outFilter1[131],
                     outFilter1[130],outFilter1[129],outFilter1[128],
                     outFilter1[127],outFilter1[126],outFilter1[125],
                     outFilter1[124],outFilter1[123],outFilter1[122],
                     outFilter1[121],outFilter1[120],outFilter1[119],
                     outFilter1[118],outFilter1[117],outFilter1[116],
                     outFilter1[115],outFilter1[114],outFilter1[113],
                     outFilter1[112],outFilter1[111],outFilter1[110],
                     outFilter1[109],outFilter1[108],outFilter1[107],
                     outFilter1[106],outFilter1[105],outFilter1[104],
                     outFilter1[103],outFilter1[102],outFilter1[101],
                     outFilter1[100],outFilter1[99],outFilter1[98],
                     outFilter1[97],outFilter1[96],outFilter1[95],outFilter1[94]
                     ,outFilter1[93],outFilter1[92],outFilter1[91],
                     outFilter1[90],outFilter1[89],outFilter1[88],outFilter1[87]
                     ,outFilter1[86],outFilter1[85],outFilter1[84],
                     outFilter1[83],outFilter1[82],outFilter1[81],outFilter1[80]
                     ,outFilter1[79],outFilter1[78],outFilter1[77],
                     outFilter1[76],outFilter1[75],outFilter1[74],outFilter1[73]
                     ,outFilter1[72],outFilter1[71],outFilter1[70],
                     outFilter1[69],outFilter1[68],outFilter1[67],outFilter1[66]
                     ,outFilter1[65],outFilter1[64],outFilter1[63],
                     outFilter1[62],outFilter1[61],outFilter1[60],outFilter1[59]
                     ,outFilter1[58],outFilter1[57],outFilter1[56],
                     outFilter1[55],outFilter1[54],outFilter1[53],outFilter1[52]
                     ,outFilter1[51],outFilter1[50],outFilter1[49],
                     outFilter1[48],outFilter1[47],outFilter1[46],outFilter1[45]
                     ,outFilter1[44],outFilter1[43],outFilter1[42],
                     outFilter1[41],outFilter1[40],outFilter1[39],outFilter1[38]
                     ,outFilter1[37],outFilter1[36],outFilter1[35],
                     outFilter1[34],outFilter1[33],outFilter1[32],outFilter1[31]
                     ,outFilter1[30],outFilter1[29],outFilter1[28],
                     outFilter1[27],outFilter1[26],outFilter1[25],outFilter1[24]
                     ,outFilter1[23],outFilter1[22],outFilter1[21],
                     outFilter1[20],outFilter1[19],outFilter1[18],outFilter1[17]
                     ,outFilter1[16],outFilter1[15],outFilter1[14],
                     outFilter1[13],outFilter1[12],outFilter1[11],outFilter1[10]
                     ,outFilter1[9],outFilter1[8],outFilter1[7],outFilter1[6],
                     outFilter1[5],outFilter1[4],outFilter1[3],outFilter1[2],
                     outFilter1[1],outFilter1[0]})) ;
    nBitRegister_1 DDF0 (.D ({NOT_IndicatorFilter_0}), .CLK (DFFCLK), .RST (
                   IndRst), .EN (secOperand_3), .Q ({IndicatorFilter[0]})) ;
    triStateBuffer_13 tsb0 (.D ({FilterAddress[12],FilterAddress[11],
                      FilterAddress[10],FilterAddress[9],FilterAddress[8],
                      FilterAddress[7],FilterAddress[6],FilterAddress[5],
                      FilterAddress[4],FilterAddress[3],FilterAddress[2],
                      FilterAddress[1],FilterAddress[0]}), .EN (tristateAddEn), 
                      .F ({DMAAddress[12],DMAAddress[11],DMAAddress[10],
                      DMAAddress[9],DMAAddress[8],DMAAddress[7],DMAAddress[6],
                      DMAAddress[5],DMAAddress[4],DMAAddress[3],DMAAddress[2],
                      DMAAddress[1],DMAAddress[0]})) ;
    my_nadder_13 adder0 (.a ({FilterAddress[12],FilterAddress[11],
                 FilterAddress[10],FilterAddress[9],FilterAddress[8],
                 FilterAddress[7],FilterAddress[6],FilterAddress[5],
                 FilterAddress[4],FilterAddress[3],FilterAddress[2],
                 FilterAddress[1],FilterAddress[0]}), .b ({secOperand_12,
                 secOperand_12,secOperand_12,secOperand_12,secOperand_12,
                 secOperand_12,secOperand_12,secOperand_12,msbNoOfFilters,
                 secOperand_3,secOperand_12,secOperand_12,secOperand_3}), .cin (
                 secOperand_12), .s ({newAddress_12,newAddress_11,newAddress_10,
                 newAddress_9,newAddress_8,newAddress_7,newAddress_6,
                 newAddress_5,newAddress_4,newAddress_3,newAddress_2,
                 newAddress_1,newAddress_0}), .cout (\$dummy [3])) ;
    triStateBuffer_13 tsb2 (.D ({newAddress_12,newAddress_11,newAddress_10,
                      newAddress_9,newAddress_8,newAddress_7,newAddress_6,
                      newAddress_5,newAddress_4,newAddress_3,newAddress_2,
                      newAddress_1,newAddress_0}), .EN (tristateAddEn), .F ({
                      UpdatedAddress[12],UpdatedAddress[11],UpdatedAddress[10],
                      UpdatedAddress[9],UpdatedAddress[8],UpdatedAddress[7],
                      UpdatedAddress[6],UpdatedAddress[5],UpdatedAddress[4],
                      UpdatedAddress[3],UpdatedAddress[2],UpdatedAddress[1],
                      UpdatedAddress[0]})) ;
    inv01 ix1459 (.Y (NOT_IndicatorFilter_0), .A (IndicatorFilter[0])) ;
    fake_vcc ix1418 (.Y (secOperand_3)) ;
    fake_gnd ix1416 (.Y (secOperand_12)) ;
    or02 ix5 (.Y (tristateAddEn), .A0 (nx2), .A1 (current_state[5])) ;
    nor02ii ix3 (.Y (nx2), .A0 (IndicatorFilter[0]), .A1 (current_state[7])) ;
    ao21 ix101 (.Y (IndRst), .A0 (current_state[10]), .A1 (nx96), .B0 (RST)) ;
    nand03 ix97 (.Y (nx96), .A0 (nx1466), .A1 (lastDepthOut), .A2 (donttrust)) ;
    or02 ix1467 (.Y (nx1466), .A0 (LastFilterIND), .A1 (nx1477)) ;
    and04 ix77 (.Y (LastFilterIND), .A0 (nx1469), .A1 (nx1471), .A2 (nx1473), .A3 (
          nx1475)) ;
    xnor2 ix1470 (.Y (nx1469), .A0 (FilterMinus_0), .A1 (FilterCounter[0])) ;
    xnor2 ix1472 (.Y (nx1471), .A0 (FilterMinus_1), .A1 (FilterCounter[1])) ;
    xnor2 ix1474 (.Y (nx1473), .A0 (FilterMinus_2), .A1 (FilterCounter[2])) ;
    xnor2 ix1476 (.Y (nx1475), .A0 (FilterMinus_3), .A1 (FilterCounter[3])) ;
    nor04 ix1478 (.Y (nx1477), .A0 (LayerInfo[1]), .A1 (LayerInfo[2]), .A2 (
          LayerInfo[3]), .A3 (nx1479)) ;
    inv01 ix1480 (.Y (nx1479), .A (LayerInfo[0])) ;
    and04 ix55 (.Y (lastDepthOut), .A0 (nx1482), .A1 (nx1484), .A2 (nx1486), .A3 (
          nx1488)) ;
    xnor2 ix1483 (.Y (nx1482), .A0 (depthcounter[0]), .A1 (depthminus_0)) ;
    xnor2 ix1485 (.Y (nx1484), .A0 (depthcounter[1]), .A1 (depthminus_1)) ;
    xnor2 ix1487 (.Y (nx1486), .A0 (depthcounter[2]), .A1 (depthminus_2)) ;
    xnor2 ix1489 (.Y (nx1488), .A0 (depthcounter[3]), .A1 (depthminus_3)) ;
    nor03_2x ix33 (.Y (donttrust), .A0 (nx1491), .A1 (nx22), .A2 (nx24)) ;
    nand03 ix1492 (.Y (nx1491), .A0 (nx1493), .A1 (nx1495), .A2 (nx1497)) ;
    xnor2 ix1494 (.Y (nx1493), .A0 (Heightminus_1), .A1 (Heightcounter[1])) ;
    xnor2 ix1496 (.Y (nx1495), .A0 (Heightminus_4), .A1 (Heightcounter[4])) ;
    xnor2 ix1498 (.Y (nx1497), .A0 (Heightminus_0), .A1 (Heightcounter[0])) ;
    xor2 ix23 (.Y (nx22), .A0 (Heightminus_2), .A1 (Heightcounter[2])) ;
    xor2 ix25 (.Y (nx24), .A0 (Heightminus_3), .A1 (Heightcounter[3])) ;
    and02 ix123 (.Y (filter2EN), .A0 (ACKF), .A1 (nx120)) ;
    mux21_ni ix121 (.Y (nx120), .A0 (nx2), .A1 (current_state[5]), .S0 (QImgStat
             )) ;
    and02 ix133 (.Y (filter1EN), .A0 (ACKF), .A1 (nx130)) ;
    mux21_ni ix131 (.Y (nx130), .A0 (current_state[5]), .A1 (nx2), .S0 (QImgStat
             )) ;
    dffr reg_DFFCLK_dup_0 (.Q (DFFCLK), .QB (\$dummy [4]), .D (secOperand_3), .CLK (
         CLK), .R (nx108)) ;
    nand02 ix109 (.Y (nx108), .A0 (ACKF), .A1 (current_state[7])) ;
endmodule


module nBitRegister_400 ( D, CLK, RST, EN, Q ) ;

    input [399:0]D ;
    input CLK ;
    input RST ;
    input EN ;
    output [399:0]Q ;

    wire nx4838, nx4848, nx4858, nx4868, nx4878, nx4888, nx4898, nx4908, nx4918, 
         nx4928, nx4938, nx4948, nx4958, nx4968, nx4978, nx4988, nx4998, nx5008, 
         nx5018, nx5028, nx5038, nx5048, nx5058, nx5068, nx5078, nx5088, nx5098, 
         nx5108, nx5118, nx5128, nx5138, nx5148, nx5158, nx5168, nx5178, nx5188, 
         nx5198, nx5208, nx5218, nx5228, nx5238, nx5248, nx5258, nx5268, nx5278, 
         nx5288, nx5298, nx5308, nx5318, nx5328, nx5338, nx5348, nx5358, nx5368, 
         nx5378, nx5388, nx5398, nx5408, nx5418, nx5428, nx5438, nx5448, nx5458, 
         nx5468, nx5478, nx5488, nx5498, nx5508, nx5518, nx5528, nx5538, nx5548, 
         nx5558, nx5568, nx5578, nx5588, nx5598, nx5608, nx5618, nx5628, nx5638, 
         nx5648, nx5658, nx5668, nx5678, nx5688, nx5698, nx5708, nx5718, nx5728, 
         nx5738, nx5748, nx5758, nx5768, nx5778, nx5788, nx5798, nx5808, nx5818, 
         nx5828, nx5838, nx5848, nx5858, nx5868, nx5878, nx5888, nx5898, nx5908, 
         nx5918, nx5928, nx5938, nx5948, nx5958, nx5968, nx5978, nx5988, nx5998, 
         nx6008, nx6018, nx6028, nx6038, nx6048, nx6058, nx6068, nx6078, nx6088, 
         nx6098, nx6108, nx6118, nx6128, nx6138, nx6148, nx6158, nx6168, nx6178, 
         nx6188, nx6198, nx6208, nx6218, nx6228, nx6238, nx6248, nx6258, nx6268, 
         nx6278, nx6288, nx6298, nx6308, nx6318, nx6328, nx6338, nx6348, nx6358, 
         nx6368, nx6378, nx6388, nx6398, nx6408, nx6418, nx6428, nx6438, nx6448, 
         nx6458, nx6468, nx6478, nx6488, nx6498, nx6508, nx6518, nx6528, nx6538, 
         nx6548, nx6558, nx6568, nx6578, nx6588, nx6598, nx6608, nx6618, nx6628, 
         nx6638, nx6648, nx6658, nx6668, nx6678, nx6688, nx6698, nx6708, nx6718, 
         nx6728, nx6738, nx6748, nx6758, nx6768, nx6778, nx6788, nx6798, nx6808, 
         nx6818, nx6828, nx6838, nx6848, nx6858, nx6868, nx6878, nx6888, nx6898, 
         nx6908, nx6918, nx6928, nx6938, nx6948, nx6958, nx6968, nx6978, nx6988, 
         nx6998, nx7008, nx7018, nx7028, nx7038, nx7048, nx7058, nx7068, nx7078, 
         nx7088, nx7098, nx7108, nx7118, nx7128, nx7138, nx7148, nx7158, nx7168, 
         nx7178, nx7188, nx7198, nx7208, nx7218, nx7228, nx7238, nx7248, nx7258, 
         nx7268, nx7278, nx7288, nx7298, nx7308, nx7318, nx7328, nx7338, nx7348, 
         nx7358, nx7368, nx7378, nx7388, nx7398, nx7408, nx7418, nx7428, nx7438, 
         nx7448, nx7458, nx7468, nx7478, nx7488, nx7498, nx7508, nx7518, nx7528, 
         nx7538, nx7548, nx7558, nx7568, nx7578, nx7588, nx7598, nx7608, nx7618, 
         nx7628, nx7638, nx7648, nx7658, nx7668, nx7678, nx7688, nx7698, nx7708, 
         nx7718, nx7728, nx7738, nx7748, nx7758, nx7768, nx7778, nx7788, nx7798, 
         nx7808, nx7818, nx7828, nx7838, nx7848, nx7858, nx7868, nx7878, nx7888, 
         nx7898, nx7908, nx7918, nx7928, nx7938, nx7948, nx7958, nx7968, nx7978, 
         nx7988, nx7998, nx8008, nx8018, nx8028, nx8038, nx8048, nx8058, nx8068, 
         nx8078, nx8088, nx8098, nx8108, nx8118, nx8128, nx8138, nx8148, nx8158, 
         nx8168, nx8178, nx8188, nx8198, nx8208, nx8218, nx8228, nx8238, nx8248, 
         nx8258, nx8268, nx8278, nx8288, nx8298, nx8308, nx8318, nx8328, nx8338, 
         nx8348, nx8358, nx8368, nx8378, nx8388, nx8398, nx8408, nx8418, nx8428, 
         nx8438, nx8448, nx8458, nx8468, nx8478, nx8488, nx8498, nx8508, nx8518, 
         nx8528, nx8538, nx8548, nx8558, nx8568, nx8578, nx8588, nx8598, nx8608, 
         nx8618, nx8628, nx8638, nx8648, nx8658, nx8668, nx8678, nx8688, nx8698, 
         nx8708, nx8718, nx8728, nx8738, nx8748, nx8758, nx8768, nx8778, nx8788, 
         nx8798, nx8808, nx8818, nx8828, nx10045, nx10047, nx10049, nx10051, 
         nx10053, nx10055, nx10057, nx10059, nx10061, nx10063, nx10065, nx10067, 
         nx10069, nx10071, nx10073, nx10075, nx10077, nx10079, nx10081, nx10083, 
         nx10085, nx10087, nx10089, nx10091, nx10093, nx10095, nx10097, nx10099, 
         nx10101, nx10103, nx10105, nx10107, nx10109, nx10111, nx10113, nx10115, 
         nx10117, nx10119, nx10121, nx10123, nx10125, nx10127, nx10129, nx10131, 
         nx10133, nx10135, nx10137, nx10139, nx10141, nx10143, nx10145, nx10147, 
         nx10149, nx10151, nx10153, nx10155, nx10157, nx10159, nx10167, nx10169, 
         nx10171, nx10173, nx10175, nx10177, nx10179, nx10181, nx10183, nx10185, 
         nx10187, nx10189, nx10191, nx10193, nx10195, nx10197, nx10199, nx10201, 
         nx10203, nx10205, nx10207, nx10209, nx10211, nx10213, nx10215, nx10217, 
         nx10219, nx10221, nx10223, nx10225, nx10227, nx10229, nx10231, nx10233, 
         nx10235, nx10237, nx10239, nx10241, nx10243, nx10245, nx10247, nx10249, 
         nx10251, nx10253, nx10255, nx10257, nx10259, nx10261, nx10263, nx10265, 
         nx10267, nx10269, nx10271, nx10273, nx10275, nx10277, nx10279, nx10281, 
         nx10283, nx10285, nx10287, nx10289, nx10291, nx10293, nx10295, nx10297, 
         nx10299, nx10301, nx10303, nx10305, nx10307, nx10309, nx10311, nx10313, 
         nx10315, nx10317, nx10319, nx10321, nx10327, nx10329;
    wire [399:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx4838), .CLK (nx10301), .R (
         RST)) ;
    mux21_ni ix4839 (.Y (nx4838), .A0 (Q[0]), .A1 (D[0]), .S0 (nx10167)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx4848), .CLK (nx10301), .R (
         RST)) ;
    mux21_ni ix4849 (.Y (nx4848), .A0 (Q[1]), .A1 (D[1]), .S0 (nx10167)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx4858), .CLK (nx10301), .R (
         RST)) ;
    mux21_ni ix4859 (.Y (nx4858), .A0 (Q[2]), .A1 (D[2]), .S0 (nx10167)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx4868), .CLK (nx10301), .R (
         RST)) ;
    mux21_ni ix4869 (.Y (nx4868), .A0 (Q[3]), .A1 (D[3]), .S0 (nx10167)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx4878), .CLK (nx10301), .R (
         RST)) ;
    mux21_ni ix4879 (.Y (nx4878), .A0 (Q[4]), .A1 (D[4]), .S0 (nx10167)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx4888), .CLK (nx10301), .R (
         RST)) ;
    mux21_ni ix4889 (.Y (nx4888), .A0 (Q[5]), .A1 (D[5]), .S0 (nx10167)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx4898), .CLK (nx10301), .R (
         RST)) ;
    mux21_ni ix4899 (.Y (nx4898), .A0 (Q[6]), .A1 (D[6]), .S0 (nx10167)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx4908), .CLK (nx10047), .R (
         RST)) ;
    mux21_ni ix4909 (.Y (nx4908), .A0 (Q[7]), .A1 (D[7]), .S0 (nx10169)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx4918), .CLK (nx10047), .R (
         RST)) ;
    mux21_ni ix4919 (.Y (nx4918), .A0 (Q[8]), .A1 (D[8]), .S0 (nx10169)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx4928), .CLK (nx10047), .R (
         RST)) ;
    mux21_ni ix4929 (.Y (nx4928), .A0 (Q[9]), .A1 (D[9]), .S0 (nx10169)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx4938), .CLK (nx10047), 
         .R (RST)) ;
    mux21_ni ix4939 (.Y (nx4938), .A0 (Q[10]), .A1 (D[10]), .S0 (nx10169)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx4948), .CLK (nx10047), 
         .R (RST)) ;
    mux21_ni ix4949 (.Y (nx4948), .A0 (Q[11]), .A1 (D[11]), .S0 (nx10169)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx4958), .CLK (nx10047), 
         .R (RST)) ;
    mux21_ni ix4959 (.Y (nx4958), .A0 (Q[12]), .A1 (D[12]), .S0 (nx10169)) ;
    dffr reg_Q_13 (.Q (Q[13]), .QB (\$dummy [13]), .D (nx4968), .CLK (nx10047), 
         .R (RST)) ;
    mux21_ni ix4969 (.Y (nx4968), .A0 (Q[13]), .A1 (D[13]), .S0 (nx10169)) ;
    dffr reg_Q_14 (.Q (Q[14]), .QB (\$dummy [14]), .D (nx4978), .CLK (nx10049), 
         .R (RST)) ;
    mux21_ni ix4979 (.Y (nx4978), .A0 (Q[14]), .A1 (D[14]), .S0 (nx10171)) ;
    dffr reg_Q_15 (.Q (Q[15]), .QB (\$dummy [15]), .D (nx4988), .CLK (nx10049), 
         .R (RST)) ;
    mux21_ni ix4989 (.Y (nx4988), .A0 (Q[15]), .A1 (D[15]), .S0 (nx10171)) ;
    dffr reg_Q_16 (.Q (Q[16]), .QB (\$dummy [16]), .D (nx4998), .CLK (nx10049), 
         .R (RST)) ;
    mux21_ni ix4999 (.Y (nx4998), .A0 (Q[16]), .A1 (D[16]), .S0 (nx10171)) ;
    dffr reg_Q_17 (.Q (Q[17]), .QB (\$dummy [17]), .D (nx5008), .CLK (nx10049), 
         .R (RST)) ;
    mux21_ni ix5009 (.Y (nx5008), .A0 (Q[17]), .A1 (D[17]), .S0 (nx10171)) ;
    dffr reg_Q_18 (.Q (Q[18]), .QB (\$dummy [18]), .D (nx5018), .CLK (nx10049), 
         .R (RST)) ;
    mux21_ni ix5019 (.Y (nx5018), .A0 (Q[18]), .A1 (D[18]), .S0 (nx10171)) ;
    dffr reg_Q_19 (.Q (Q[19]), .QB (\$dummy [19]), .D (nx5028), .CLK (nx10049), 
         .R (RST)) ;
    mux21_ni ix5029 (.Y (nx5028), .A0 (Q[19]), .A1 (D[19]), .S0 (nx10171)) ;
    dffr reg_Q_20 (.Q (Q[20]), .QB (\$dummy [20]), .D (nx5038), .CLK (nx10049), 
         .R (RST)) ;
    mux21_ni ix5039 (.Y (nx5038), .A0 (Q[20]), .A1 (D[20]), .S0 (nx10171)) ;
    dffr reg_Q_21 (.Q (Q[21]), .QB (\$dummy [21]), .D (nx5048), .CLK (nx10051), 
         .R (RST)) ;
    mux21_ni ix5049 (.Y (nx5048), .A0 (Q[21]), .A1 (D[21]), .S0 (nx10173)) ;
    dffr reg_Q_22 (.Q (Q[22]), .QB (\$dummy [22]), .D (nx5058), .CLK (nx10051), 
         .R (RST)) ;
    mux21_ni ix5059 (.Y (nx5058), .A0 (Q[22]), .A1 (D[22]), .S0 (nx10173)) ;
    dffr reg_Q_23 (.Q (Q[23]), .QB (\$dummy [23]), .D (nx5068), .CLK (nx10051), 
         .R (RST)) ;
    mux21_ni ix5069 (.Y (nx5068), .A0 (Q[23]), .A1 (D[23]), .S0 (nx10173)) ;
    dffr reg_Q_24 (.Q (Q[24]), .QB (\$dummy [24]), .D (nx5078), .CLK (nx10051), 
         .R (RST)) ;
    mux21_ni ix5079 (.Y (nx5078), .A0 (Q[24]), .A1 (D[24]), .S0 (nx10173)) ;
    dffr reg_Q_25 (.Q (Q[25]), .QB (\$dummy [25]), .D (nx5088), .CLK (nx10051), 
         .R (RST)) ;
    mux21_ni ix5089 (.Y (nx5088), .A0 (Q[25]), .A1 (D[25]), .S0 (nx10173)) ;
    dffr reg_Q_26 (.Q (Q[26]), .QB (\$dummy [26]), .D (nx5098), .CLK (nx10051), 
         .R (RST)) ;
    mux21_ni ix5099 (.Y (nx5098), .A0 (Q[26]), .A1 (D[26]), .S0 (nx10173)) ;
    dffr reg_Q_27 (.Q (Q[27]), .QB (\$dummy [27]), .D (nx5108), .CLK (nx10051), 
         .R (RST)) ;
    mux21_ni ix5109 (.Y (nx5108), .A0 (Q[27]), .A1 (D[27]), .S0 (nx10173)) ;
    dffr reg_Q_28 (.Q (Q[28]), .QB (\$dummy [28]), .D (nx5118), .CLK (nx10053), 
         .R (RST)) ;
    mux21_ni ix5119 (.Y (nx5118), .A0 (Q[28]), .A1 (D[28]), .S0 (nx10175)) ;
    dffr reg_Q_29 (.Q (Q[29]), .QB (\$dummy [29]), .D (nx5128), .CLK (nx10053), 
         .R (RST)) ;
    mux21_ni ix5129 (.Y (nx5128), .A0 (Q[29]), .A1 (D[29]), .S0 (nx10175)) ;
    dffr reg_Q_30 (.Q (Q[30]), .QB (\$dummy [30]), .D (nx5138), .CLK (nx10053), 
         .R (RST)) ;
    mux21_ni ix5139 (.Y (nx5138), .A0 (Q[30]), .A1 (D[30]), .S0 (nx10175)) ;
    dffr reg_Q_31 (.Q (Q[31]), .QB (\$dummy [31]), .D (nx5148), .CLK (nx10053), 
         .R (RST)) ;
    mux21_ni ix5149 (.Y (nx5148), .A0 (Q[31]), .A1 (D[31]), .S0 (nx10175)) ;
    dffr reg_Q_32 (.Q (Q[32]), .QB (\$dummy [32]), .D (nx5158), .CLK (nx10053), 
         .R (RST)) ;
    mux21_ni ix5159 (.Y (nx5158), .A0 (Q[32]), .A1 (D[32]), .S0 (nx10175)) ;
    dffr reg_Q_33 (.Q (Q[33]), .QB (\$dummy [33]), .D (nx5168), .CLK (nx10053), 
         .R (RST)) ;
    mux21_ni ix5169 (.Y (nx5168), .A0 (Q[33]), .A1 (D[33]), .S0 (nx10175)) ;
    dffr reg_Q_34 (.Q (Q[34]), .QB (\$dummy [34]), .D (nx5178), .CLK (nx10053), 
         .R (RST)) ;
    mux21_ni ix5179 (.Y (nx5178), .A0 (Q[34]), .A1 (D[34]), .S0 (nx10175)) ;
    dffr reg_Q_35 (.Q (Q[35]), .QB (\$dummy [35]), .D (nx5188), .CLK (nx10055), 
         .R (RST)) ;
    mux21_ni ix5189 (.Y (nx5188), .A0 (Q[35]), .A1 (D[35]), .S0 (nx10177)) ;
    dffr reg_Q_36 (.Q (Q[36]), .QB (\$dummy [36]), .D (nx5198), .CLK (nx10055), 
         .R (RST)) ;
    mux21_ni ix5199 (.Y (nx5198), .A0 (Q[36]), .A1 (D[36]), .S0 (nx10177)) ;
    dffr reg_Q_37 (.Q (Q[37]), .QB (\$dummy [37]), .D (nx5208), .CLK (nx10055), 
         .R (RST)) ;
    mux21_ni ix5209 (.Y (nx5208), .A0 (Q[37]), .A1 (D[37]), .S0 (nx10177)) ;
    dffr reg_Q_38 (.Q (Q[38]), .QB (\$dummy [38]), .D (nx5218), .CLK (nx10055), 
         .R (RST)) ;
    mux21_ni ix5219 (.Y (nx5218), .A0 (Q[38]), .A1 (D[38]), .S0 (nx10177)) ;
    dffr reg_Q_39 (.Q (Q[39]), .QB (\$dummy [39]), .D (nx5228), .CLK (nx10055), 
         .R (RST)) ;
    mux21_ni ix5229 (.Y (nx5228), .A0 (Q[39]), .A1 (D[39]), .S0 (nx10177)) ;
    dffr reg_Q_40 (.Q (Q[40]), .QB (\$dummy [40]), .D (nx5238), .CLK (nx10055), 
         .R (RST)) ;
    mux21_ni ix5239 (.Y (nx5238), .A0 (Q[40]), .A1 (D[40]), .S0 (nx10177)) ;
    dffr reg_Q_41 (.Q (Q[41]), .QB (\$dummy [41]), .D (nx5248), .CLK (nx10055), 
         .R (RST)) ;
    mux21_ni ix5249 (.Y (nx5248), .A0 (Q[41]), .A1 (D[41]), .S0 (nx10177)) ;
    dffr reg_Q_42 (.Q (Q[42]), .QB (\$dummy [42]), .D (nx5258), .CLK (nx10057), 
         .R (RST)) ;
    mux21_ni ix5259 (.Y (nx5258), .A0 (Q[42]), .A1 (D[42]), .S0 (nx10179)) ;
    dffr reg_Q_43 (.Q (Q[43]), .QB (\$dummy [43]), .D (nx5268), .CLK (nx10057), 
         .R (RST)) ;
    mux21_ni ix5269 (.Y (nx5268), .A0 (Q[43]), .A1 (D[43]), .S0 (nx10179)) ;
    dffr reg_Q_44 (.Q (Q[44]), .QB (\$dummy [44]), .D (nx5278), .CLK (nx10057), 
         .R (RST)) ;
    mux21_ni ix5279 (.Y (nx5278), .A0 (Q[44]), .A1 (D[44]), .S0 (nx10179)) ;
    dffr reg_Q_45 (.Q (Q[45]), .QB (\$dummy [45]), .D (nx5288), .CLK (nx10057), 
         .R (RST)) ;
    mux21_ni ix5289 (.Y (nx5288), .A0 (Q[45]), .A1 (D[45]), .S0 (nx10179)) ;
    dffr reg_Q_46 (.Q (Q[46]), .QB (\$dummy [46]), .D (nx5298), .CLK (nx10057), 
         .R (RST)) ;
    mux21_ni ix5299 (.Y (nx5298), .A0 (Q[46]), .A1 (D[46]), .S0 (nx10179)) ;
    dffr reg_Q_47 (.Q (Q[47]), .QB (\$dummy [47]), .D (nx5308), .CLK (nx10057), 
         .R (RST)) ;
    mux21_ni ix5309 (.Y (nx5308), .A0 (Q[47]), .A1 (D[47]), .S0 (nx10179)) ;
    dffr reg_Q_48 (.Q (Q[48]), .QB (\$dummy [48]), .D (nx5318), .CLK (nx10057), 
         .R (RST)) ;
    mux21_ni ix5319 (.Y (nx5318), .A0 (Q[48]), .A1 (D[48]), .S0 (nx10179)) ;
    dffr reg_Q_49 (.Q (Q[49]), .QB (\$dummy [49]), .D (nx5328), .CLK (nx10059), 
         .R (RST)) ;
    mux21_ni ix5329 (.Y (nx5328), .A0 (Q[49]), .A1 (D[49]), .S0 (nx10181)) ;
    dffr reg_Q_50 (.Q (Q[50]), .QB (\$dummy [50]), .D (nx5338), .CLK (nx10059), 
         .R (RST)) ;
    mux21_ni ix5339 (.Y (nx5338), .A0 (Q[50]), .A1 (D[50]), .S0 (nx10181)) ;
    dffr reg_Q_51 (.Q (Q[51]), .QB (\$dummy [51]), .D (nx5348), .CLK (nx10059), 
         .R (RST)) ;
    mux21_ni ix5349 (.Y (nx5348), .A0 (Q[51]), .A1 (D[51]), .S0 (nx10181)) ;
    dffr reg_Q_52 (.Q (Q[52]), .QB (\$dummy [52]), .D (nx5358), .CLK (nx10059), 
         .R (RST)) ;
    mux21_ni ix5359 (.Y (nx5358), .A0 (Q[52]), .A1 (D[52]), .S0 (nx10181)) ;
    dffr reg_Q_53 (.Q (Q[53]), .QB (\$dummy [53]), .D (nx5368), .CLK (nx10059), 
         .R (RST)) ;
    mux21_ni ix5369 (.Y (nx5368), .A0 (Q[53]), .A1 (D[53]), .S0 (nx10181)) ;
    dffr reg_Q_54 (.Q (Q[54]), .QB (\$dummy [54]), .D (nx5378), .CLK (nx10059), 
         .R (RST)) ;
    mux21_ni ix5379 (.Y (nx5378), .A0 (Q[54]), .A1 (D[54]), .S0 (nx10181)) ;
    dffr reg_Q_55 (.Q (Q[55]), .QB (\$dummy [55]), .D (nx5388), .CLK (nx10059), 
         .R (RST)) ;
    mux21_ni ix5389 (.Y (nx5388), .A0 (Q[55]), .A1 (D[55]), .S0 (nx10181)) ;
    dffr reg_Q_56 (.Q (Q[56]), .QB (\$dummy [56]), .D (nx5398), .CLK (nx10061), 
         .R (RST)) ;
    mux21_ni ix5399 (.Y (nx5398), .A0 (Q[56]), .A1 (D[56]), .S0 (nx10183)) ;
    dffr reg_Q_57 (.Q (Q[57]), .QB (\$dummy [57]), .D (nx5408), .CLK (nx10061), 
         .R (RST)) ;
    mux21_ni ix5409 (.Y (nx5408), .A0 (Q[57]), .A1 (D[57]), .S0 (nx10183)) ;
    dffr reg_Q_58 (.Q (Q[58]), .QB (\$dummy [58]), .D (nx5418), .CLK (nx10061), 
         .R (RST)) ;
    mux21_ni ix5419 (.Y (nx5418), .A0 (Q[58]), .A1 (D[58]), .S0 (nx10183)) ;
    dffr reg_Q_59 (.Q (Q[59]), .QB (\$dummy [59]), .D (nx5428), .CLK (nx10061), 
         .R (RST)) ;
    mux21_ni ix5429 (.Y (nx5428), .A0 (Q[59]), .A1 (D[59]), .S0 (nx10183)) ;
    dffr reg_Q_60 (.Q (Q[60]), .QB (\$dummy [60]), .D (nx5438), .CLK (nx10061), 
         .R (RST)) ;
    mux21_ni ix5439 (.Y (nx5438), .A0 (Q[60]), .A1 (D[60]), .S0 (nx10183)) ;
    dffr reg_Q_61 (.Q (Q[61]), .QB (\$dummy [61]), .D (nx5448), .CLK (nx10061), 
         .R (RST)) ;
    mux21_ni ix5449 (.Y (nx5448), .A0 (Q[61]), .A1 (D[61]), .S0 (nx10183)) ;
    dffr reg_Q_62 (.Q (Q[62]), .QB (\$dummy [62]), .D (nx5458), .CLK (nx10061), 
         .R (RST)) ;
    mux21_ni ix5459 (.Y (nx5458), .A0 (Q[62]), .A1 (D[62]), .S0 (nx10183)) ;
    dffr reg_Q_63 (.Q (Q[63]), .QB (\$dummy [63]), .D (nx5468), .CLK (nx10063), 
         .R (RST)) ;
    mux21_ni ix5469 (.Y (nx5468), .A0 (Q[63]), .A1 (D[63]), .S0 (nx10185)) ;
    dffr reg_Q_64 (.Q (Q[64]), .QB (\$dummy [64]), .D (nx5478), .CLK (nx10063), 
         .R (RST)) ;
    mux21_ni ix5479 (.Y (nx5478), .A0 (Q[64]), .A1 (D[64]), .S0 (nx10185)) ;
    dffr reg_Q_65 (.Q (Q[65]), .QB (\$dummy [65]), .D (nx5488), .CLK (nx10063), 
         .R (RST)) ;
    mux21_ni ix5489 (.Y (nx5488), .A0 (Q[65]), .A1 (D[65]), .S0 (nx10185)) ;
    dffr reg_Q_66 (.Q (Q[66]), .QB (\$dummy [66]), .D (nx5498), .CLK (nx10063), 
         .R (RST)) ;
    mux21_ni ix5499 (.Y (nx5498), .A0 (Q[66]), .A1 (D[66]), .S0 (nx10185)) ;
    dffr reg_Q_67 (.Q (Q[67]), .QB (\$dummy [67]), .D (nx5508), .CLK (nx10063), 
         .R (RST)) ;
    mux21_ni ix5509 (.Y (nx5508), .A0 (Q[67]), .A1 (D[67]), .S0 (nx10185)) ;
    dffr reg_Q_68 (.Q (Q[68]), .QB (\$dummy [68]), .D (nx5518), .CLK (nx10063), 
         .R (RST)) ;
    mux21_ni ix5519 (.Y (nx5518), .A0 (Q[68]), .A1 (D[68]), .S0 (nx10185)) ;
    dffr reg_Q_69 (.Q (Q[69]), .QB (\$dummy [69]), .D (nx5528), .CLK (nx10063), 
         .R (RST)) ;
    mux21_ni ix5529 (.Y (nx5528), .A0 (Q[69]), .A1 (D[69]), .S0 (nx10185)) ;
    dffr reg_Q_70 (.Q (Q[70]), .QB (\$dummy [70]), .D (nx5538), .CLK (nx10065), 
         .R (RST)) ;
    mux21_ni ix5539 (.Y (nx5538), .A0 (Q[70]), .A1 (D[70]), .S0 (nx10187)) ;
    dffr reg_Q_71 (.Q (Q[71]), .QB (\$dummy [71]), .D (nx5548), .CLK (nx10065), 
         .R (RST)) ;
    mux21_ni ix5549 (.Y (nx5548), .A0 (Q[71]), .A1 (D[71]), .S0 (nx10187)) ;
    dffr reg_Q_72 (.Q (Q[72]), .QB (\$dummy [72]), .D (nx5558), .CLK (nx10065), 
         .R (RST)) ;
    mux21_ni ix5559 (.Y (nx5558), .A0 (Q[72]), .A1 (D[72]), .S0 (nx10187)) ;
    dffr reg_Q_73 (.Q (Q[73]), .QB (\$dummy [73]), .D (nx5568), .CLK (nx10065), 
         .R (RST)) ;
    mux21_ni ix5569 (.Y (nx5568), .A0 (Q[73]), .A1 (D[73]), .S0 (nx10187)) ;
    dffr reg_Q_74 (.Q (Q[74]), .QB (\$dummy [74]), .D (nx5578), .CLK (nx10065), 
         .R (RST)) ;
    mux21_ni ix5579 (.Y (nx5578), .A0 (Q[74]), .A1 (D[74]), .S0 (nx10187)) ;
    dffr reg_Q_75 (.Q (Q[75]), .QB (\$dummy [75]), .D (nx5588), .CLK (nx10065), 
         .R (RST)) ;
    mux21_ni ix5589 (.Y (nx5588), .A0 (Q[75]), .A1 (D[75]), .S0 (nx10187)) ;
    dffr reg_Q_76 (.Q (Q[76]), .QB (\$dummy [76]), .D (nx5598), .CLK (nx10065), 
         .R (RST)) ;
    mux21_ni ix5599 (.Y (nx5598), .A0 (Q[76]), .A1 (D[76]), .S0 (nx10187)) ;
    dffr reg_Q_77 (.Q (Q[77]), .QB (\$dummy [77]), .D (nx5608), .CLK (nx10067), 
         .R (RST)) ;
    mux21_ni ix5609 (.Y (nx5608), .A0 (Q[77]), .A1 (D[77]), .S0 (nx10189)) ;
    dffr reg_Q_78 (.Q (Q[78]), .QB (\$dummy [78]), .D (nx5618), .CLK (nx10067), 
         .R (RST)) ;
    mux21_ni ix5619 (.Y (nx5618), .A0 (Q[78]), .A1 (D[78]), .S0 (nx10189)) ;
    dffr reg_Q_79 (.Q (Q[79]), .QB (\$dummy [79]), .D (nx5628), .CLK (nx10067), 
         .R (RST)) ;
    mux21_ni ix5629 (.Y (nx5628), .A0 (Q[79]), .A1 (D[79]), .S0 (nx10189)) ;
    dffr reg_Q_80 (.Q (Q[80]), .QB (\$dummy [80]), .D (nx5638), .CLK (nx10067), 
         .R (RST)) ;
    mux21_ni ix5639 (.Y (nx5638), .A0 (Q[80]), .A1 (D[80]), .S0 (nx10189)) ;
    dffr reg_Q_81 (.Q (Q[81]), .QB (\$dummy [81]), .D (nx5648), .CLK (nx10067), 
         .R (RST)) ;
    mux21_ni ix5649 (.Y (nx5648), .A0 (Q[81]), .A1 (D[81]), .S0 (nx10189)) ;
    dffr reg_Q_82 (.Q (Q[82]), .QB (\$dummy [82]), .D (nx5658), .CLK (nx10067), 
         .R (RST)) ;
    mux21_ni ix5659 (.Y (nx5658), .A0 (Q[82]), .A1 (D[82]), .S0 (nx10189)) ;
    dffr reg_Q_83 (.Q (Q[83]), .QB (\$dummy [83]), .D (nx5668), .CLK (nx10067), 
         .R (RST)) ;
    mux21_ni ix5669 (.Y (nx5668), .A0 (Q[83]), .A1 (D[83]), .S0 (nx10189)) ;
    dffr reg_Q_84 (.Q (Q[84]), .QB (\$dummy [84]), .D (nx5678), .CLK (nx10069), 
         .R (RST)) ;
    mux21_ni ix5679 (.Y (nx5678), .A0 (Q[84]), .A1 (D[84]), .S0 (nx10191)) ;
    dffr reg_Q_85 (.Q (Q[85]), .QB (\$dummy [85]), .D (nx5688), .CLK (nx10069), 
         .R (RST)) ;
    mux21_ni ix5689 (.Y (nx5688), .A0 (Q[85]), .A1 (D[85]), .S0 (nx10191)) ;
    dffr reg_Q_86 (.Q (Q[86]), .QB (\$dummy [86]), .D (nx5698), .CLK (nx10069), 
         .R (RST)) ;
    mux21_ni ix5699 (.Y (nx5698), .A0 (Q[86]), .A1 (D[86]), .S0 (nx10191)) ;
    dffr reg_Q_87 (.Q (Q[87]), .QB (\$dummy [87]), .D (nx5708), .CLK (nx10069), 
         .R (RST)) ;
    mux21_ni ix5709 (.Y (nx5708), .A0 (Q[87]), .A1 (D[87]), .S0 (nx10191)) ;
    dffr reg_Q_88 (.Q (Q[88]), .QB (\$dummy [88]), .D (nx5718), .CLK (nx10069), 
         .R (RST)) ;
    mux21_ni ix5719 (.Y (nx5718), .A0 (Q[88]), .A1 (D[88]), .S0 (nx10191)) ;
    dffr reg_Q_89 (.Q (Q[89]), .QB (\$dummy [89]), .D (nx5728), .CLK (nx10069), 
         .R (RST)) ;
    mux21_ni ix5729 (.Y (nx5728), .A0 (Q[89]), .A1 (D[89]), .S0 (nx10191)) ;
    dffr reg_Q_90 (.Q (Q[90]), .QB (\$dummy [90]), .D (nx5738), .CLK (nx10069), 
         .R (RST)) ;
    mux21_ni ix5739 (.Y (nx5738), .A0 (Q[90]), .A1 (D[90]), .S0 (nx10191)) ;
    dffr reg_Q_91 (.Q (Q[91]), .QB (\$dummy [91]), .D (nx5748), .CLK (nx10071), 
         .R (RST)) ;
    mux21_ni ix5749 (.Y (nx5748), .A0 (Q[91]), .A1 (D[91]), .S0 (nx10193)) ;
    dffr reg_Q_92 (.Q (Q[92]), .QB (\$dummy [92]), .D (nx5758), .CLK (nx10071), 
         .R (RST)) ;
    mux21_ni ix5759 (.Y (nx5758), .A0 (Q[92]), .A1 (D[92]), .S0 (nx10193)) ;
    dffr reg_Q_93 (.Q (Q[93]), .QB (\$dummy [93]), .D (nx5768), .CLK (nx10071), 
         .R (RST)) ;
    mux21_ni ix5769 (.Y (nx5768), .A0 (Q[93]), .A1 (D[93]), .S0 (nx10193)) ;
    dffr reg_Q_94 (.Q (Q[94]), .QB (\$dummy [94]), .D (nx5778), .CLK (nx10071), 
         .R (RST)) ;
    mux21_ni ix5779 (.Y (nx5778), .A0 (Q[94]), .A1 (D[94]), .S0 (nx10193)) ;
    dffr reg_Q_95 (.Q (Q[95]), .QB (\$dummy [95]), .D (nx5788), .CLK (nx10071), 
         .R (RST)) ;
    mux21_ni ix5789 (.Y (nx5788), .A0 (Q[95]), .A1 (D[95]), .S0 (nx10193)) ;
    dffr reg_Q_96 (.Q (Q[96]), .QB (\$dummy [96]), .D (nx5798), .CLK (nx10071), 
         .R (RST)) ;
    mux21_ni ix5799 (.Y (nx5798), .A0 (Q[96]), .A1 (D[96]), .S0 (nx10193)) ;
    dffr reg_Q_97 (.Q (Q[97]), .QB (\$dummy [97]), .D (nx5808), .CLK (nx10071), 
         .R (RST)) ;
    mux21_ni ix5809 (.Y (nx5808), .A0 (Q[97]), .A1 (D[97]), .S0 (nx10193)) ;
    dffr reg_Q_98 (.Q (Q[98]), .QB (\$dummy [98]), .D (nx5818), .CLK (nx10073), 
         .R (RST)) ;
    mux21_ni ix5819 (.Y (nx5818), .A0 (Q[98]), .A1 (D[98]), .S0 (nx10195)) ;
    dffr reg_Q_99 (.Q (Q[99]), .QB (\$dummy [99]), .D (nx5828), .CLK (nx10073), 
         .R (RST)) ;
    mux21_ni ix5829 (.Y (nx5828), .A0 (Q[99]), .A1 (D[99]), .S0 (nx10195)) ;
    dffr reg_Q_100 (.Q (Q[100]), .QB (\$dummy [100]), .D (nx5838), .CLK (nx10073
         ), .R (RST)) ;
    mux21_ni ix5839 (.Y (nx5838), .A0 (Q[100]), .A1 (D[100]), .S0 (nx10195)) ;
    dffr reg_Q_101 (.Q (Q[101]), .QB (\$dummy [101]), .D (nx5848), .CLK (nx10073
         ), .R (RST)) ;
    mux21_ni ix5849 (.Y (nx5848), .A0 (Q[101]), .A1 (D[101]), .S0 (nx10195)) ;
    dffr reg_Q_102 (.Q (Q[102]), .QB (\$dummy [102]), .D (nx5858), .CLK (nx10073
         ), .R (RST)) ;
    mux21_ni ix5859 (.Y (nx5858), .A0 (Q[102]), .A1 (D[102]), .S0 (nx10195)) ;
    dffr reg_Q_103 (.Q (Q[103]), .QB (\$dummy [103]), .D (nx5868), .CLK (nx10073
         ), .R (RST)) ;
    mux21_ni ix5869 (.Y (nx5868), .A0 (Q[103]), .A1 (D[103]), .S0 (nx10195)) ;
    dffr reg_Q_104 (.Q (Q[104]), .QB (\$dummy [104]), .D (nx5878), .CLK (nx10073
         ), .R (RST)) ;
    mux21_ni ix5879 (.Y (nx5878), .A0 (Q[104]), .A1 (D[104]), .S0 (nx10195)) ;
    dffr reg_Q_105 (.Q (Q[105]), .QB (\$dummy [105]), .D (nx5888), .CLK (nx10075
         ), .R (RST)) ;
    mux21_ni ix5889 (.Y (nx5888), .A0 (Q[105]), .A1 (D[105]), .S0 (nx10197)) ;
    dffr reg_Q_106 (.Q (Q[106]), .QB (\$dummy [106]), .D (nx5898), .CLK (nx10075
         ), .R (RST)) ;
    mux21_ni ix5899 (.Y (nx5898), .A0 (Q[106]), .A1 (D[106]), .S0 (nx10197)) ;
    dffr reg_Q_107 (.Q (Q[107]), .QB (\$dummy [107]), .D (nx5908), .CLK (nx10075
         ), .R (RST)) ;
    mux21_ni ix5909 (.Y (nx5908), .A0 (Q[107]), .A1 (D[107]), .S0 (nx10197)) ;
    dffr reg_Q_108 (.Q (Q[108]), .QB (\$dummy [108]), .D (nx5918), .CLK (nx10075
         ), .R (RST)) ;
    mux21_ni ix5919 (.Y (nx5918), .A0 (Q[108]), .A1 (D[108]), .S0 (nx10197)) ;
    dffr reg_Q_109 (.Q (Q[109]), .QB (\$dummy [109]), .D (nx5928), .CLK (nx10075
         ), .R (RST)) ;
    mux21_ni ix5929 (.Y (nx5928), .A0 (Q[109]), .A1 (D[109]), .S0 (nx10197)) ;
    dffr reg_Q_110 (.Q (Q[110]), .QB (\$dummy [110]), .D (nx5938), .CLK (nx10075
         ), .R (RST)) ;
    mux21_ni ix5939 (.Y (nx5938), .A0 (Q[110]), .A1 (D[110]), .S0 (nx10197)) ;
    dffr reg_Q_111 (.Q (Q[111]), .QB (\$dummy [111]), .D (nx5948), .CLK (nx10075
         ), .R (RST)) ;
    mux21_ni ix5949 (.Y (nx5948), .A0 (Q[111]), .A1 (D[111]), .S0 (nx10197)) ;
    dffr reg_Q_112 (.Q (Q[112]), .QB (\$dummy [112]), .D (nx5958), .CLK (nx10077
         ), .R (RST)) ;
    mux21_ni ix5959 (.Y (nx5958), .A0 (Q[112]), .A1 (D[112]), .S0 (nx10199)) ;
    dffr reg_Q_113 (.Q (Q[113]), .QB (\$dummy [113]), .D (nx5968), .CLK (nx10077
         ), .R (RST)) ;
    mux21_ni ix5969 (.Y (nx5968), .A0 (Q[113]), .A1 (D[113]), .S0 (nx10199)) ;
    dffr reg_Q_114 (.Q (Q[114]), .QB (\$dummy [114]), .D (nx5978), .CLK (nx10077
         ), .R (RST)) ;
    mux21_ni ix5979 (.Y (nx5978), .A0 (Q[114]), .A1 (D[114]), .S0 (nx10199)) ;
    dffr reg_Q_115 (.Q (Q[115]), .QB (\$dummy [115]), .D (nx5988), .CLK (nx10077
         ), .R (RST)) ;
    mux21_ni ix5989 (.Y (nx5988), .A0 (Q[115]), .A1 (D[115]), .S0 (nx10199)) ;
    dffr reg_Q_116 (.Q (Q[116]), .QB (\$dummy [116]), .D (nx5998), .CLK (nx10077
         ), .R (RST)) ;
    mux21_ni ix5999 (.Y (nx5998), .A0 (Q[116]), .A1 (D[116]), .S0 (nx10199)) ;
    dffr reg_Q_117 (.Q (Q[117]), .QB (\$dummy [117]), .D (nx6008), .CLK (nx10077
         ), .R (RST)) ;
    mux21_ni ix6009 (.Y (nx6008), .A0 (Q[117]), .A1 (D[117]), .S0 (nx10199)) ;
    dffr reg_Q_118 (.Q (Q[118]), .QB (\$dummy [118]), .D (nx6018), .CLK (nx10077
         ), .R (RST)) ;
    mux21_ni ix6019 (.Y (nx6018), .A0 (Q[118]), .A1 (D[118]), .S0 (nx10199)) ;
    dffr reg_Q_119 (.Q (Q[119]), .QB (\$dummy [119]), .D (nx6028), .CLK (nx10079
         ), .R (RST)) ;
    mux21_ni ix6029 (.Y (nx6028), .A0 (Q[119]), .A1 (D[119]), .S0 (nx10201)) ;
    dffr reg_Q_120 (.Q (Q[120]), .QB (\$dummy [120]), .D (nx6038), .CLK (nx10079
         ), .R (RST)) ;
    mux21_ni ix6039 (.Y (nx6038), .A0 (Q[120]), .A1 (D[120]), .S0 (nx10201)) ;
    dffr reg_Q_121 (.Q (Q[121]), .QB (\$dummy [121]), .D (nx6048), .CLK (nx10079
         ), .R (RST)) ;
    mux21_ni ix6049 (.Y (nx6048), .A0 (Q[121]), .A1 (D[121]), .S0 (nx10201)) ;
    dffr reg_Q_122 (.Q (Q[122]), .QB (\$dummy [122]), .D (nx6058), .CLK (nx10079
         ), .R (RST)) ;
    mux21_ni ix6059 (.Y (nx6058), .A0 (Q[122]), .A1 (D[122]), .S0 (nx10201)) ;
    dffr reg_Q_123 (.Q (Q[123]), .QB (\$dummy [123]), .D (nx6068), .CLK (nx10079
         ), .R (RST)) ;
    mux21_ni ix6069 (.Y (nx6068), .A0 (Q[123]), .A1 (D[123]), .S0 (nx10201)) ;
    dffr reg_Q_124 (.Q (Q[124]), .QB (\$dummy [124]), .D (nx6078), .CLK (nx10079
         ), .R (RST)) ;
    mux21_ni ix6079 (.Y (nx6078), .A0 (Q[124]), .A1 (D[124]), .S0 (nx10201)) ;
    dffr reg_Q_125 (.Q (Q[125]), .QB (\$dummy [125]), .D (nx6088), .CLK (nx10079
         ), .R (RST)) ;
    mux21_ni ix6089 (.Y (nx6088), .A0 (Q[125]), .A1 (D[125]), .S0 (nx10201)) ;
    dffr reg_Q_126 (.Q (Q[126]), .QB (\$dummy [126]), .D (nx6098), .CLK (nx10081
         ), .R (RST)) ;
    mux21_ni ix6099 (.Y (nx6098), .A0 (Q[126]), .A1 (D[126]), .S0 (nx10203)) ;
    dffr reg_Q_127 (.Q (Q[127]), .QB (\$dummy [127]), .D (nx6108), .CLK (nx10081
         ), .R (RST)) ;
    mux21_ni ix6109 (.Y (nx6108), .A0 (Q[127]), .A1 (D[127]), .S0 (nx10203)) ;
    dffr reg_Q_128 (.Q (Q[128]), .QB (\$dummy [128]), .D (nx6118), .CLK (nx10081
         ), .R (RST)) ;
    mux21_ni ix6119 (.Y (nx6118), .A0 (Q[128]), .A1 (D[128]), .S0 (nx10203)) ;
    dffr reg_Q_129 (.Q (Q[129]), .QB (\$dummy [129]), .D (nx6128), .CLK (nx10081
         ), .R (RST)) ;
    mux21_ni ix6129 (.Y (nx6128), .A0 (Q[129]), .A1 (D[129]), .S0 (nx10203)) ;
    dffr reg_Q_130 (.Q (Q[130]), .QB (\$dummy [130]), .D (nx6138), .CLK (nx10081
         ), .R (RST)) ;
    mux21_ni ix6139 (.Y (nx6138), .A0 (Q[130]), .A1 (D[130]), .S0 (nx10203)) ;
    dffr reg_Q_131 (.Q (Q[131]), .QB (\$dummy [131]), .D (nx6148), .CLK (nx10081
         ), .R (RST)) ;
    mux21_ni ix6149 (.Y (nx6148), .A0 (Q[131]), .A1 (D[131]), .S0 (nx10203)) ;
    dffr reg_Q_132 (.Q (Q[132]), .QB (\$dummy [132]), .D (nx6158), .CLK (nx10081
         ), .R (RST)) ;
    mux21_ni ix6159 (.Y (nx6158), .A0 (Q[132]), .A1 (D[132]), .S0 (nx10203)) ;
    dffr reg_Q_133 (.Q (Q[133]), .QB (\$dummy [133]), .D (nx6168), .CLK (nx10083
         ), .R (RST)) ;
    mux21_ni ix6169 (.Y (nx6168), .A0 (Q[133]), .A1 (D[133]), .S0 (nx10205)) ;
    dffr reg_Q_134 (.Q (Q[134]), .QB (\$dummy [134]), .D (nx6178), .CLK (nx10083
         ), .R (RST)) ;
    mux21_ni ix6179 (.Y (nx6178), .A0 (Q[134]), .A1 (D[134]), .S0 (nx10205)) ;
    dffr reg_Q_135 (.Q (Q[135]), .QB (\$dummy [135]), .D (nx6188), .CLK (nx10083
         ), .R (RST)) ;
    mux21_ni ix6189 (.Y (nx6188), .A0 (Q[135]), .A1 (D[135]), .S0 (nx10205)) ;
    dffr reg_Q_136 (.Q (Q[136]), .QB (\$dummy [136]), .D (nx6198), .CLK (nx10083
         ), .R (RST)) ;
    mux21_ni ix6199 (.Y (nx6198), .A0 (Q[136]), .A1 (D[136]), .S0 (nx10205)) ;
    dffr reg_Q_137 (.Q (Q[137]), .QB (\$dummy [137]), .D (nx6208), .CLK (nx10083
         ), .R (RST)) ;
    mux21_ni ix6209 (.Y (nx6208), .A0 (Q[137]), .A1 (D[137]), .S0 (nx10205)) ;
    dffr reg_Q_138 (.Q (Q[138]), .QB (\$dummy [138]), .D (nx6218), .CLK (nx10083
         ), .R (RST)) ;
    mux21_ni ix6219 (.Y (nx6218), .A0 (Q[138]), .A1 (D[138]), .S0 (nx10205)) ;
    dffr reg_Q_139 (.Q (Q[139]), .QB (\$dummy [139]), .D (nx6228), .CLK (nx10083
         ), .R (RST)) ;
    mux21_ni ix6229 (.Y (nx6228), .A0 (Q[139]), .A1 (D[139]), .S0 (nx10205)) ;
    dffr reg_Q_140 (.Q (Q[140]), .QB (\$dummy [140]), .D (nx6238), .CLK (nx10085
         ), .R (RST)) ;
    mux21_ni ix6239 (.Y (nx6238), .A0 (Q[140]), .A1 (D[140]), .S0 (nx10207)) ;
    dffr reg_Q_141 (.Q (Q[141]), .QB (\$dummy [141]), .D (nx6248), .CLK (nx10085
         ), .R (RST)) ;
    mux21_ni ix6249 (.Y (nx6248), .A0 (Q[141]), .A1 (D[141]), .S0 (nx10207)) ;
    dffr reg_Q_142 (.Q (Q[142]), .QB (\$dummy [142]), .D (nx6258), .CLK (nx10085
         ), .R (RST)) ;
    mux21_ni ix6259 (.Y (nx6258), .A0 (Q[142]), .A1 (D[142]), .S0 (nx10207)) ;
    dffr reg_Q_143 (.Q (Q[143]), .QB (\$dummy [143]), .D (nx6268), .CLK (nx10085
         ), .R (RST)) ;
    mux21_ni ix6269 (.Y (nx6268), .A0 (Q[143]), .A1 (D[143]), .S0 (nx10207)) ;
    dffr reg_Q_144 (.Q (Q[144]), .QB (\$dummy [144]), .D (nx6278), .CLK (nx10085
         ), .R (RST)) ;
    mux21_ni ix6279 (.Y (nx6278), .A0 (Q[144]), .A1 (D[144]), .S0 (nx10207)) ;
    dffr reg_Q_145 (.Q (Q[145]), .QB (\$dummy [145]), .D (nx6288), .CLK (nx10085
         ), .R (RST)) ;
    mux21_ni ix6289 (.Y (nx6288), .A0 (Q[145]), .A1 (D[145]), .S0 (nx10207)) ;
    dffr reg_Q_146 (.Q (Q[146]), .QB (\$dummy [146]), .D (nx6298), .CLK (nx10085
         ), .R (RST)) ;
    mux21_ni ix6299 (.Y (nx6298), .A0 (Q[146]), .A1 (D[146]), .S0 (nx10207)) ;
    dffr reg_Q_147 (.Q (Q[147]), .QB (\$dummy [147]), .D (nx6308), .CLK (nx10087
         ), .R (RST)) ;
    mux21_ni ix6309 (.Y (nx6308), .A0 (Q[147]), .A1 (D[147]), .S0 (nx10209)) ;
    dffr reg_Q_148 (.Q (Q[148]), .QB (\$dummy [148]), .D (nx6318), .CLK (nx10087
         ), .R (RST)) ;
    mux21_ni ix6319 (.Y (nx6318), .A0 (Q[148]), .A1 (D[148]), .S0 (nx10209)) ;
    dffr reg_Q_149 (.Q (Q[149]), .QB (\$dummy [149]), .D (nx6328), .CLK (nx10087
         ), .R (RST)) ;
    mux21_ni ix6329 (.Y (nx6328), .A0 (Q[149]), .A1 (D[149]), .S0 (nx10209)) ;
    dffr reg_Q_150 (.Q (Q[150]), .QB (\$dummy [150]), .D (nx6338), .CLK (nx10087
         ), .R (RST)) ;
    mux21_ni ix6339 (.Y (nx6338), .A0 (Q[150]), .A1 (D[150]), .S0 (nx10209)) ;
    dffr reg_Q_151 (.Q (Q[151]), .QB (\$dummy [151]), .D (nx6348), .CLK (nx10087
         ), .R (RST)) ;
    mux21_ni ix6349 (.Y (nx6348), .A0 (Q[151]), .A1 (D[151]), .S0 (nx10209)) ;
    dffr reg_Q_152 (.Q (Q[152]), .QB (\$dummy [152]), .D (nx6358), .CLK (nx10087
         ), .R (RST)) ;
    mux21_ni ix6359 (.Y (nx6358), .A0 (Q[152]), .A1 (D[152]), .S0 (nx10209)) ;
    dffr reg_Q_153 (.Q (Q[153]), .QB (\$dummy [153]), .D (nx6368), .CLK (nx10087
         ), .R (RST)) ;
    mux21_ni ix6369 (.Y (nx6368), .A0 (Q[153]), .A1 (D[153]), .S0 (nx10209)) ;
    dffr reg_Q_154 (.Q (Q[154]), .QB (\$dummy [154]), .D (nx6378), .CLK (nx10089
         ), .R (RST)) ;
    mux21_ni ix6379 (.Y (nx6378), .A0 (Q[154]), .A1 (D[154]), .S0 (nx10211)) ;
    dffr reg_Q_155 (.Q (Q[155]), .QB (\$dummy [155]), .D (nx6388), .CLK (nx10089
         ), .R (RST)) ;
    mux21_ni ix6389 (.Y (nx6388), .A0 (Q[155]), .A1 (D[155]), .S0 (nx10211)) ;
    dffr reg_Q_156 (.Q (Q[156]), .QB (\$dummy [156]), .D (nx6398), .CLK (nx10089
         ), .R (RST)) ;
    mux21_ni ix6399 (.Y (nx6398), .A0 (Q[156]), .A1 (D[156]), .S0 (nx10211)) ;
    dffr reg_Q_157 (.Q (Q[157]), .QB (\$dummy [157]), .D (nx6408), .CLK (nx10089
         ), .R (RST)) ;
    mux21_ni ix6409 (.Y (nx6408), .A0 (Q[157]), .A1 (D[157]), .S0 (nx10211)) ;
    dffr reg_Q_158 (.Q (Q[158]), .QB (\$dummy [158]), .D (nx6418), .CLK (nx10089
         ), .R (RST)) ;
    mux21_ni ix6419 (.Y (nx6418), .A0 (Q[158]), .A1 (D[158]), .S0 (nx10211)) ;
    dffr reg_Q_159 (.Q (Q[159]), .QB (\$dummy [159]), .D (nx6428), .CLK (nx10089
         ), .R (RST)) ;
    mux21_ni ix6429 (.Y (nx6428), .A0 (Q[159]), .A1 (D[159]), .S0 (nx10211)) ;
    dffr reg_Q_160 (.Q (Q[160]), .QB (\$dummy [160]), .D (nx6438), .CLK (nx10089
         ), .R (RST)) ;
    mux21_ni ix6439 (.Y (nx6438), .A0 (Q[160]), .A1 (D[160]), .S0 (nx10211)) ;
    dffr reg_Q_161 (.Q (Q[161]), .QB (\$dummy [161]), .D (nx6448), .CLK (nx10091
         ), .R (RST)) ;
    mux21_ni ix6449 (.Y (nx6448), .A0 (Q[161]), .A1 (D[161]), .S0 (nx10213)) ;
    dffr reg_Q_162 (.Q (Q[162]), .QB (\$dummy [162]), .D (nx6458), .CLK (nx10091
         ), .R (RST)) ;
    mux21_ni ix6459 (.Y (nx6458), .A0 (Q[162]), .A1 (D[162]), .S0 (nx10213)) ;
    dffr reg_Q_163 (.Q (Q[163]), .QB (\$dummy [163]), .D (nx6468), .CLK (nx10091
         ), .R (RST)) ;
    mux21_ni ix6469 (.Y (nx6468), .A0 (Q[163]), .A1 (D[163]), .S0 (nx10213)) ;
    dffr reg_Q_164 (.Q (Q[164]), .QB (\$dummy [164]), .D (nx6478), .CLK (nx10091
         ), .R (RST)) ;
    mux21_ni ix6479 (.Y (nx6478), .A0 (Q[164]), .A1 (D[164]), .S0 (nx10213)) ;
    dffr reg_Q_165 (.Q (Q[165]), .QB (\$dummy [165]), .D (nx6488), .CLK (nx10091
         ), .R (RST)) ;
    mux21_ni ix6489 (.Y (nx6488), .A0 (Q[165]), .A1 (D[165]), .S0 (nx10213)) ;
    dffr reg_Q_166 (.Q (Q[166]), .QB (\$dummy [166]), .D (nx6498), .CLK (nx10091
         ), .R (RST)) ;
    mux21_ni ix6499 (.Y (nx6498), .A0 (Q[166]), .A1 (D[166]), .S0 (nx10213)) ;
    dffr reg_Q_167 (.Q (Q[167]), .QB (\$dummy [167]), .D (nx6508), .CLK (nx10091
         ), .R (RST)) ;
    mux21_ni ix6509 (.Y (nx6508), .A0 (Q[167]), .A1 (D[167]), .S0 (nx10213)) ;
    dffr reg_Q_168 (.Q (Q[168]), .QB (\$dummy [168]), .D (nx6518), .CLK (nx10093
         ), .R (RST)) ;
    mux21_ni ix6519 (.Y (nx6518), .A0 (Q[168]), .A1 (D[168]), .S0 (nx10215)) ;
    dffr reg_Q_169 (.Q (Q[169]), .QB (\$dummy [169]), .D (nx6528), .CLK (nx10093
         ), .R (RST)) ;
    mux21_ni ix6529 (.Y (nx6528), .A0 (Q[169]), .A1 (D[169]), .S0 (nx10215)) ;
    dffr reg_Q_170 (.Q (Q[170]), .QB (\$dummy [170]), .D (nx6538), .CLK (nx10093
         ), .R (RST)) ;
    mux21_ni ix6539 (.Y (nx6538), .A0 (Q[170]), .A1 (D[170]), .S0 (nx10215)) ;
    dffr reg_Q_171 (.Q (Q[171]), .QB (\$dummy [171]), .D (nx6548), .CLK (nx10093
         ), .R (RST)) ;
    mux21_ni ix6549 (.Y (nx6548), .A0 (Q[171]), .A1 (D[171]), .S0 (nx10215)) ;
    dffr reg_Q_172 (.Q (Q[172]), .QB (\$dummy [172]), .D (nx6558), .CLK (nx10093
         ), .R (RST)) ;
    mux21_ni ix6559 (.Y (nx6558), .A0 (Q[172]), .A1 (D[172]), .S0 (nx10215)) ;
    dffr reg_Q_173 (.Q (Q[173]), .QB (\$dummy [173]), .D (nx6568), .CLK (nx10093
         ), .R (RST)) ;
    mux21_ni ix6569 (.Y (nx6568), .A0 (Q[173]), .A1 (D[173]), .S0 (nx10215)) ;
    dffr reg_Q_174 (.Q (Q[174]), .QB (\$dummy [174]), .D (nx6578), .CLK (nx10093
         ), .R (RST)) ;
    mux21_ni ix6579 (.Y (nx6578), .A0 (Q[174]), .A1 (D[174]), .S0 (nx10215)) ;
    dffr reg_Q_175 (.Q (Q[175]), .QB (\$dummy [175]), .D (nx6588), .CLK (nx10095
         ), .R (RST)) ;
    mux21_ni ix6589 (.Y (nx6588), .A0 (Q[175]), .A1 (D[175]), .S0 (nx10217)) ;
    dffr reg_Q_176 (.Q (Q[176]), .QB (\$dummy [176]), .D (nx6598), .CLK (nx10095
         ), .R (RST)) ;
    mux21_ni ix6599 (.Y (nx6598), .A0 (Q[176]), .A1 (D[176]), .S0 (nx10217)) ;
    dffr reg_Q_177 (.Q (Q[177]), .QB (\$dummy [177]), .D (nx6608), .CLK (nx10095
         ), .R (RST)) ;
    mux21_ni ix6609 (.Y (nx6608), .A0 (Q[177]), .A1 (D[177]), .S0 (nx10217)) ;
    dffr reg_Q_178 (.Q (Q[178]), .QB (\$dummy [178]), .D (nx6618), .CLK (nx10095
         ), .R (RST)) ;
    mux21_ni ix6619 (.Y (nx6618), .A0 (Q[178]), .A1 (D[178]), .S0 (nx10217)) ;
    dffr reg_Q_179 (.Q (Q[179]), .QB (\$dummy [179]), .D (nx6628), .CLK (nx10095
         ), .R (RST)) ;
    mux21_ni ix6629 (.Y (nx6628), .A0 (Q[179]), .A1 (D[179]), .S0 (nx10217)) ;
    dffr reg_Q_180 (.Q (Q[180]), .QB (\$dummy [180]), .D (nx6638), .CLK (nx10095
         ), .R (RST)) ;
    mux21_ni ix6639 (.Y (nx6638), .A0 (Q[180]), .A1 (D[180]), .S0 (nx10217)) ;
    dffr reg_Q_181 (.Q (Q[181]), .QB (\$dummy [181]), .D (nx6648), .CLK (nx10095
         ), .R (RST)) ;
    mux21_ni ix6649 (.Y (nx6648), .A0 (Q[181]), .A1 (D[181]), .S0 (nx10217)) ;
    dffr reg_Q_182 (.Q (Q[182]), .QB (\$dummy [182]), .D (nx6658), .CLK (nx10097
         ), .R (RST)) ;
    mux21_ni ix6659 (.Y (nx6658), .A0 (Q[182]), .A1 (D[182]), .S0 (nx10219)) ;
    dffr reg_Q_183 (.Q (Q[183]), .QB (\$dummy [183]), .D (nx6668), .CLK (nx10097
         ), .R (RST)) ;
    mux21_ni ix6669 (.Y (nx6668), .A0 (Q[183]), .A1 (D[183]), .S0 (nx10219)) ;
    dffr reg_Q_184 (.Q (Q[184]), .QB (\$dummy [184]), .D (nx6678), .CLK (nx10097
         ), .R (RST)) ;
    mux21_ni ix6679 (.Y (nx6678), .A0 (Q[184]), .A1 (D[184]), .S0 (nx10219)) ;
    dffr reg_Q_185 (.Q (Q[185]), .QB (\$dummy [185]), .D (nx6688), .CLK (nx10097
         ), .R (RST)) ;
    mux21_ni ix6689 (.Y (nx6688), .A0 (Q[185]), .A1 (D[185]), .S0 (nx10219)) ;
    dffr reg_Q_186 (.Q (Q[186]), .QB (\$dummy [186]), .D (nx6698), .CLK (nx10097
         ), .R (RST)) ;
    mux21_ni ix6699 (.Y (nx6698), .A0 (Q[186]), .A1 (D[186]), .S0 (nx10219)) ;
    dffr reg_Q_187 (.Q (Q[187]), .QB (\$dummy [187]), .D (nx6708), .CLK (nx10097
         ), .R (RST)) ;
    mux21_ni ix6709 (.Y (nx6708), .A0 (Q[187]), .A1 (D[187]), .S0 (nx10219)) ;
    dffr reg_Q_188 (.Q (Q[188]), .QB (\$dummy [188]), .D (nx6718), .CLK (nx10097
         ), .R (RST)) ;
    mux21_ni ix6719 (.Y (nx6718), .A0 (Q[188]), .A1 (D[188]), .S0 (nx10219)) ;
    dffr reg_Q_189 (.Q (Q[189]), .QB (\$dummy [189]), .D (nx6728), .CLK (nx10099
         ), .R (RST)) ;
    mux21_ni ix6729 (.Y (nx6728), .A0 (Q[189]), .A1 (D[189]), .S0 (nx10221)) ;
    dffr reg_Q_190 (.Q (Q[190]), .QB (\$dummy [190]), .D (nx6738), .CLK (nx10099
         ), .R (RST)) ;
    mux21_ni ix6739 (.Y (nx6738), .A0 (Q[190]), .A1 (D[190]), .S0 (nx10221)) ;
    dffr reg_Q_191 (.Q (Q[191]), .QB (\$dummy [191]), .D (nx6748), .CLK (nx10099
         ), .R (RST)) ;
    mux21_ni ix6749 (.Y (nx6748), .A0 (Q[191]), .A1 (D[191]), .S0 (nx10221)) ;
    dffr reg_Q_192 (.Q (Q[192]), .QB (\$dummy [192]), .D (nx6758), .CLK (nx10099
         ), .R (RST)) ;
    mux21_ni ix6759 (.Y (nx6758), .A0 (Q[192]), .A1 (D[192]), .S0 (nx10221)) ;
    dffr reg_Q_193 (.Q (Q[193]), .QB (\$dummy [193]), .D (nx6768), .CLK (nx10099
         ), .R (RST)) ;
    mux21_ni ix6769 (.Y (nx6768), .A0 (Q[193]), .A1 (D[193]), .S0 (nx10221)) ;
    dffr reg_Q_194 (.Q (Q[194]), .QB (\$dummy [194]), .D (nx6778), .CLK (nx10099
         ), .R (RST)) ;
    mux21_ni ix6779 (.Y (nx6778), .A0 (Q[194]), .A1 (D[194]), .S0 (nx10221)) ;
    dffr reg_Q_195 (.Q (Q[195]), .QB (\$dummy [195]), .D (nx6788), .CLK (nx10099
         ), .R (RST)) ;
    mux21_ni ix6789 (.Y (nx6788), .A0 (Q[195]), .A1 (D[195]), .S0 (nx10221)) ;
    dffr reg_Q_196 (.Q (Q[196]), .QB (\$dummy [196]), .D (nx6798), .CLK (nx10101
         ), .R (RST)) ;
    mux21_ni ix6799 (.Y (nx6798), .A0 (Q[196]), .A1 (D[196]), .S0 (nx10223)) ;
    dffr reg_Q_197 (.Q (Q[197]), .QB (\$dummy [197]), .D (nx6808), .CLK (nx10101
         ), .R (RST)) ;
    mux21_ni ix6809 (.Y (nx6808), .A0 (Q[197]), .A1 (D[197]), .S0 (nx10223)) ;
    dffr reg_Q_198 (.Q (Q[198]), .QB (\$dummy [198]), .D (nx6818), .CLK (nx10101
         ), .R (RST)) ;
    mux21_ni ix6819 (.Y (nx6818), .A0 (Q[198]), .A1 (D[198]), .S0 (nx10223)) ;
    dffr reg_Q_199 (.Q (Q[199]), .QB (\$dummy [199]), .D (nx6828), .CLK (nx10101
         ), .R (RST)) ;
    mux21_ni ix6829 (.Y (nx6828), .A0 (Q[199]), .A1 (D[199]), .S0 (nx10223)) ;
    dffr reg_Q_200 (.Q (Q[200]), .QB (\$dummy [200]), .D (nx6838), .CLK (nx10101
         ), .R (RST)) ;
    mux21_ni ix6839 (.Y (nx6838), .A0 (Q[200]), .A1 (D[200]), .S0 (nx10223)) ;
    dffr reg_Q_201 (.Q (Q[201]), .QB (\$dummy [201]), .D (nx6848), .CLK (nx10101
         ), .R (RST)) ;
    mux21_ni ix6849 (.Y (nx6848), .A0 (Q[201]), .A1 (D[201]), .S0 (nx10223)) ;
    dffr reg_Q_202 (.Q (Q[202]), .QB (\$dummy [202]), .D (nx6858), .CLK (nx10101
         ), .R (RST)) ;
    mux21_ni ix6859 (.Y (nx6858), .A0 (Q[202]), .A1 (D[202]), .S0 (nx10223)) ;
    dffr reg_Q_203 (.Q (Q[203]), .QB (\$dummy [203]), .D (nx6868), .CLK (nx10103
         ), .R (RST)) ;
    mux21_ni ix6869 (.Y (nx6868), .A0 (Q[203]), .A1 (D[203]), .S0 (nx10225)) ;
    dffr reg_Q_204 (.Q (Q[204]), .QB (\$dummy [204]), .D (nx6878), .CLK (nx10103
         ), .R (RST)) ;
    mux21_ni ix6879 (.Y (nx6878), .A0 (Q[204]), .A1 (D[204]), .S0 (nx10225)) ;
    dffr reg_Q_205 (.Q (Q[205]), .QB (\$dummy [205]), .D (nx6888), .CLK (nx10103
         ), .R (RST)) ;
    mux21_ni ix6889 (.Y (nx6888), .A0 (Q[205]), .A1 (D[205]), .S0 (nx10225)) ;
    dffr reg_Q_206 (.Q (Q[206]), .QB (\$dummy [206]), .D (nx6898), .CLK (nx10103
         ), .R (RST)) ;
    mux21_ni ix6899 (.Y (nx6898), .A0 (Q[206]), .A1 (D[206]), .S0 (nx10225)) ;
    dffr reg_Q_207 (.Q (Q[207]), .QB (\$dummy [207]), .D (nx6908), .CLK (nx10103
         ), .R (RST)) ;
    mux21_ni ix6909 (.Y (nx6908), .A0 (Q[207]), .A1 (D[207]), .S0 (nx10225)) ;
    dffr reg_Q_208 (.Q (Q[208]), .QB (\$dummy [208]), .D (nx6918), .CLK (nx10103
         ), .R (RST)) ;
    mux21_ni ix6919 (.Y (nx6918), .A0 (Q[208]), .A1 (D[208]), .S0 (nx10225)) ;
    dffr reg_Q_209 (.Q (Q[209]), .QB (\$dummy [209]), .D (nx6928), .CLK (nx10103
         ), .R (RST)) ;
    mux21_ni ix6929 (.Y (nx6928), .A0 (Q[209]), .A1 (D[209]), .S0 (nx10225)) ;
    dffr reg_Q_210 (.Q (Q[210]), .QB (\$dummy [210]), .D (nx6938), .CLK (nx10105
         ), .R (RST)) ;
    mux21_ni ix6939 (.Y (nx6938), .A0 (Q[210]), .A1 (D[210]), .S0 (nx10227)) ;
    dffr reg_Q_211 (.Q (Q[211]), .QB (\$dummy [211]), .D (nx6948), .CLK (nx10105
         ), .R (RST)) ;
    mux21_ni ix6949 (.Y (nx6948), .A0 (Q[211]), .A1 (D[211]), .S0 (nx10227)) ;
    dffr reg_Q_212 (.Q (Q[212]), .QB (\$dummy [212]), .D (nx6958), .CLK (nx10105
         ), .R (RST)) ;
    mux21_ni ix6959 (.Y (nx6958), .A0 (Q[212]), .A1 (D[212]), .S0 (nx10227)) ;
    dffr reg_Q_213 (.Q (Q[213]), .QB (\$dummy [213]), .D (nx6968), .CLK (nx10105
         ), .R (RST)) ;
    mux21_ni ix6969 (.Y (nx6968), .A0 (Q[213]), .A1 (D[213]), .S0 (nx10227)) ;
    dffr reg_Q_214 (.Q (Q[214]), .QB (\$dummy [214]), .D (nx6978), .CLK (nx10105
         ), .R (RST)) ;
    mux21_ni ix6979 (.Y (nx6978), .A0 (Q[214]), .A1 (D[214]), .S0 (nx10227)) ;
    dffr reg_Q_215 (.Q (Q[215]), .QB (\$dummy [215]), .D (nx6988), .CLK (nx10105
         ), .R (RST)) ;
    mux21_ni ix6989 (.Y (nx6988), .A0 (Q[215]), .A1 (D[215]), .S0 (nx10227)) ;
    dffr reg_Q_216 (.Q (Q[216]), .QB (\$dummy [216]), .D (nx6998), .CLK (nx10105
         ), .R (RST)) ;
    mux21_ni ix6999 (.Y (nx6998), .A0 (Q[216]), .A1 (D[216]), .S0 (nx10227)) ;
    dffr reg_Q_217 (.Q (Q[217]), .QB (\$dummy [217]), .D (nx7008), .CLK (nx10107
         ), .R (RST)) ;
    mux21_ni ix7009 (.Y (nx7008), .A0 (Q[217]), .A1 (D[217]), .S0 (nx10229)) ;
    dffr reg_Q_218 (.Q (Q[218]), .QB (\$dummy [218]), .D (nx7018), .CLK (nx10107
         ), .R (RST)) ;
    mux21_ni ix7019 (.Y (nx7018), .A0 (Q[218]), .A1 (D[218]), .S0 (nx10229)) ;
    dffr reg_Q_219 (.Q (Q[219]), .QB (\$dummy [219]), .D (nx7028), .CLK (nx10107
         ), .R (RST)) ;
    mux21_ni ix7029 (.Y (nx7028), .A0 (Q[219]), .A1 (D[219]), .S0 (nx10229)) ;
    dffr reg_Q_220 (.Q (Q[220]), .QB (\$dummy [220]), .D (nx7038), .CLK (nx10107
         ), .R (RST)) ;
    mux21_ni ix7039 (.Y (nx7038), .A0 (Q[220]), .A1 (D[220]), .S0 (nx10229)) ;
    dffr reg_Q_221 (.Q (Q[221]), .QB (\$dummy [221]), .D (nx7048), .CLK (nx10107
         ), .R (RST)) ;
    mux21_ni ix7049 (.Y (nx7048), .A0 (Q[221]), .A1 (D[221]), .S0 (nx10229)) ;
    dffr reg_Q_222 (.Q (Q[222]), .QB (\$dummy [222]), .D (nx7058), .CLK (nx10107
         ), .R (RST)) ;
    mux21_ni ix7059 (.Y (nx7058), .A0 (Q[222]), .A1 (D[222]), .S0 (nx10229)) ;
    dffr reg_Q_223 (.Q (Q[223]), .QB (\$dummy [223]), .D (nx7068), .CLK (nx10107
         ), .R (RST)) ;
    mux21_ni ix7069 (.Y (nx7068), .A0 (Q[223]), .A1 (D[223]), .S0 (nx10229)) ;
    dffr reg_Q_224 (.Q (Q[224]), .QB (\$dummy [224]), .D (nx7078), .CLK (nx10109
         ), .R (RST)) ;
    mux21_ni ix7079 (.Y (nx7078), .A0 (Q[224]), .A1 (D[224]), .S0 (nx10231)) ;
    dffr reg_Q_225 (.Q (Q[225]), .QB (\$dummy [225]), .D (nx7088), .CLK (nx10109
         ), .R (RST)) ;
    mux21_ni ix7089 (.Y (nx7088), .A0 (Q[225]), .A1 (D[225]), .S0 (nx10231)) ;
    dffr reg_Q_226 (.Q (Q[226]), .QB (\$dummy [226]), .D (nx7098), .CLK (nx10109
         ), .R (RST)) ;
    mux21_ni ix7099 (.Y (nx7098), .A0 (Q[226]), .A1 (D[226]), .S0 (nx10231)) ;
    dffr reg_Q_227 (.Q (Q[227]), .QB (\$dummy [227]), .D (nx7108), .CLK (nx10109
         ), .R (RST)) ;
    mux21_ni ix7109 (.Y (nx7108), .A0 (Q[227]), .A1 (D[227]), .S0 (nx10231)) ;
    dffr reg_Q_228 (.Q (Q[228]), .QB (\$dummy [228]), .D (nx7118), .CLK (nx10109
         ), .R (RST)) ;
    mux21_ni ix7119 (.Y (nx7118), .A0 (Q[228]), .A1 (D[228]), .S0 (nx10231)) ;
    dffr reg_Q_229 (.Q (Q[229]), .QB (\$dummy [229]), .D (nx7128), .CLK (nx10109
         ), .R (RST)) ;
    mux21_ni ix7129 (.Y (nx7128), .A0 (Q[229]), .A1 (D[229]), .S0 (nx10231)) ;
    dffr reg_Q_230 (.Q (Q[230]), .QB (\$dummy [230]), .D (nx7138), .CLK (nx10109
         ), .R (RST)) ;
    mux21_ni ix7139 (.Y (nx7138), .A0 (Q[230]), .A1 (D[230]), .S0 (nx10231)) ;
    dffr reg_Q_231 (.Q (Q[231]), .QB (\$dummy [231]), .D (nx7148), .CLK (nx10111
         ), .R (RST)) ;
    mux21_ni ix7149 (.Y (nx7148), .A0 (Q[231]), .A1 (D[231]), .S0 (nx10233)) ;
    dffr reg_Q_232 (.Q (Q[232]), .QB (\$dummy [232]), .D (nx7158), .CLK (nx10111
         ), .R (RST)) ;
    mux21_ni ix7159 (.Y (nx7158), .A0 (Q[232]), .A1 (D[232]), .S0 (nx10233)) ;
    dffr reg_Q_233 (.Q (Q[233]), .QB (\$dummy [233]), .D (nx7168), .CLK (nx10111
         ), .R (RST)) ;
    mux21_ni ix7169 (.Y (nx7168), .A0 (Q[233]), .A1 (D[233]), .S0 (nx10233)) ;
    dffr reg_Q_234 (.Q (Q[234]), .QB (\$dummy [234]), .D (nx7178), .CLK (nx10111
         ), .R (RST)) ;
    mux21_ni ix7179 (.Y (nx7178), .A0 (Q[234]), .A1 (D[234]), .S0 (nx10233)) ;
    dffr reg_Q_235 (.Q (Q[235]), .QB (\$dummy [235]), .D (nx7188), .CLK (nx10111
         ), .R (RST)) ;
    mux21_ni ix7189 (.Y (nx7188), .A0 (Q[235]), .A1 (D[235]), .S0 (nx10233)) ;
    dffr reg_Q_236 (.Q (Q[236]), .QB (\$dummy [236]), .D (nx7198), .CLK (nx10111
         ), .R (RST)) ;
    mux21_ni ix7199 (.Y (nx7198), .A0 (Q[236]), .A1 (D[236]), .S0 (nx10233)) ;
    dffr reg_Q_237 (.Q (Q[237]), .QB (\$dummy [237]), .D (nx7208), .CLK (nx10111
         ), .R (RST)) ;
    mux21_ni ix7209 (.Y (nx7208), .A0 (Q[237]), .A1 (D[237]), .S0 (nx10233)) ;
    dffr reg_Q_238 (.Q (Q[238]), .QB (\$dummy [238]), .D (nx7218), .CLK (nx10113
         ), .R (RST)) ;
    mux21_ni ix7219 (.Y (nx7218), .A0 (Q[238]), .A1 (D[238]), .S0 (nx10235)) ;
    dffr reg_Q_239 (.Q (Q[239]), .QB (\$dummy [239]), .D (nx7228), .CLK (nx10113
         ), .R (RST)) ;
    mux21_ni ix7229 (.Y (nx7228), .A0 (Q[239]), .A1 (D[239]), .S0 (nx10235)) ;
    dffr reg_Q_240 (.Q (Q[240]), .QB (\$dummy [240]), .D (nx7238), .CLK (nx10113
         ), .R (RST)) ;
    mux21_ni ix7239 (.Y (nx7238), .A0 (Q[240]), .A1 (D[240]), .S0 (nx10235)) ;
    dffr reg_Q_241 (.Q (Q[241]), .QB (\$dummy [241]), .D (nx7248), .CLK (nx10113
         ), .R (RST)) ;
    mux21_ni ix7249 (.Y (nx7248), .A0 (Q[241]), .A1 (D[241]), .S0 (nx10235)) ;
    dffr reg_Q_242 (.Q (Q[242]), .QB (\$dummy [242]), .D (nx7258), .CLK (nx10113
         ), .R (RST)) ;
    mux21_ni ix7259 (.Y (nx7258), .A0 (Q[242]), .A1 (D[242]), .S0 (nx10235)) ;
    dffr reg_Q_243 (.Q (Q[243]), .QB (\$dummy [243]), .D (nx7268), .CLK (nx10113
         ), .R (RST)) ;
    mux21_ni ix7269 (.Y (nx7268), .A0 (Q[243]), .A1 (D[243]), .S0 (nx10235)) ;
    dffr reg_Q_244 (.Q (Q[244]), .QB (\$dummy [244]), .D (nx7278), .CLK (nx10113
         ), .R (RST)) ;
    mux21_ni ix7279 (.Y (nx7278), .A0 (Q[244]), .A1 (D[244]), .S0 (nx10235)) ;
    dffr reg_Q_245 (.Q (Q[245]), .QB (\$dummy [245]), .D (nx7288), .CLK (nx10115
         ), .R (RST)) ;
    mux21_ni ix7289 (.Y (nx7288), .A0 (Q[245]), .A1 (D[245]), .S0 (nx10237)) ;
    dffr reg_Q_246 (.Q (Q[246]), .QB (\$dummy [246]), .D (nx7298), .CLK (nx10115
         ), .R (RST)) ;
    mux21_ni ix7299 (.Y (nx7298), .A0 (Q[246]), .A1 (D[246]), .S0 (nx10237)) ;
    dffr reg_Q_247 (.Q (Q[247]), .QB (\$dummy [247]), .D (nx7308), .CLK (nx10115
         ), .R (RST)) ;
    mux21_ni ix7309 (.Y (nx7308), .A0 (Q[247]), .A1 (D[247]), .S0 (nx10237)) ;
    dffr reg_Q_248 (.Q (Q[248]), .QB (\$dummy [248]), .D (nx7318), .CLK (nx10115
         ), .R (RST)) ;
    mux21_ni ix7319 (.Y (nx7318), .A0 (Q[248]), .A1 (D[248]), .S0 (nx10237)) ;
    dffr reg_Q_249 (.Q (Q[249]), .QB (\$dummy [249]), .D (nx7328), .CLK (nx10115
         ), .R (RST)) ;
    mux21_ni ix7329 (.Y (nx7328), .A0 (Q[249]), .A1 (D[249]), .S0 (nx10237)) ;
    dffr reg_Q_250 (.Q (Q[250]), .QB (\$dummy [250]), .D (nx7338), .CLK (nx10115
         ), .R (RST)) ;
    mux21_ni ix7339 (.Y (nx7338), .A0 (Q[250]), .A1 (D[250]), .S0 (nx10237)) ;
    dffr reg_Q_251 (.Q (Q[251]), .QB (\$dummy [251]), .D (nx7348), .CLK (nx10115
         ), .R (RST)) ;
    mux21_ni ix7349 (.Y (nx7348), .A0 (Q[251]), .A1 (D[251]), .S0 (nx10237)) ;
    dffr reg_Q_252 (.Q (Q[252]), .QB (\$dummy [252]), .D (nx7358), .CLK (nx10117
         ), .R (RST)) ;
    mux21_ni ix7359 (.Y (nx7358), .A0 (Q[252]), .A1 (D[252]), .S0 (nx10239)) ;
    dffr reg_Q_253 (.Q (Q[253]), .QB (\$dummy [253]), .D (nx7368), .CLK (nx10117
         ), .R (RST)) ;
    mux21_ni ix7369 (.Y (nx7368), .A0 (Q[253]), .A1 (D[253]), .S0 (nx10239)) ;
    dffr reg_Q_254 (.Q (Q[254]), .QB (\$dummy [254]), .D (nx7378), .CLK (nx10117
         ), .R (RST)) ;
    mux21_ni ix7379 (.Y (nx7378), .A0 (Q[254]), .A1 (D[254]), .S0 (nx10239)) ;
    dffr reg_Q_255 (.Q (Q[255]), .QB (\$dummy [255]), .D (nx7388), .CLK (nx10117
         ), .R (RST)) ;
    mux21_ni ix7389 (.Y (nx7388), .A0 (Q[255]), .A1 (D[255]), .S0 (nx10239)) ;
    dffr reg_Q_256 (.Q (Q[256]), .QB (\$dummy [256]), .D (nx7398), .CLK (nx10117
         ), .R (RST)) ;
    mux21_ni ix7399 (.Y (nx7398), .A0 (Q[256]), .A1 (D[256]), .S0 (nx10239)) ;
    dffr reg_Q_257 (.Q (Q[257]), .QB (\$dummy [257]), .D (nx7408), .CLK (nx10117
         ), .R (RST)) ;
    mux21_ni ix7409 (.Y (nx7408), .A0 (Q[257]), .A1 (D[257]), .S0 (nx10239)) ;
    dffr reg_Q_258 (.Q (Q[258]), .QB (\$dummy [258]), .D (nx7418), .CLK (nx10117
         ), .R (RST)) ;
    mux21_ni ix7419 (.Y (nx7418), .A0 (Q[258]), .A1 (D[258]), .S0 (nx10239)) ;
    dffr reg_Q_259 (.Q (Q[259]), .QB (\$dummy [259]), .D (nx7428), .CLK (nx10119
         ), .R (RST)) ;
    mux21_ni ix7429 (.Y (nx7428), .A0 (Q[259]), .A1 (D[259]), .S0 (nx10241)) ;
    dffr reg_Q_260 (.Q (Q[260]), .QB (\$dummy [260]), .D (nx7438), .CLK (nx10119
         ), .R (RST)) ;
    mux21_ni ix7439 (.Y (nx7438), .A0 (Q[260]), .A1 (D[260]), .S0 (nx10241)) ;
    dffr reg_Q_261 (.Q (Q[261]), .QB (\$dummy [261]), .D (nx7448), .CLK (nx10119
         ), .R (RST)) ;
    mux21_ni ix7449 (.Y (nx7448), .A0 (Q[261]), .A1 (D[261]), .S0 (nx10241)) ;
    dffr reg_Q_262 (.Q (Q[262]), .QB (\$dummy [262]), .D (nx7458), .CLK (nx10119
         ), .R (RST)) ;
    mux21_ni ix7459 (.Y (nx7458), .A0 (Q[262]), .A1 (D[262]), .S0 (nx10241)) ;
    dffr reg_Q_263 (.Q (Q[263]), .QB (\$dummy [263]), .D (nx7468), .CLK (nx10119
         ), .R (RST)) ;
    mux21_ni ix7469 (.Y (nx7468), .A0 (Q[263]), .A1 (D[263]), .S0 (nx10241)) ;
    dffr reg_Q_264 (.Q (Q[264]), .QB (\$dummy [264]), .D (nx7478), .CLK (nx10119
         ), .R (RST)) ;
    mux21_ni ix7479 (.Y (nx7478), .A0 (Q[264]), .A1 (D[264]), .S0 (nx10241)) ;
    dffr reg_Q_265 (.Q (Q[265]), .QB (\$dummy [265]), .D (nx7488), .CLK (nx10119
         ), .R (RST)) ;
    mux21_ni ix7489 (.Y (nx7488), .A0 (Q[265]), .A1 (D[265]), .S0 (nx10241)) ;
    dffr reg_Q_266 (.Q (Q[266]), .QB (\$dummy [266]), .D (nx7498), .CLK (nx10121
         ), .R (RST)) ;
    mux21_ni ix7499 (.Y (nx7498), .A0 (Q[266]), .A1 (D[266]), .S0 (nx10243)) ;
    dffr reg_Q_267 (.Q (Q[267]), .QB (\$dummy [267]), .D (nx7508), .CLK (nx10121
         ), .R (RST)) ;
    mux21_ni ix7509 (.Y (nx7508), .A0 (Q[267]), .A1 (D[267]), .S0 (nx10243)) ;
    dffr reg_Q_268 (.Q (Q[268]), .QB (\$dummy [268]), .D (nx7518), .CLK (nx10121
         ), .R (RST)) ;
    mux21_ni ix7519 (.Y (nx7518), .A0 (Q[268]), .A1 (D[268]), .S0 (nx10243)) ;
    dffr reg_Q_269 (.Q (Q[269]), .QB (\$dummy [269]), .D (nx7528), .CLK (nx10121
         ), .R (RST)) ;
    mux21_ni ix7529 (.Y (nx7528), .A0 (Q[269]), .A1 (D[269]), .S0 (nx10243)) ;
    dffr reg_Q_270 (.Q (Q[270]), .QB (\$dummy [270]), .D (nx7538), .CLK (nx10121
         ), .R (RST)) ;
    mux21_ni ix7539 (.Y (nx7538), .A0 (Q[270]), .A1 (D[270]), .S0 (nx10243)) ;
    dffr reg_Q_271 (.Q (Q[271]), .QB (\$dummy [271]), .D (nx7548), .CLK (nx10121
         ), .R (RST)) ;
    mux21_ni ix7549 (.Y (nx7548), .A0 (Q[271]), .A1 (D[271]), .S0 (nx10243)) ;
    dffr reg_Q_272 (.Q (Q[272]), .QB (\$dummy [272]), .D (nx7558), .CLK (nx10121
         ), .R (RST)) ;
    mux21_ni ix7559 (.Y (nx7558), .A0 (Q[272]), .A1 (D[272]), .S0 (nx10243)) ;
    dffr reg_Q_273 (.Q (Q[273]), .QB (\$dummy [273]), .D (nx7568), .CLK (nx10123
         ), .R (RST)) ;
    mux21_ni ix7569 (.Y (nx7568), .A0 (Q[273]), .A1 (D[273]), .S0 (nx10245)) ;
    dffr reg_Q_274 (.Q (Q[274]), .QB (\$dummy [274]), .D (nx7578), .CLK (nx10123
         ), .R (RST)) ;
    mux21_ni ix7579 (.Y (nx7578), .A0 (Q[274]), .A1 (D[274]), .S0 (nx10245)) ;
    dffr reg_Q_275 (.Q (Q[275]), .QB (\$dummy [275]), .D (nx7588), .CLK (nx10123
         ), .R (RST)) ;
    mux21_ni ix7589 (.Y (nx7588), .A0 (Q[275]), .A1 (D[275]), .S0 (nx10245)) ;
    dffr reg_Q_276 (.Q (Q[276]), .QB (\$dummy [276]), .D (nx7598), .CLK (nx10123
         ), .R (RST)) ;
    mux21_ni ix7599 (.Y (nx7598), .A0 (Q[276]), .A1 (D[276]), .S0 (nx10245)) ;
    dffr reg_Q_277 (.Q (Q[277]), .QB (\$dummy [277]), .D (nx7608), .CLK (nx10123
         ), .R (RST)) ;
    mux21_ni ix7609 (.Y (nx7608), .A0 (Q[277]), .A1 (D[277]), .S0 (nx10245)) ;
    dffr reg_Q_278 (.Q (Q[278]), .QB (\$dummy [278]), .D (nx7618), .CLK (nx10123
         ), .R (RST)) ;
    mux21_ni ix7619 (.Y (nx7618), .A0 (Q[278]), .A1 (D[278]), .S0 (nx10245)) ;
    dffr reg_Q_279 (.Q (Q[279]), .QB (\$dummy [279]), .D (nx7628), .CLK (nx10123
         ), .R (RST)) ;
    mux21_ni ix7629 (.Y (nx7628), .A0 (Q[279]), .A1 (D[279]), .S0 (nx10245)) ;
    dffr reg_Q_280 (.Q (Q[280]), .QB (\$dummy [280]), .D (nx7638), .CLK (nx10125
         ), .R (RST)) ;
    mux21_ni ix7639 (.Y (nx7638), .A0 (Q[280]), .A1 (D[280]), .S0 (nx10247)) ;
    dffr reg_Q_281 (.Q (Q[281]), .QB (\$dummy [281]), .D (nx7648), .CLK (nx10125
         ), .R (RST)) ;
    mux21_ni ix7649 (.Y (nx7648), .A0 (Q[281]), .A1 (D[281]), .S0 (nx10247)) ;
    dffr reg_Q_282 (.Q (Q[282]), .QB (\$dummy [282]), .D (nx7658), .CLK (nx10125
         ), .R (RST)) ;
    mux21_ni ix7659 (.Y (nx7658), .A0 (Q[282]), .A1 (D[282]), .S0 (nx10247)) ;
    dffr reg_Q_283 (.Q (Q[283]), .QB (\$dummy [283]), .D (nx7668), .CLK (nx10125
         ), .R (RST)) ;
    mux21_ni ix7669 (.Y (nx7668), .A0 (Q[283]), .A1 (D[283]), .S0 (nx10247)) ;
    dffr reg_Q_284 (.Q (Q[284]), .QB (\$dummy [284]), .D (nx7678), .CLK (nx10125
         ), .R (RST)) ;
    mux21_ni ix7679 (.Y (nx7678), .A0 (Q[284]), .A1 (D[284]), .S0 (nx10247)) ;
    dffr reg_Q_285 (.Q (Q[285]), .QB (\$dummy [285]), .D (nx7688), .CLK (nx10125
         ), .R (RST)) ;
    mux21_ni ix7689 (.Y (nx7688), .A0 (Q[285]), .A1 (D[285]), .S0 (nx10247)) ;
    dffr reg_Q_286 (.Q (Q[286]), .QB (\$dummy [286]), .D (nx7698), .CLK (nx10125
         ), .R (RST)) ;
    mux21_ni ix7699 (.Y (nx7698), .A0 (Q[286]), .A1 (D[286]), .S0 (nx10247)) ;
    dffr reg_Q_287 (.Q (Q[287]), .QB (\$dummy [287]), .D (nx7708), .CLK (nx10127
         ), .R (RST)) ;
    mux21_ni ix7709 (.Y (nx7708), .A0 (Q[287]), .A1 (D[287]), .S0 (nx10249)) ;
    dffr reg_Q_288 (.Q (Q[288]), .QB (\$dummy [288]), .D (nx7718), .CLK (nx10127
         ), .R (RST)) ;
    mux21_ni ix7719 (.Y (nx7718), .A0 (Q[288]), .A1 (D[288]), .S0 (nx10249)) ;
    dffr reg_Q_289 (.Q (Q[289]), .QB (\$dummy [289]), .D (nx7728), .CLK (nx10127
         ), .R (RST)) ;
    mux21_ni ix7729 (.Y (nx7728), .A0 (Q[289]), .A1 (D[289]), .S0 (nx10249)) ;
    dffr reg_Q_290 (.Q (Q[290]), .QB (\$dummy [290]), .D (nx7738), .CLK (nx10127
         ), .R (RST)) ;
    mux21_ni ix7739 (.Y (nx7738), .A0 (Q[290]), .A1 (D[290]), .S0 (nx10249)) ;
    dffr reg_Q_291 (.Q (Q[291]), .QB (\$dummy [291]), .D (nx7748), .CLK (nx10127
         ), .R (RST)) ;
    mux21_ni ix7749 (.Y (nx7748), .A0 (Q[291]), .A1 (D[291]), .S0 (nx10249)) ;
    dffr reg_Q_292 (.Q (Q[292]), .QB (\$dummy [292]), .D (nx7758), .CLK (nx10127
         ), .R (RST)) ;
    mux21_ni ix7759 (.Y (nx7758), .A0 (Q[292]), .A1 (D[292]), .S0 (nx10249)) ;
    dffr reg_Q_293 (.Q (Q[293]), .QB (\$dummy [293]), .D (nx7768), .CLK (nx10127
         ), .R (RST)) ;
    mux21_ni ix7769 (.Y (nx7768), .A0 (Q[293]), .A1 (D[293]), .S0 (nx10249)) ;
    dffr reg_Q_294 (.Q (Q[294]), .QB (\$dummy [294]), .D (nx7778), .CLK (nx10129
         ), .R (RST)) ;
    mux21_ni ix7779 (.Y (nx7778), .A0 (Q[294]), .A1 (D[294]), .S0 (nx10251)) ;
    dffr reg_Q_295 (.Q (Q[295]), .QB (\$dummy [295]), .D (nx7788), .CLK (nx10129
         ), .R (RST)) ;
    mux21_ni ix7789 (.Y (nx7788), .A0 (Q[295]), .A1 (D[295]), .S0 (nx10251)) ;
    dffr reg_Q_296 (.Q (Q[296]), .QB (\$dummy [296]), .D (nx7798), .CLK (nx10129
         ), .R (RST)) ;
    mux21_ni ix7799 (.Y (nx7798), .A0 (Q[296]), .A1 (D[296]), .S0 (nx10251)) ;
    dffr reg_Q_297 (.Q (Q[297]), .QB (\$dummy [297]), .D (nx7808), .CLK (nx10129
         ), .R (RST)) ;
    mux21_ni ix7809 (.Y (nx7808), .A0 (Q[297]), .A1 (D[297]), .S0 (nx10251)) ;
    dffr reg_Q_298 (.Q (Q[298]), .QB (\$dummy [298]), .D (nx7818), .CLK (nx10129
         ), .R (RST)) ;
    mux21_ni ix7819 (.Y (nx7818), .A0 (Q[298]), .A1 (D[298]), .S0 (nx10251)) ;
    dffr reg_Q_299 (.Q (Q[299]), .QB (\$dummy [299]), .D (nx7828), .CLK (nx10129
         ), .R (RST)) ;
    mux21_ni ix7829 (.Y (nx7828), .A0 (Q[299]), .A1 (D[299]), .S0 (nx10251)) ;
    dffr reg_Q_300 (.Q (Q[300]), .QB (\$dummy [300]), .D (nx7838), .CLK (nx10129
         ), .R (RST)) ;
    mux21_ni ix7839 (.Y (nx7838), .A0 (Q[300]), .A1 (D[300]), .S0 (nx10251)) ;
    dffr reg_Q_301 (.Q (Q[301]), .QB (\$dummy [301]), .D (nx7848), .CLK (nx10131
         ), .R (RST)) ;
    mux21_ni ix7849 (.Y (nx7848), .A0 (Q[301]), .A1 (D[301]), .S0 (nx10253)) ;
    dffr reg_Q_302 (.Q (Q[302]), .QB (\$dummy [302]), .D (nx7858), .CLK (nx10131
         ), .R (RST)) ;
    mux21_ni ix7859 (.Y (nx7858), .A0 (Q[302]), .A1 (D[302]), .S0 (nx10253)) ;
    dffr reg_Q_303 (.Q (Q[303]), .QB (\$dummy [303]), .D (nx7868), .CLK (nx10131
         ), .R (RST)) ;
    mux21_ni ix7869 (.Y (nx7868), .A0 (Q[303]), .A1 (D[303]), .S0 (nx10253)) ;
    dffr reg_Q_304 (.Q (Q[304]), .QB (\$dummy [304]), .D (nx7878), .CLK (nx10131
         ), .R (RST)) ;
    mux21_ni ix7879 (.Y (nx7878), .A0 (Q[304]), .A1 (D[304]), .S0 (nx10253)) ;
    dffr reg_Q_305 (.Q (Q[305]), .QB (\$dummy [305]), .D (nx7888), .CLK (nx10131
         ), .R (RST)) ;
    mux21_ni ix7889 (.Y (nx7888), .A0 (Q[305]), .A1 (D[305]), .S0 (nx10253)) ;
    dffr reg_Q_306 (.Q (Q[306]), .QB (\$dummy [306]), .D (nx7898), .CLK (nx10131
         ), .R (RST)) ;
    mux21_ni ix7899 (.Y (nx7898), .A0 (Q[306]), .A1 (D[306]), .S0 (nx10253)) ;
    dffr reg_Q_307 (.Q (Q[307]), .QB (\$dummy [307]), .D (nx7908), .CLK (nx10131
         ), .R (RST)) ;
    mux21_ni ix7909 (.Y (nx7908), .A0 (Q[307]), .A1 (D[307]), .S0 (nx10253)) ;
    dffr reg_Q_308 (.Q (Q[308]), .QB (\$dummy [308]), .D (nx7918), .CLK (nx10133
         ), .R (RST)) ;
    mux21_ni ix7919 (.Y (nx7918), .A0 (Q[308]), .A1 (D[308]), .S0 (nx10255)) ;
    dffr reg_Q_309 (.Q (Q[309]), .QB (\$dummy [309]), .D (nx7928), .CLK (nx10133
         ), .R (RST)) ;
    mux21_ni ix7929 (.Y (nx7928), .A0 (Q[309]), .A1 (D[309]), .S0 (nx10255)) ;
    dffr reg_Q_310 (.Q (Q[310]), .QB (\$dummy [310]), .D (nx7938), .CLK (nx10133
         ), .R (RST)) ;
    mux21_ni ix7939 (.Y (nx7938), .A0 (Q[310]), .A1 (D[310]), .S0 (nx10255)) ;
    dffr reg_Q_311 (.Q (Q[311]), .QB (\$dummy [311]), .D (nx7948), .CLK (nx10133
         ), .R (RST)) ;
    mux21_ni ix7949 (.Y (nx7948), .A0 (Q[311]), .A1 (D[311]), .S0 (nx10255)) ;
    dffr reg_Q_312 (.Q (Q[312]), .QB (\$dummy [312]), .D (nx7958), .CLK (nx10133
         ), .R (RST)) ;
    mux21_ni ix7959 (.Y (nx7958), .A0 (Q[312]), .A1 (D[312]), .S0 (nx10255)) ;
    dffr reg_Q_313 (.Q (Q[313]), .QB (\$dummy [313]), .D (nx7968), .CLK (nx10133
         ), .R (RST)) ;
    mux21_ni ix7969 (.Y (nx7968), .A0 (Q[313]), .A1 (D[313]), .S0 (nx10255)) ;
    dffr reg_Q_314 (.Q (Q[314]), .QB (\$dummy [314]), .D (nx7978), .CLK (nx10133
         ), .R (RST)) ;
    mux21_ni ix7979 (.Y (nx7978), .A0 (Q[314]), .A1 (D[314]), .S0 (nx10255)) ;
    dffr reg_Q_315 (.Q (Q[315]), .QB (\$dummy [315]), .D (nx7988), .CLK (nx10135
         ), .R (RST)) ;
    mux21_ni ix7989 (.Y (nx7988), .A0 (Q[315]), .A1 (D[315]), .S0 (nx10257)) ;
    dffr reg_Q_316 (.Q (Q[316]), .QB (\$dummy [316]), .D (nx7998), .CLK (nx10135
         ), .R (RST)) ;
    mux21_ni ix7999 (.Y (nx7998), .A0 (Q[316]), .A1 (D[316]), .S0 (nx10257)) ;
    dffr reg_Q_317 (.Q (Q[317]), .QB (\$dummy [317]), .D (nx8008), .CLK (nx10135
         ), .R (RST)) ;
    mux21_ni ix8009 (.Y (nx8008), .A0 (Q[317]), .A1 (D[317]), .S0 (nx10257)) ;
    dffr reg_Q_318 (.Q (Q[318]), .QB (\$dummy [318]), .D (nx8018), .CLK (nx10135
         ), .R (RST)) ;
    mux21_ni ix8019 (.Y (nx8018), .A0 (Q[318]), .A1 (D[318]), .S0 (nx10257)) ;
    dffr reg_Q_319 (.Q (Q[319]), .QB (\$dummy [319]), .D (nx8028), .CLK (nx10135
         ), .R (RST)) ;
    mux21_ni ix8029 (.Y (nx8028), .A0 (Q[319]), .A1 (D[319]), .S0 (nx10257)) ;
    dffr reg_Q_320 (.Q (Q[320]), .QB (\$dummy [320]), .D (nx8038), .CLK (nx10135
         ), .R (RST)) ;
    mux21_ni ix8039 (.Y (nx8038), .A0 (Q[320]), .A1 (D[320]), .S0 (nx10257)) ;
    dffr reg_Q_321 (.Q (Q[321]), .QB (\$dummy [321]), .D (nx8048), .CLK (nx10135
         ), .R (RST)) ;
    mux21_ni ix8049 (.Y (nx8048), .A0 (Q[321]), .A1 (D[321]), .S0 (nx10257)) ;
    dffr reg_Q_322 (.Q (Q[322]), .QB (\$dummy [322]), .D (nx8058), .CLK (nx10137
         ), .R (RST)) ;
    mux21_ni ix8059 (.Y (nx8058), .A0 (Q[322]), .A1 (D[322]), .S0 (nx10259)) ;
    dffr reg_Q_323 (.Q (Q[323]), .QB (\$dummy [323]), .D (nx8068), .CLK (nx10137
         ), .R (RST)) ;
    mux21_ni ix8069 (.Y (nx8068), .A0 (Q[323]), .A1 (D[323]), .S0 (nx10259)) ;
    dffr reg_Q_324 (.Q (Q[324]), .QB (\$dummy [324]), .D (nx8078), .CLK (nx10137
         ), .R (RST)) ;
    mux21_ni ix8079 (.Y (nx8078), .A0 (Q[324]), .A1 (D[324]), .S0 (nx10259)) ;
    dffr reg_Q_325 (.Q (Q[325]), .QB (\$dummy [325]), .D (nx8088), .CLK (nx10137
         ), .R (RST)) ;
    mux21_ni ix8089 (.Y (nx8088), .A0 (Q[325]), .A1 (D[325]), .S0 (nx10259)) ;
    dffr reg_Q_326 (.Q (Q[326]), .QB (\$dummy [326]), .D (nx8098), .CLK (nx10137
         ), .R (RST)) ;
    mux21_ni ix8099 (.Y (nx8098), .A0 (Q[326]), .A1 (D[326]), .S0 (nx10259)) ;
    dffr reg_Q_327 (.Q (Q[327]), .QB (\$dummy [327]), .D (nx8108), .CLK (nx10137
         ), .R (RST)) ;
    mux21_ni ix8109 (.Y (nx8108), .A0 (Q[327]), .A1 (D[327]), .S0 (nx10259)) ;
    dffr reg_Q_328 (.Q (Q[328]), .QB (\$dummy [328]), .D (nx8118), .CLK (nx10137
         ), .R (RST)) ;
    mux21_ni ix8119 (.Y (nx8118), .A0 (Q[328]), .A1 (D[328]), .S0 (nx10259)) ;
    dffr reg_Q_329 (.Q (Q[329]), .QB (\$dummy [329]), .D (nx8128), .CLK (nx10139
         ), .R (RST)) ;
    mux21_ni ix8129 (.Y (nx8128), .A0 (Q[329]), .A1 (D[329]), .S0 (nx10261)) ;
    dffr reg_Q_330 (.Q (Q[330]), .QB (\$dummy [330]), .D (nx8138), .CLK (nx10139
         ), .R (RST)) ;
    mux21_ni ix8139 (.Y (nx8138), .A0 (Q[330]), .A1 (D[330]), .S0 (nx10261)) ;
    dffr reg_Q_331 (.Q (Q[331]), .QB (\$dummy [331]), .D (nx8148), .CLK (nx10139
         ), .R (RST)) ;
    mux21_ni ix8149 (.Y (nx8148), .A0 (Q[331]), .A1 (D[331]), .S0 (nx10261)) ;
    dffr reg_Q_332 (.Q (Q[332]), .QB (\$dummy [332]), .D (nx8158), .CLK (nx10139
         ), .R (RST)) ;
    mux21_ni ix8159 (.Y (nx8158), .A0 (Q[332]), .A1 (D[332]), .S0 (nx10261)) ;
    dffr reg_Q_333 (.Q (Q[333]), .QB (\$dummy [333]), .D (nx8168), .CLK (nx10139
         ), .R (RST)) ;
    mux21_ni ix8169 (.Y (nx8168), .A0 (Q[333]), .A1 (D[333]), .S0 (nx10261)) ;
    dffr reg_Q_334 (.Q (Q[334]), .QB (\$dummy [334]), .D (nx8178), .CLK (nx10139
         ), .R (RST)) ;
    mux21_ni ix8179 (.Y (nx8178), .A0 (Q[334]), .A1 (D[334]), .S0 (nx10261)) ;
    dffr reg_Q_335 (.Q (Q[335]), .QB (\$dummy [335]), .D (nx8188), .CLK (nx10139
         ), .R (RST)) ;
    mux21_ni ix8189 (.Y (nx8188), .A0 (Q[335]), .A1 (D[335]), .S0 (nx10261)) ;
    dffr reg_Q_336 (.Q (Q[336]), .QB (\$dummy [336]), .D (nx8198), .CLK (nx10141
         ), .R (RST)) ;
    mux21_ni ix8199 (.Y (nx8198), .A0 (Q[336]), .A1 (D[336]), .S0 (nx10263)) ;
    dffr reg_Q_337 (.Q (Q[337]), .QB (\$dummy [337]), .D (nx8208), .CLK (nx10141
         ), .R (RST)) ;
    mux21_ni ix8209 (.Y (nx8208), .A0 (Q[337]), .A1 (D[337]), .S0 (nx10263)) ;
    dffr reg_Q_338 (.Q (Q[338]), .QB (\$dummy [338]), .D (nx8218), .CLK (nx10141
         ), .R (RST)) ;
    mux21_ni ix8219 (.Y (nx8218), .A0 (Q[338]), .A1 (D[338]), .S0 (nx10263)) ;
    dffr reg_Q_339 (.Q (Q[339]), .QB (\$dummy [339]), .D (nx8228), .CLK (nx10141
         ), .R (RST)) ;
    mux21_ni ix8229 (.Y (nx8228), .A0 (Q[339]), .A1 (D[339]), .S0 (nx10263)) ;
    dffr reg_Q_340 (.Q (Q[340]), .QB (\$dummy [340]), .D (nx8238), .CLK (nx10141
         ), .R (RST)) ;
    mux21_ni ix8239 (.Y (nx8238), .A0 (Q[340]), .A1 (D[340]), .S0 (nx10263)) ;
    dffr reg_Q_341 (.Q (Q[341]), .QB (\$dummy [341]), .D (nx8248), .CLK (nx10141
         ), .R (RST)) ;
    mux21_ni ix8249 (.Y (nx8248), .A0 (Q[341]), .A1 (D[341]), .S0 (nx10263)) ;
    dffr reg_Q_342 (.Q (Q[342]), .QB (\$dummy [342]), .D (nx8258), .CLK (nx10141
         ), .R (RST)) ;
    mux21_ni ix8259 (.Y (nx8258), .A0 (Q[342]), .A1 (D[342]), .S0 (nx10263)) ;
    dffr reg_Q_343 (.Q (Q[343]), .QB (\$dummy [343]), .D (nx8268), .CLK (nx10143
         ), .R (RST)) ;
    mux21_ni ix8269 (.Y (nx8268), .A0 (Q[343]), .A1 (D[343]), .S0 (nx10265)) ;
    dffr reg_Q_344 (.Q (Q[344]), .QB (\$dummy [344]), .D (nx8278), .CLK (nx10143
         ), .R (RST)) ;
    mux21_ni ix8279 (.Y (nx8278), .A0 (Q[344]), .A1 (D[344]), .S0 (nx10265)) ;
    dffr reg_Q_345 (.Q (Q[345]), .QB (\$dummy [345]), .D (nx8288), .CLK (nx10143
         ), .R (RST)) ;
    mux21_ni ix8289 (.Y (nx8288), .A0 (Q[345]), .A1 (D[345]), .S0 (nx10265)) ;
    dffr reg_Q_346 (.Q (Q[346]), .QB (\$dummy [346]), .D (nx8298), .CLK (nx10143
         ), .R (RST)) ;
    mux21_ni ix8299 (.Y (nx8298), .A0 (Q[346]), .A1 (D[346]), .S0 (nx10265)) ;
    dffr reg_Q_347 (.Q (Q[347]), .QB (\$dummy [347]), .D (nx8308), .CLK (nx10143
         ), .R (RST)) ;
    mux21_ni ix8309 (.Y (nx8308), .A0 (Q[347]), .A1 (D[347]), .S0 (nx10265)) ;
    dffr reg_Q_348 (.Q (Q[348]), .QB (\$dummy [348]), .D (nx8318), .CLK (nx10143
         ), .R (RST)) ;
    mux21_ni ix8319 (.Y (nx8318), .A0 (Q[348]), .A1 (D[348]), .S0 (nx10265)) ;
    dffr reg_Q_349 (.Q (Q[349]), .QB (\$dummy [349]), .D (nx8328), .CLK (nx10143
         ), .R (RST)) ;
    mux21_ni ix8329 (.Y (nx8328), .A0 (Q[349]), .A1 (D[349]), .S0 (nx10265)) ;
    dffr reg_Q_350 (.Q (Q[350]), .QB (\$dummy [350]), .D (nx8338), .CLK (nx10145
         ), .R (RST)) ;
    mux21_ni ix8339 (.Y (nx8338), .A0 (Q[350]), .A1 (D[350]), .S0 (nx10267)) ;
    dffr reg_Q_351 (.Q (Q[351]), .QB (\$dummy [351]), .D (nx8348), .CLK (nx10145
         ), .R (RST)) ;
    mux21_ni ix8349 (.Y (nx8348), .A0 (Q[351]), .A1 (D[351]), .S0 (nx10267)) ;
    dffr reg_Q_352 (.Q (Q[352]), .QB (\$dummy [352]), .D (nx8358), .CLK (nx10145
         ), .R (RST)) ;
    mux21_ni ix8359 (.Y (nx8358), .A0 (Q[352]), .A1 (D[352]), .S0 (nx10267)) ;
    dffr reg_Q_353 (.Q (Q[353]), .QB (\$dummy [353]), .D (nx8368), .CLK (nx10145
         ), .R (RST)) ;
    mux21_ni ix8369 (.Y (nx8368), .A0 (Q[353]), .A1 (D[353]), .S0 (nx10267)) ;
    dffr reg_Q_354 (.Q (Q[354]), .QB (\$dummy [354]), .D (nx8378), .CLK (nx10145
         ), .R (RST)) ;
    mux21_ni ix8379 (.Y (nx8378), .A0 (Q[354]), .A1 (D[354]), .S0 (nx10267)) ;
    dffr reg_Q_355 (.Q (Q[355]), .QB (\$dummy [355]), .D (nx8388), .CLK (nx10145
         ), .R (RST)) ;
    mux21_ni ix8389 (.Y (nx8388), .A0 (Q[355]), .A1 (D[355]), .S0 (nx10267)) ;
    dffr reg_Q_356 (.Q (Q[356]), .QB (\$dummy [356]), .D (nx8398), .CLK (nx10145
         ), .R (RST)) ;
    mux21_ni ix8399 (.Y (nx8398), .A0 (Q[356]), .A1 (D[356]), .S0 (nx10267)) ;
    dffr reg_Q_357 (.Q (Q[357]), .QB (\$dummy [357]), .D (nx8408), .CLK (nx10147
         ), .R (RST)) ;
    mux21_ni ix8409 (.Y (nx8408), .A0 (Q[357]), .A1 (D[357]), .S0 (nx10269)) ;
    dffr reg_Q_358 (.Q (Q[358]), .QB (\$dummy [358]), .D (nx8418), .CLK (nx10147
         ), .R (RST)) ;
    mux21_ni ix8419 (.Y (nx8418), .A0 (Q[358]), .A1 (D[358]), .S0 (nx10269)) ;
    dffr reg_Q_359 (.Q (Q[359]), .QB (\$dummy [359]), .D (nx8428), .CLK (nx10147
         ), .R (RST)) ;
    mux21_ni ix8429 (.Y (nx8428), .A0 (Q[359]), .A1 (D[359]), .S0 (nx10269)) ;
    dffr reg_Q_360 (.Q (Q[360]), .QB (\$dummy [360]), .D (nx8438), .CLK (nx10147
         ), .R (RST)) ;
    mux21_ni ix8439 (.Y (nx8438), .A0 (Q[360]), .A1 (D[360]), .S0 (nx10269)) ;
    dffr reg_Q_361 (.Q (Q[361]), .QB (\$dummy [361]), .D (nx8448), .CLK (nx10147
         ), .R (RST)) ;
    mux21_ni ix8449 (.Y (nx8448), .A0 (Q[361]), .A1 (D[361]), .S0 (nx10269)) ;
    dffr reg_Q_362 (.Q (Q[362]), .QB (\$dummy [362]), .D (nx8458), .CLK (nx10147
         ), .R (RST)) ;
    mux21_ni ix8459 (.Y (nx8458), .A0 (Q[362]), .A1 (D[362]), .S0 (nx10269)) ;
    dffr reg_Q_363 (.Q (Q[363]), .QB (\$dummy [363]), .D (nx8468), .CLK (nx10147
         ), .R (RST)) ;
    mux21_ni ix8469 (.Y (nx8468), .A0 (Q[363]), .A1 (D[363]), .S0 (nx10269)) ;
    dffr reg_Q_364 (.Q (Q[364]), .QB (\$dummy [364]), .D (nx8478), .CLK (nx10149
         ), .R (RST)) ;
    mux21_ni ix8479 (.Y (nx8478), .A0 (Q[364]), .A1 (D[364]), .S0 (nx10271)) ;
    dffr reg_Q_365 (.Q (Q[365]), .QB (\$dummy [365]), .D (nx8488), .CLK (nx10149
         ), .R (RST)) ;
    mux21_ni ix8489 (.Y (nx8488), .A0 (Q[365]), .A1 (D[365]), .S0 (nx10271)) ;
    dffr reg_Q_366 (.Q (Q[366]), .QB (\$dummy [366]), .D (nx8498), .CLK (nx10149
         ), .R (RST)) ;
    mux21_ni ix8499 (.Y (nx8498), .A0 (Q[366]), .A1 (D[366]), .S0 (nx10271)) ;
    dffr reg_Q_367 (.Q (Q[367]), .QB (\$dummy [367]), .D (nx8508), .CLK (nx10149
         ), .R (RST)) ;
    mux21_ni ix8509 (.Y (nx8508), .A0 (Q[367]), .A1 (D[367]), .S0 (nx10271)) ;
    dffr reg_Q_368 (.Q (Q[368]), .QB (\$dummy [368]), .D (nx8518), .CLK (nx10149
         ), .R (RST)) ;
    mux21_ni ix8519 (.Y (nx8518), .A0 (Q[368]), .A1 (D[368]), .S0 (nx10271)) ;
    dffr reg_Q_369 (.Q (Q[369]), .QB (\$dummy [369]), .D (nx8528), .CLK (nx10149
         ), .R (RST)) ;
    mux21_ni ix8529 (.Y (nx8528), .A0 (Q[369]), .A1 (D[369]), .S0 (nx10271)) ;
    dffr reg_Q_370 (.Q (Q[370]), .QB (\$dummy [370]), .D (nx8538), .CLK (nx10149
         ), .R (RST)) ;
    mux21_ni ix8539 (.Y (nx8538), .A0 (Q[370]), .A1 (D[370]), .S0 (nx10271)) ;
    dffr reg_Q_371 (.Q (Q[371]), .QB (\$dummy [371]), .D (nx8548), .CLK (nx10151
         ), .R (RST)) ;
    mux21_ni ix8549 (.Y (nx8548), .A0 (Q[371]), .A1 (D[371]), .S0 (nx10273)) ;
    dffr reg_Q_372 (.Q (Q[372]), .QB (\$dummy [372]), .D (nx8558), .CLK (nx10151
         ), .R (RST)) ;
    mux21_ni ix8559 (.Y (nx8558), .A0 (Q[372]), .A1 (D[372]), .S0 (nx10273)) ;
    dffr reg_Q_373 (.Q (Q[373]), .QB (\$dummy [373]), .D (nx8568), .CLK (nx10151
         ), .R (RST)) ;
    mux21_ni ix8569 (.Y (nx8568), .A0 (Q[373]), .A1 (D[373]), .S0 (nx10273)) ;
    dffr reg_Q_374 (.Q (Q[374]), .QB (\$dummy [374]), .D (nx8578), .CLK (nx10151
         ), .R (RST)) ;
    mux21_ni ix8579 (.Y (nx8578), .A0 (Q[374]), .A1 (D[374]), .S0 (nx10273)) ;
    dffr reg_Q_375 (.Q (Q[375]), .QB (\$dummy [375]), .D (nx8588), .CLK (nx10151
         ), .R (RST)) ;
    mux21_ni ix8589 (.Y (nx8588), .A0 (Q[375]), .A1 (D[375]), .S0 (nx10273)) ;
    dffr reg_Q_376 (.Q (Q[376]), .QB (\$dummy [376]), .D (nx8598), .CLK (nx10151
         ), .R (RST)) ;
    mux21_ni ix8599 (.Y (nx8598), .A0 (Q[376]), .A1 (D[376]), .S0 (nx10273)) ;
    dffr reg_Q_377 (.Q (Q[377]), .QB (\$dummy [377]), .D (nx8608), .CLK (nx10151
         ), .R (RST)) ;
    mux21_ni ix8609 (.Y (nx8608), .A0 (Q[377]), .A1 (D[377]), .S0 (nx10273)) ;
    dffr reg_Q_378 (.Q (Q[378]), .QB (\$dummy [378]), .D (nx8618), .CLK (nx10153
         ), .R (RST)) ;
    mux21_ni ix8619 (.Y (nx8618), .A0 (Q[378]), .A1 (D[378]), .S0 (nx10275)) ;
    dffr reg_Q_379 (.Q (Q[379]), .QB (\$dummy [379]), .D (nx8628), .CLK (nx10153
         ), .R (RST)) ;
    mux21_ni ix8629 (.Y (nx8628), .A0 (Q[379]), .A1 (D[379]), .S0 (nx10275)) ;
    dffr reg_Q_380 (.Q (Q[380]), .QB (\$dummy [380]), .D (nx8638), .CLK (nx10153
         ), .R (RST)) ;
    mux21_ni ix8639 (.Y (nx8638), .A0 (Q[380]), .A1 (D[380]), .S0 (nx10275)) ;
    dffr reg_Q_381 (.Q (Q[381]), .QB (\$dummy [381]), .D (nx8648), .CLK (nx10153
         ), .R (RST)) ;
    mux21_ni ix8649 (.Y (nx8648), .A0 (Q[381]), .A1 (D[381]), .S0 (nx10275)) ;
    dffr reg_Q_382 (.Q (Q[382]), .QB (\$dummy [382]), .D (nx8658), .CLK (nx10153
         ), .R (RST)) ;
    mux21_ni ix8659 (.Y (nx8658), .A0 (Q[382]), .A1 (D[382]), .S0 (nx10275)) ;
    dffr reg_Q_383 (.Q (Q[383]), .QB (\$dummy [383]), .D (nx8668), .CLK (nx10153
         ), .R (RST)) ;
    mux21_ni ix8669 (.Y (nx8668), .A0 (Q[383]), .A1 (D[383]), .S0 (nx10275)) ;
    dffr reg_Q_384 (.Q (Q[384]), .QB (\$dummy [384]), .D (nx8678), .CLK (nx10153
         ), .R (RST)) ;
    mux21_ni ix8679 (.Y (nx8678), .A0 (Q[384]), .A1 (D[384]), .S0 (nx10275)) ;
    dffr reg_Q_385 (.Q (Q[385]), .QB (\$dummy [385]), .D (nx8688), .CLK (nx10155
         ), .R (RST)) ;
    mux21_ni ix8689 (.Y (nx8688), .A0 (Q[385]), .A1 (D[385]), .S0 (nx10277)) ;
    dffr reg_Q_386 (.Q (Q[386]), .QB (\$dummy [386]), .D (nx8698), .CLK (nx10155
         ), .R (RST)) ;
    mux21_ni ix8699 (.Y (nx8698), .A0 (Q[386]), .A1 (D[386]), .S0 (nx10277)) ;
    dffr reg_Q_387 (.Q (Q[387]), .QB (\$dummy [387]), .D (nx8708), .CLK (nx10155
         ), .R (RST)) ;
    mux21_ni ix8709 (.Y (nx8708), .A0 (Q[387]), .A1 (D[387]), .S0 (nx10277)) ;
    dffr reg_Q_388 (.Q (Q[388]), .QB (\$dummy [388]), .D (nx8718), .CLK (nx10155
         ), .R (RST)) ;
    mux21_ni ix8719 (.Y (nx8718), .A0 (Q[388]), .A1 (D[388]), .S0 (nx10277)) ;
    dffr reg_Q_389 (.Q (Q[389]), .QB (\$dummy [389]), .D (nx8728), .CLK (nx10155
         ), .R (RST)) ;
    mux21_ni ix8729 (.Y (nx8728), .A0 (Q[389]), .A1 (D[389]), .S0 (nx10277)) ;
    dffr reg_Q_390 (.Q (Q[390]), .QB (\$dummy [390]), .D (nx8738), .CLK (nx10155
         ), .R (RST)) ;
    mux21_ni ix8739 (.Y (nx8738), .A0 (Q[390]), .A1 (D[390]), .S0 (nx10277)) ;
    dffr reg_Q_391 (.Q (Q[391]), .QB (\$dummy [391]), .D (nx8748), .CLK (nx10155
         ), .R (RST)) ;
    mux21_ni ix8749 (.Y (nx8748), .A0 (Q[391]), .A1 (D[391]), .S0 (nx10277)) ;
    dffr reg_Q_392 (.Q (Q[392]), .QB (\$dummy [392]), .D (nx8758), .CLK (nx10157
         ), .R (RST)) ;
    mux21_ni ix8759 (.Y (nx8758), .A0 (Q[392]), .A1 (D[392]), .S0 (nx10279)) ;
    dffr reg_Q_393 (.Q (Q[393]), .QB (\$dummy [393]), .D (nx8768), .CLK (nx10157
         ), .R (RST)) ;
    mux21_ni ix8769 (.Y (nx8768), .A0 (Q[393]), .A1 (D[393]), .S0 (nx10279)) ;
    dffr reg_Q_394 (.Q (Q[394]), .QB (\$dummy [394]), .D (nx8778), .CLK (nx10157
         ), .R (RST)) ;
    mux21_ni ix8779 (.Y (nx8778), .A0 (Q[394]), .A1 (D[394]), .S0 (nx10279)) ;
    dffr reg_Q_395 (.Q (Q[395]), .QB (\$dummy [395]), .D (nx8788), .CLK (nx10157
         ), .R (RST)) ;
    mux21_ni ix8789 (.Y (nx8788), .A0 (Q[395]), .A1 (D[395]), .S0 (nx10279)) ;
    dffr reg_Q_396 (.Q (Q[396]), .QB (\$dummy [396]), .D (nx8798), .CLK (nx10157
         ), .R (RST)) ;
    mux21_ni ix8799 (.Y (nx8798), .A0 (Q[396]), .A1 (D[396]), .S0 (nx10279)) ;
    dffr reg_Q_397 (.Q (Q[397]), .QB (\$dummy [397]), .D (nx8808), .CLK (nx10157
         ), .R (RST)) ;
    mux21_ni ix8809 (.Y (nx8808), .A0 (Q[397]), .A1 (D[397]), .S0 (nx10279)) ;
    dffr reg_Q_398 (.Q (Q[398]), .QB (\$dummy [398]), .D (nx8818), .CLK (nx10157
         ), .R (RST)) ;
    mux21_ni ix8819 (.Y (nx8818), .A0 (Q[398]), .A1 (D[398]), .S0 (nx10279)) ;
    dffr reg_Q_399 (.Q (Q[399]), .QB (\$dummy [399]), .D (nx8828), .CLK (nx10159
         ), .R (RST)) ;
    mux21_ni ix8829 (.Y (nx8828), .A0 (Q[399]), .A1 (D[399]), .S0 (nx10281)) ;
    inv02 ix10044 (.Y (nx10045), .A (CLK)) ;
    inv02 ix10046 (.Y (nx10047), .A (nx10283)) ;
    inv02 ix10048 (.Y (nx10049), .A (nx10283)) ;
    inv02 ix10050 (.Y (nx10051), .A (nx10283)) ;
    inv02 ix10052 (.Y (nx10053), .A (nx10283)) ;
    inv02 ix10054 (.Y (nx10055), .A (nx10283)) ;
    inv02 ix10056 (.Y (nx10057), .A (nx10283)) ;
    inv02 ix10058 (.Y (nx10059), .A (nx10283)) ;
    inv02 ix10060 (.Y (nx10061), .A (nx10285)) ;
    inv02 ix10062 (.Y (nx10063), .A (nx10285)) ;
    inv02 ix10064 (.Y (nx10065), .A (nx10285)) ;
    inv02 ix10066 (.Y (nx10067), .A (nx10285)) ;
    inv02 ix10068 (.Y (nx10069), .A (nx10285)) ;
    inv02 ix10070 (.Y (nx10071), .A (nx10285)) ;
    inv02 ix10072 (.Y (nx10073), .A (nx10285)) ;
    inv02 ix10074 (.Y (nx10075), .A (nx10287)) ;
    inv02 ix10076 (.Y (nx10077), .A (nx10287)) ;
    inv02 ix10078 (.Y (nx10079), .A (nx10287)) ;
    inv02 ix10080 (.Y (nx10081), .A (nx10287)) ;
    inv02 ix10082 (.Y (nx10083), .A (nx10287)) ;
    inv02 ix10084 (.Y (nx10085), .A (nx10287)) ;
    inv02 ix10086 (.Y (nx10087), .A (nx10287)) ;
    inv02 ix10088 (.Y (nx10089), .A (nx10289)) ;
    inv02 ix10090 (.Y (nx10091), .A (nx10289)) ;
    inv02 ix10092 (.Y (nx10093), .A (nx10289)) ;
    inv02 ix10094 (.Y (nx10095), .A (nx10289)) ;
    inv02 ix10096 (.Y (nx10097), .A (nx10289)) ;
    inv02 ix10098 (.Y (nx10099), .A (nx10289)) ;
    inv02 ix10100 (.Y (nx10101), .A (nx10289)) ;
    inv02 ix10102 (.Y (nx10103), .A (nx10291)) ;
    inv02 ix10104 (.Y (nx10105), .A (nx10291)) ;
    inv02 ix10106 (.Y (nx10107), .A (nx10291)) ;
    inv02 ix10108 (.Y (nx10109), .A (nx10291)) ;
    inv02 ix10110 (.Y (nx10111), .A (nx10291)) ;
    inv02 ix10112 (.Y (nx10113), .A (nx10291)) ;
    inv02 ix10114 (.Y (nx10115), .A (nx10291)) ;
    inv02 ix10116 (.Y (nx10117), .A (nx10293)) ;
    inv02 ix10118 (.Y (nx10119), .A (nx10293)) ;
    inv02 ix10120 (.Y (nx10121), .A (nx10293)) ;
    inv02 ix10122 (.Y (nx10123), .A (nx10293)) ;
    inv02 ix10124 (.Y (nx10125), .A (nx10293)) ;
    inv02 ix10126 (.Y (nx10127), .A (nx10293)) ;
    inv02 ix10128 (.Y (nx10129), .A (nx10293)) ;
    inv02 ix10130 (.Y (nx10131), .A (nx10295)) ;
    inv02 ix10132 (.Y (nx10133), .A (nx10295)) ;
    inv02 ix10134 (.Y (nx10135), .A (nx10295)) ;
    inv02 ix10136 (.Y (nx10137), .A (nx10295)) ;
    inv02 ix10138 (.Y (nx10139), .A (nx10295)) ;
    inv02 ix10140 (.Y (nx10141), .A (nx10295)) ;
    inv02 ix10142 (.Y (nx10143), .A (nx10295)) ;
    inv02 ix10144 (.Y (nx10145), .A (nx10297)) ;
    inv02 ix10146 (.Y (nx10147), .A (nx10297)) ;
    inv02 ix10148 (.Y (nx10149), .A (nx10297)) ;
    inv02 ix10150 (.Y (nx10151), .A (nx10297)) ;
    inv02 ix10152 (.Y (nx10153), .A (nx10297)) ;
    inv02 ix10154 (.Y (nx10155), .A (nx10297)) ;
    inv02 ix10156 (.Y (nx10157), .A (nx10297)) ;
    inv02 ix10158 (.Y (nx10159), .A (nx10299)) ;
    inv02 ix10166 (.Y (nx10167), .A (nx10305)) ;
    inv02 ix10168 (.Y (nx10169), .A (nx10305)) ;
    inv02 ix10170 (.Y (nx10171), .A (nx10305)) ;
    inv02 ix10172 (.Y (nx10173), .A (nx10305)) ;
    inv02 ix10174 (.Y (nx10175), .A (nx10305)) ;
    inv02 ix10176 (.Y (nx10177), .A (nx10305)) ;
    inv02 ix10178 (.Y (nx10179), .A (nx10305)) ;
    inv02 ix10180 (.Y (nx10181), .A (nx10307)) ;
    inv02 ix10182 (.Y (nx10183), .A (nx10307)) ;
    inv02 ix10184 (.Y (nx10185), .A (nx10307)) ;
    inv02 ix10186 (.Y (nx10187), .A (nx10307)) ;
    inv02 ix10188 (.Y (nx10189), .A (nx10307)) ;
    inv02 ix10190 (.Y (nx10191), .A (nx10307)) ;
    inv02 ix10192 (.Y (nx10193), .A (nx10307)) ;
    inv02 ix10194 (.Y (nx10195), .A (nx10309)) ;
    inv02 ix10196 (.Y (nx10197), .A (nx10309)) ;
    inv02 ix10198 (.Y (nx10199), .A (nx10309)) ;
    inv02 ix10200 (.Y (nx10201), .A (nx10309)) ;
    inv02 ix10202 (.Y (nx10203), .A (nx10309)) ;
    inv02 ix10204 (.Y (nx10205), .A (nx10309)) ;
    inv02 ix10206 (.Y (nx10207), .A (nx10309)) ;
    inv02 ix10208 (.Y (nx10209), .A (nx10311)) ;
    inv02 ix10210 (.Y (nx10211), .A (nx10311)) ;
    inv02 ix10212 (.Y (nx10213), .A (nx10311)) ;
    inv02 ix10214 (.Y (nx10215), .A (nx10311)) ;
    inv02 ix10216 (.Y (nx10217), .A (nx10311)) ;
    inv02 ix10218 (.Y (nx10219), .A (nx10311)) ;
    inv02 ix10220 (.Y (nx10221), .A (nx10311)) ;
    inv02 ix10222 (.Y (nx10223), .A (nx10313)) ;
    inv02 ix10224 (.Y (nx10225), .A (nx10313)) ;
    inv02 ix10226 (.Y (nx10227), .A (nx10313)) ;
    inv02 ix10228 (.Y (nx10229), .A (nx10313)) ;
    inv02 ix10230 (.Y (nx10231), .A (nx10313)) ;
    inv02 ix10232 (.Y (nx10233), .A (nx10313)) ;
    inv02 ix10234 (.Y (nx10235), .A (nx10313)) ;
    inv02 ix10236 (.Y (nx10237), .A (nx10315)) ;
    inv02 ix10238 (.Y (nx10239), .A (nx10315)) ;
    inv02 ix10240 (.Y (nx10241), .A (nx10315)) ;
    inv02 ix10242 (.Y (nx10243), .A (nx10315)) ;
    inv02 ix10244 (.Y (nx10245), .A (nx10315)) ;
    inv02 ix10246 (.Y (nx10247), .A (nx10315)) ;
    inv02 ix10248 (.Y (nx10249), .A (nx10315)) ;
    inv02 ix10250 (.Y (nx10251), .A (nx10317)) ;
    inv02 ix10252 (.Y (nx10253), .A (nx10317)) ;
    inv02 ix10254 (.Y (nx10255), .A (nx10317)) ;
    inv02 ix10256 (.Y (nx10257), .A (nx10317)) ;
    inv02 ix10258 (.Y (nx10259), .A (nx10317)) ;
    inv02 ix10260 (.Y (nx10261), .A (nx10317)) ;
    inv02 ix10262 (.Y (nx10263), .A (nx10317)) ;
    inv02 ix10264 (.Y (nx10265), .A (nx10319)) ;
    inv02 ix10266 (.Y (nx10267), .A (nx10319)) ;
    inv02 ix10268 (.Y (nx10269), .A (nx10319)) ;
    inv02 ix10270 (.Y (nx10271), .A (nx10319)) ;
    inv02 ix10272 (.Y (nx10273), .A (nx10319)) ;
    inv02 ix10274 (.Y (nx10275), .A (nx10319)) ;
    inv02 ix10276 (.Y (nx10277), .A (nx10319)) ;
    inv02 ix10278 (.Y (nx10279), .A (nx10321)) ;
    inv02 ix10280 (.Y (nx10281), .A (nx10321)) ;
    inv02 ix10282 (.Y (nx10283), .A (nx10303)) ;
    inv02 ix10284 (.Y (nx10285), .A (nx10303)) ;
    inv02 ix10286 (.Y (nx10287), .A (nx10303)) ;
    inv02 ix10288 (.Y (nx10289), .A (nx10303)) ;
    inv02 ix10290 (.Y (nx10291), .A (nx10303)) ;
    inv02 ix10292 (.Y (nx10293), .A (nx10303)) ;
    inv02 ix10294 (.Y (nx10295), .A (nx10303)) ;
    inv02 ix10296 (.Y (nx10297), .A (nx10045)) ;
    inv02 ix10298 (.Y (nx10299), .A (nx10045)) ;
    inv02 ix10300 (.Y (nx10301), .A (CLK)) ;
    inv02 ix10302 (.Y (nx10303), .A (CLK)) ;
    inv02 ix10304 (.Y (nx10305), .A (EN)) ;
    inv02 ix10306 (.Y (nx10307), .A (nx10327)) ;
    inv02 ix10308 (.Y (nx10309), .A (nx10327)) ;
    inv02 ix10310 (.Y (nx10311), .A (nx10327)) ;
    inv02 ix10312 (.Y (nx10313), .A (nx10327)) ;
    inv02 ix10314 (.Y (nx10315), .A (nx10327)) ;
    inv02 ix10316 (.Y (nx10317), .A (nx10329)) ;
    inv02 ix10318 (.Y (nx10319), .A (nx10329)) ;
    inv02 ix10320 (.Y (nx10321), .A (nx10329)) ;
    inv01 ix10326 (.Y (nx10327), .A (nx10305)) ;
    inv01 ix10328 (.Y (nx10329), .A (nx10305)) ;
endmodule


module my_nadder_4 ( a, b, cin, s, cout ) ;

    input [3:0]a ;
    input [3:0]b ;
    input cin ;
    output [3:0]s ;
    output cout ;

    wire temp_2, temp_1, temp_0;



    my_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (s[0]), .cout (temp_0)) ;
    my_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (s[1]), .cout (
             temp_1)) ;
    my_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (s[2]), .cout (
             temp_2)) ;
    my_adder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (s[3]), .cout (
             cout)) ;
endmodule


module ReadBias ( current_state, BIAS, FilterAddress, DMAAddressToFilter, 
                  UpdatedAddress, changerAdd, CLK, RST, LayerInfo, outBias0, 
                  outBias1, outBias2, outBias3, outBias4, outBias5, outBias6, 
                  outBias7, ACKF ) ;

    input [14:0]current_state ;
    input [399:0]BIAS ;
    input [12:0]FilterAddress ;
    output [12:0]DMAAddressToFilter ;
    output [12:0]UpdatedAddress ;
    output [12:0]changerAdd ;
    input CLK ;
    input RST ;
    input [15:0]LayerInfo ;
    output [15:0]outBias0 ;
    output [15:0]outBias1 ;
    output [15:0]outBias2 ;
    output [15:0]outBias3 ;
    output [15:0]outBias4 ;
    output [15:0]outBias5 ;
    output [15:0]outBias6 ;
    output [15:0]outBias7 ;
    input ACKF ;

    wire upAddress_12, upAddress_11, upAddress_10, upAddress_9, upAddress_8, 
         upAddress_7, upAddress_6, upAddress_5, upAddress_4, upAddress_3, 
         upAddress_2, upAddress_1, upAddress_0, BiasEnable, Zeros_8, nx370, 
         nx372, nx374, nx376, nx378;
    wire [0:0] \$dummy ;




    nBitRegister_16 B0 (.D ({BIAS[15],BIAS[14],BIAS[13],BIAS[12],BIAS[11],
                    BIAS[10],BIAS[9],BIAS[8],BIAS[7],BIAS[6],BIAS[5],BIAS[4],
                    BIAS[3],BIAS[2],BIAS[1],BIAS[0]}), .CLK (nx372), .RST (RST)
                    , .EN (BiasEnable), .Q ({outBias0[15],outBias0[14],
                    outBias0[13],outBias0[12],outBias0[11],outBias0[10],
                    outBias0[9],outBias0[8],outBias0[7],outBias0[6],outBias0[5],
                    outBias0[4],outBias0[3],outBias0[2],outBias0[1],outBias0[0]}
                    )) ;
    nBitRegister_16 B1 (.D ({BIAS[31],BIAS[30],BIAS[29],BIAS[28],BIAS[27],
                    BIAS[26],BIAS[25],BIAS[24],BIAS[23],BIAS[22],BIAS[21],
                    BIAS[20],BIAS[19],BIAS[18],BIAS[17],BIAS[16]}), .CLK (nx372)
                    , .RST (RST), .EN (BiasEnable), .Q ({outBias1[15],
                    outBias1[14],outBias1[13],outBias1[12],outBias1[11],
                    outBias1[10],outBias1[9],outBias1[8],outBias1[7],outBias1[6]
                    ,outBias1[5],outBias1[4],outBias1[3],outBias1[2],outBias1[1]
                    ,outBias1[0]})) ;
    nBitRegister_16 B2 (.D ({BIAS[47],BIAS[46],BIAS[45],BIAS[44],BIAS[43],
                    BIAS[42],BIAS[41],BIAS[40],BIAS[39],BIAS[38],BIAS[37],
                    BIAS[36],BIAS[35],BIAS[34],BIAS[33],BIAS[32]}), .CLK (nx374)
                    , .RST (RST), .EN (BiasEnable), .Q ({outBias2[15],
                    outBias2[14],outBias2[13],outBias2[12],outBias2[11],
                    outBias2[10],outBias2[9],outBias2[8],outBias2[7],outBias2[6]
                    ,outBias2[5],outBias2[4],outBias2[3],outBias2[2],outBias2[1]
                    ,outBias2[0]})) ;
    nBitRegister_16 B3 (.D ({BIAS[63],BIAS[62],BIAS[61],BIAS[60],BIAS[59],
                    BIAS[58],BIAS[57],BIAS[56],BIAS[55],BIAS[54],BIAS[53],
                    BIAS[52],BIAS[51],BIAS[50],BIAS[49],BIAS[48]}), .CLK (nx374)
                    , .RST (RST), .EN (BiasEnable), .Q ({outBias3[15],
                    outBias3[14],outBias3[13],outBias3[12],outBias3[11],
                    outBias3[10],outBias3[9],outBias3[8],outBias3[7],outBias3[6]
                    ,outBias3[5],outBias3[4],outBias3[3],outBias3[2],outBias3[1]
                    ,outBias3[0]})) ;
    nBitRegister_16 B4 (.D ({BIAS[79],BIAS[78],BIAS[77],BIAS[76],BIAS[75],
                    BIAS[74],BIAS[73],BIAS[72],BIAS[71],BIAS[70],BIAS[69],
                    BIAS[68],BIAS[67],BIAS[66],BIAS[65],BIAS[64]}), .CLK (nx376)
                    , .RST (RST), .EN (BiasEnable), .Q ({outBias4[15],
                    outBias4[14],outBias4[13],outBias4[12],outBias4[11],
                    outBias4[10],outBias4[9],outBias4[8],outBias4[7],outBias4[6]
                    ,outBias4[5],outBias4[4],outBias4[3],outBias4[2],outBias4[1]
                    ,outBias4[0]})) ;
    nBitRegister_16 B5 (.D ({BIAS[95],BIAS[94],BIAS[93],BIAS[92],BIAS[91],
                    BIAS[90],BIAS[89],BIAS[88],BIAS[87],BIAS[86],BIAS[85],
                    BIAS[84],BIAS[83],BIAS[82],BIAS[81],BIAS[80]}), .CLK (nx376)
                    , .RST (RST), .EN (BiasEnable), .Q ({outBias5[15],
                    outBias5[14],outBias5[13],outBias5[12],outBias5[11],
                    outBias5[10],outBias5[9],outBias5[8],outBias5[7],outBias5[6]
                    ,outBias5[5],outBias5[4],outBias5[3],outBias5[2],outBias5[1]
                    ,outBias5[0]})) ;
    nBitRegister_16 B6 (.D ({BIAS[111],BIAS[110],BIAS[109],BIAS[108],BIAS[107],
                    BIAS[106],BIAS[105],BIAS[104],BIAS[103],BIAS[102],BIAS[101],
                    BIAS[100],BIAS[99],BIAS[98],BIAS[97],BIAS[96]}), .CLK (nx378
                    ), .RST (RST), .EN (BiasEnable), .Q ({outBias6[15],
                    outBias6[14],outBias6[13],outBias6[12],outBias6[11],
                    outBias6[10],outBias6[9],outBias6[8],outBias6[7],outBias6[6]
                    ,outBias6[5],outBias6[4],outBias6[3],outBias6[2],outBias6[1]
                    ,outBias6[0]})) ;
    nBitRegister_16 B7 (.D ({BIAS[127],BIAS[126],BIAS[125],BIAS[124],BIAS[123],
                    BIAS[122],BIAS[121],BIAS[120],BIAS[119],BIAS[118],BIAS[117],
                    BIAS[116],BIAS[115],BIAS[114],BIAS[113],BIAS[112]}), .CLK (
                    nx378), .RST (RST), .EN (BiasEnable), .Q ({outBias7[15],
                    outBias7[14],outBias7[13],outBias7[12],outBias7[11],
                    outBias7[10],outBias7[9],outBias7[8],outBias7[7],outBias7[6]
                    ,outBias7[5],outBias7[4],outBias7[3],outBias7[2],outBias7[1]
                    ,outBias7[0]})) ;
    triStateBuffer_13 tsb0 (.D ({FilterAddress[12],FilterAddress[11],
                      FilterAddress[10],FilterAddress[9],FilterAddress[8],
                      FilterAddress[7],FilterAddress[6],FilterAddress[5],
                      FilterAddress[4],FilterAddress[3],FilterAddress[2],
                      FilterAddress[1],FilterAddress[0]}), .EN (current_state[4]
                      ), .F ({DMAAddressToFilter[12],DMAAddressToFilter[11],
                      DMAAddressToFilter[10],DMAAddressToFilter[9],
                      DMAAddressToFilter[8],DMAAddressToFilter[7],
                      DMAAddressToFilter[6],DMAAddressToFilter[5],
                      DMAAddressToFilter[4],DMAAddressToFilter[3],
                      DMAAddressToFilter[2],DMAAddressToFilter[1],
                      DMAAddressToFilter[0]})) ;
    my_nadder_13 adder0 (.a ({FilterAddress[12],FilterAddress[11],
                 FilterAddress[10],FilterAddress[9],FilterAddress[8],
                 FilterAddress[7],FilterAddress[6],FilterAddress[5],
                 FilterAddress[4],FilterAddress[3],FilterAddress[2],
                 FilterAddress[1],FilterAddress[0]}), .b ({Zeros_8,Zeros_8,
                 Zeros_8,Zeros_8,Zeros_8,Zeros_8,Zeros_8,Zeros_8,Zeros_8,
                 LayerInfo[3],LayerInfo[2],LayerInfo[1],LayerInfo[0]}), .cin (
                 Zeros_8), .s ({upAddress_12,upAddress_11,upAddress_10,
                 upAddress_9,upAddress_8,upAddress_7,upAddress_6,upAddress_5,
                 upAddress_4,upAddress_3,upAddress_2,upAddress_1,upAddress_0}), 
                 .cout (\$dummy [0])) ;
    triStateBuffer_13 TriStateAdd (.D ({upAddress_12,upAddress_11,upAddress_10,
                      upAddress_9,upAddress_8,upAddress_7,upAddress_6,
                      upAddress_5,upAddress_4,upAddress_3,upAddress_2,
                      upAddress_1,upAddress_0}), .EN (current_state[4]), .F ({
                      UpdatedAddress[12],UpdatedAddress[11],UpdatedAddress[10],
                      UpdatedAddress[9],UpdatedAddress[8],UpdatedAddress[7],
                      UpdatedAddress[6],UpdatedAddress[5],UpdatedAddress[4],
                      UpdatedAddress[3],UpdatedAddress[2],UpdatedAddress[1],
                      UpdatedAddress[0]})) ;
    triStateBuffer_13 TriStateAddchanger (.D ({upAddress_12,upAddress_11,
                      upAddress_10,upAddress_9,upAddress_8,upAddress_7,
                      upAddress_6,upAddress_5,upAddress_4,upAddress_3,
                      upAddress_2,upAddress_1,upAddress_0}), .EN (
                      current_state[4]), .F ({changerAdd[12],changerAdd[11],
                      changerAdd[10],changerAdd[9],changerAdd[8],changerAdd[7],
                      changerAdd[6],changerAdd[5],changerAdd[4],changerAdd[3],
                      changerAdd[2],changerAdd[1],changerAdd[0]})) ;
    fake_gnd ix355 (.Y (Zeros_8)) ;
    and02 ix1 (.Y (BiasEnable), .A0 (ACKF), .A1 (current_state[4])) ;
    inv01 ix369 (.Y (nx370), .A (CLK)) ;
    inv02 ix371 (.Y (nx372), .A (nx370)) ;
    inv02 ix373 (.Y (nx374), .A (nx370)) ;
    inv02 ix375 (.Y (nx376), .A (nx370)) ;
    inv02 ix377 (.Y (nx378), .A (nx370)) ;
endmodule


module CalculateInfo ( WSquareOut, CounOut, LayerInfoIn, clk, rst, current_state, 
                       ACK, ACKI, Wmin1 ) ;

    output [9:0]WSquareOut ;
    output [1:0]CounOut ;
    input [15:0]LayerInfoIn ;
    input clk ;
    input rst ;
    input [14:0]current_state ;
    output ACK ;
    input ACKI ;
    output [4:0]Wmin1 ;

    wire CountereEN, CountereRST, GND0, PWR, nx0, nx2, nx12, nx38, nx42, nx46, 
         nx48, nx54, nx58, nx60, nx86, nx88, nx110, nx116, nx130, nx132, nx146, 
         nx148, nx172, nx180, nx182, nx190, nx192, nx206, nx208, nx232, nx236, 
         nx240, nx274, nx290, nx111, nx123, nx129, nx131, nx139, nx141, nx143, 
         nx147, nx157, nx159, nx161, nx163, nx167, nx173, nx183, nx185, nx187, 
         nx189, nx191, nx195, nx197, nx199, nx201, nx203, nx205, nx207, nx209, 
         nx211, nx213, nx215, nx217, nx219, nx227, nx231, nx239, nx241, nx243, 
         nx245, nx247, nx255, nx263, nx265, nx267, nx279, nx291, nx293, nx295, 
         nx297;
    wire [1:0] \$dummy ;




    my_nadder_5 adder (.a ({LayerInfoIn[8],LayerInfoIn[7],LayerInfoIn[6],nx291,
                nx295}), .b ({PWR,PWR,PWR,PWR,PWR}), .cin (GND0), .s ({Wmin1[4],
                Wmin1[3],Wmin1[2],Wmin1[1],Wmin1[0]}), .cout (\$dummy [0])) ;
    Counter_2 EndCounter (.enable (CountereEN), .reset (CountereRST), .clk (clk)
              , .load (GND0), .\output  ({CounOut[1],CounOut[0]}), .\input  ({
              GND0,GND0})) ;
    fake_vcc ix81 (.Y (PWR)) ;
    fake_gnd ix79 (.Y (GND0)) ;
    ao221 ix285 (.Y (CountereRST), .A0 (CounOut[1]), .A1 (nx111), .B0 (ACKI), .B1 (
          nx274), .C0 (rst)) ;
    inv01 ix112 (.Y (nx111), .A (CounOut[0])) ;
    or02 ix275 (.Y (nx274), .A0 (current_state[2]), .A1 (current_state[4])) ;
    nor02_2x ix301 (.Y (CountereEN), .A0 (ACK), .A1 (nx123)) ;
    dffs_ni reg_ACKW_dup_1 (.Q (ACK), .QB (\$dummy [1]), .D (GND0), .CLK (clk), 
            .S (nx290)) ;
    nor02ii ix291 (.Y (nx290), .A0 (CounOut[1]), .A1 (CounOut[0])) ;
    nor02_2x ix124 (.Y (nx123), .A0 (current_state[2]), .A1 (current_state[4])
             ) ;
    and02 ix215 (.Y (WSquareOut[0]), .A0 (Wmin1[0]), .A1 (nx295)) ;
    nor02ii ix273 (.Y (WSquareOut[1]), .A0 (nx129), .A1 (nx131)) ;
    aoi22 ix130 (.Y (nx129), .A0 (nx291), .A1 (Wmin1[0]), .B0 (Wmin1[1]), .B1 (
          nx295)) ;
    nand03 ix132 (.Y (nx131), .A0 (WSquareOut[0]), .A1 (nx291), .A2 (Wmin1[1])
           ) ;
    xnor2 ix263 (.Y (WSquareOut[2]), .A0 (nx131), .A1 (nx208)) ;
    xnor2 ix209 (.Y (nx208), .A0 (nx206), .A1 (nx143)) ;
    nor02ii ix207 (.Y (nx206), .A0 (nx139), .A1 (nx141)) ;
    aoi22 ix140 (.Y (nx139), .A0 (Wmin1[2]), .A1 (nx295), .B0 (nx291), .B1 (
          Wmin1[1])) ;
    nand04 ix142 (.Y (nx141), .A0 (nx291), .A1 (Wmin1[1]), .A2 (Wmin1[2]), .A3 (
           nx295)) ;
    nand02 ix144 (.Y (nx143), .A0 (LayerInfoIn[6]), .A1 (Wmin1[0])) ;
    xnor2 ix261 (.Y (WSquareOut[3]), .A0 (nx147), .A1 (nx192)) ;
    mux21_ni ix148 (.Y (nx147), .A0 (nx143), .A1 (nx131), .S0 (nx208)) ;
    xnor2 ix193 (.Y (nx192), .A0 (nx190), .A1 (nx163)) ;
    xnor2 ix191 (.Y (nx190), .A0 (nx141), .A1 (nx148)) ;
    xnor2 ix149 (.Y (nx148), .A0 (nx146), .A1 (nx161)) ;
    nor02ii ix147 (.Y (nx146), .A0 (nx157), .A1 (nx159)) ;
    aoi22 ix158 (.Y (nx157), .A0 (nx291), .A1 (Wmin1[2]), .B0 (Wmin1[3]), .B1 (
          nx295)) ;
    nand04 ix160 (.Y (nx159), .A0 (Wmin1[3]), .A1 (nx297), .A2 (nx293), .A3 (
           Wmin1[2])) ;
    nand02 ix162 (.Y (nx161), .A0 (LayerInfoIn[6]), .A1 (Wmin1[1])) ;
    nand02 ix164 (.Y (nx163), .A0 (LayerInfoIn[7]), .A1 (Wmin1[0])) ;
    xnor2 ix259 (.Y (WSquareOut[4]), .A0 (nx167), .A1 (nx182)) ;
    mux21_ni ix168 (.Y (nx167), .A0 (nx163), .A1 (nx147), .S0 (nx192)) ;
    xnor2 ix183 (.Y (nx182), .A0 (nx180), .A1 (nx191)) ;
    xnor2 ix181 (.Y (nx180), .A0 (nx173), .A1 (nx132)) ;
    mux21_ni ix174 (.Y (nx173), .A0 (nx161), .A1 (nx141), .S0 (nx148)) ;
    xnor2 ix133 (.Y (nx132), .A0 (nx130), .A1 (nx189)) ;
    xnor2 ix131 (.Y (nx130), .A0 (nx159), .A1 (nx88)) ;
    xnor2 ix89 (.Y (nx88), .A0 (nx86), .A1 (nx187)) ;
    nor02ii ix87 (.Y (nx86), .A0 (nx183), .A1 (nx185)) ;
    aoi22 ix184 (.Y (nx183), .A0 (nx293), .A1 (Wmin1[3]), .B0 (Wmin1[4]), .B1 (
          nx297)) ;
    nand04 ix186 (.Y (nx185), .A0 (nx293), .A1 (Wmin1[4]), .A2 (Wmin1[3]), .A3 (
           nx297)) ;
    nand02 ix188 (.Y (nx187), .A0 (LayerInfoIn[6]), .A1 (Wmin1[2])) ;
    nand02 ix190 (.Y (nx189), .A0 (LayerInfoIn[7]), .A1 (Wmin1[1])) ;
    nand02 ix192 (.Y (nx191), .A0 (LayerInfoIn[8]), .A1 (Wmin1[0])) ;
    xor2 ix257 (.Y (WSquareOut[5]), .A0 (nx195), .A1 (nx197)) ;
    mux21_ni ix196 (.Y (nx195), .A0 (nx191), .A1 (nx167), .S0 (nx182)) ;
    xnor2 ix198 (.Y (nx197), .A0 (nx199), .A1 (nx201)) ;
    mux21_ni ix200 (.Y (nx199), .A0 (nx189), .A1 (nx173), .S0 (nx132)) ;
    xnor2 ix202 (.Y (nx201), .A0 (nx203), .A1 (nx219)) ;
    xnor2 ix204 (.Y (nx203), .A0 (nx205), .A1 (nx207)) ;
    mux21_ni ix206 (.Y (nx205), .A0 (nx187), .A1 (nx159), .S0 (nx88)) ;
    xnor2 ix208 (.Y (nx207), .A0 (nx209), .A1 (nx217)) ;
    xnor2 ix210 (.Y (nx209), .A0 (nx185), .A1 (nx211)) ;
    xnor2 ix212 (.Y (nx211), .A0 (nx213), .A1 (nx215)) ;
    nand02 ix214 (.Y (nx213), .A0 (nx293), .A1 (Wmin1[4])) ;
    nand02 ix216 (.Y (nx215), .A0 (LayerInfoIn[6]), .A1 (Wmin1[3])) ;
    nand02 ix218 (.Y (nx217), .A0 (LayerInfoIn[7]), .A1 (Wmin1[2])) ;
    nand02 ix220 (.Y (nx219), .A0 (LayerInfoIn[8]), .A1 (Wmin1[1])) ;
    xor2 ix251 (.Y (WSquareOut[6]), .A0 (nx232), .A1 (nx172)) ;
    nor02_2x ix233 (.Y (nx232), .A0 (nx195), .A1 (nx197)) ;
    xnor2 ix173 (.Y (nx172), .A0 (nx227), .A1 (nx116)) ;
    mux21_ni ix228 (.Y (nx227), .A0 (nx199), .A1 (nx219), .S0 (nx201)) ;
    xnor2 ix117 (.Y (nx116), .A0 (nx231), .A1 (nx60)) ;
    mux21_ni ix232 (.Y (nx231), .A0 (nx205), .A1 (nx217), .S0 (nx207)) ;
    xnor2 ix61 (.Y (nx60), .A0 (nx58), .A1 (nx247)) ;
    xnor2 ix59 (.Y (nx58), .A0 (nx38), .A1 (nx241)) ;
    aoi21 ix39 (.Y (nx38), .A0 (nx239), .A1 (nx215), .B0 (nx213)) ;
    nand02 ix240 (.Y (nx239), .A0 (Wmin1[3]), .A1 (nx297)) ;
    xnor2 ix242 (.Y (nx241), .A0 (nx243), .A1 (nx245)) ;
    nand02 ix244 (.Y (nx243), .A0 (LayerInfoIn[6]), .A1 (Wmin1[4])) ;
    nand02 ix246 (.Y (nx245), .A0 (LayerInfoIn[7]), .A1 (Wmin1[3])) ;
    nand02 ix248 (.Y (nx247), .A0 (LayerInfoIn[8]), .A1 (Wmin1[2])) ;
    xor2 ix249 (.Y (WSquareOut[7]), .A0 (nx236), .A1 (nx110)) ;
    mux21_ni ix237 (.Y (nx236), .A0 (nx116), .A1 (nx232), .S0 (nx172)) ;
    xnor2 ix111 (.Y (nx110), .A0 (nx255), .A1 (nx54)) ;
    mux21_ni ix256 (.Y (nx255), .A0 (nx247), .A1 (nx231), .S0 (nx60)) ;
    xnor2 ix55 (.Y (nx54), .A0 (nx42), .A1 (nx263)) ;
    mux21_ni ix43 (.Y (nx42), .A0 (nx38), .A1 (nx12), .S0 (nx241)) ;
    xnor2 ix264 (.Y (nx263), .A0 (nx265), .A1 (nx267)) ;
    nand02 ix266 (.Y (nx265), .A0 (LayerInfoIn[7]), .A1 (Wmin1[4])) ;
    nand02 ix268 (.Y (nx267), .A0 (LayerInfoIn[8]), .A1 (Wmin1[3])) ;
    xor2 ix247 (.Y (WSquareOut[8]), .A0 (nx240), .A1 (nx48)) ;
    mux21_ni ix241 (.Y (nx240), .A0 (nx54), .A1 (nx236), .S0 (nx110)) ;
    xnor2 ix49 (.Y (nx48), .A0 (nx46), .A1 (nx279)) ;
    mux21_ni ix47 (.Y (nx46), .A0 (nx42), .A1 (nx2), .S0 (nx263)) ;
    nand02 ix280 (.Y (nx279), .A0 (LayerInfoIn[8]), .A1 (Wmin1[4])) ;
    mux21_ni ix245 (.Y (WSquareOut[9]), .A0 (nx0), .A1 (nx240), .S0 (nx48)) ;
    inv01 ix13 (.Y (nx12), .A (nx245)) ;
    inv01 ix3 (.Y (nx2), .A (nx267)) ;
    inv01 ix1 (.Y (nx0), .A (nx279)) ;
    buf02 ix289 (.Y (nx291), .A (LayerInfoIn[5])) ;
    buf02 ix292 (.Y (nx293), .A (LayerInfoIn[5])) ;
    buf02 ix294 (.Y (nx295), .A (LayerInfoIn[4])) ;
    buf02 ix296 (.Y (nx297), .A (LayerInfoIn[4])) ;
endmodule


module Counter_2 ( enable, reset, clk, load, \output , \input  ) ;

    input enable ;
    input reset ;
    input clk ;
    input load ;
    output [1:0]\output  ;
    input [1:0]\input  ;

    wire addResult_1, addResult_0, one_0, one_1, nx28, NOT_clk, nx8, nx12, nx22, 
         nx20, nx25, nx85, nx95, nx104;
    wire [4:0] \$dummy ;




    my_nadder_2 A1 (.a ({\output [1],\output [0]}), .b ({one_1,one_0}), .cin (
                one_1), .s ({addResult_1,addResult_0}), .cout (\$dummy [0])) ;
    fake_gnd ix68 (.Y (one_1)) ;
    fake_vcc ix66 (.Y (one_0)) ;
    dffsr_ni reg_toOutput_0__dup_1 (.Q (\output [0]), .QB (\$dummy [1]), .D (
             nx85), .CLK (clk), .S (nx8), .R (nx12)) ;
    mux21_ni ix86 (.Y (nx85), .A0 (\output [0]), .A1 (addResult_0), .S0 (enable)
             ) ;
    nor02ii ix9 (.Y (nx8), .A0 (nx104), .A1 (nx28)) ;
    nor02_2x ix105 (.Y (nx104), .A0 (reset), .A1 (load)) ;
    dffr ix29 (.Q (nx28), .QB (\$dummy [2]), .D (\input [0]), .CLK (NOT_clk), .R (
         reset)) ;
    inv01 ix108 (.Y (NOT_clk), .A (clk)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (nx28), .A1 (nx104)) ;
    dffsr_ni reg_toOutput_1__dup_1 (.Q (\output [1]), .QB (\$dummy [3]), .D (
             nx95), .CLK (clk), .S (nx20), .R (nx25)) ;
    mux21_ni ix96 (.Y (nx95), .A0 (\output [1]), .A1 (addResult_1), .S0 (enable)
             ) ;
    nor02ii ix21 (.Y (nx20), .A0 (nx104), .A1 (nx22)) ;
    dffr ix23 (.Q (nx22), .QB (\$dummy [4]), .D (\input [1]), .CLK (NOT_clk), .R (
         reset)) ;
    nor02_2x ix26 (.Y (nx25), .A0 (nx22), .A1 (nx104)) ;
endmodule


module my_nadder_2 ( a, b, cin, s, cout ) ;

    input [1:0]a ;
    input [1:0]b ;
    input cin ;
    output [1:0]s ;
    output cout ;

    wire temp_0;



    my_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (s[0]), .cout (temp_0)) ;
    my_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (s[1]), .cout (
             cout)) ;
endmodule


module my_nadder_5 ( a, b, cin, s, cout ) ;

    input [4:0]a ;
    input [4:0]b ;
    input cin ;
    output [4:0]s ;
    output cout ;

    wire temp_3, temp_2, temp_1, temp_0;



    my_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (s[0]), .cout (temp_0)) ;
    my_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (s[1]), .cout (
             temp_1)) ;
    my_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (s[2]), .cout (
             temp_2)) ;
    my_adder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (s[3]), .cout (
             temp_3)) ;
    my_adder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (s[4]), .cout (
             cout)) ;
endmodule


module ReadLayerInfo ( LayerInfoIn, ImgWidthIn, FilterAdd, ImgAdd, clk, rst, 
                       ACKF, ACKI, current_state, LayerInfoOut, ImgWidthOut, 
                       FilterAddToDMA, ImgAddToDMA ) ;

    input [15:0]LayerInfoIn ;
    input [15:0]ImgWidthIn ;
    input [12:0]FilterAdd ;
    input [12:0]ImgAdd ;
    input clk ;
    input rst ;
    input ACKF ;
    input ACKI ;
    input [14:0]current_state ;
    output [15:0]LayerInfoOut ;
    output [15:0]ImgWidthOut ;
    output [12:0]FilterAddToDMA ;
    output [12:0]ImgAddToDMA ;

    wire LayerInfEN, ImgWidthEN;



    nBitRegister_16 LayerInf (.D ({LayerInfoIn[15],LayerInfoIn[14],
                    LayerInfoIn[13],LayerInfoIn[12],LayerInfoIn[11],
                    LayerInfoIn[10],LayerInfoIn[9],LayerInfoIn[8],LayerInfoIn[7]
                    ,LayerInfoIn[6],LayerInfoIn[5],LayerInfoIn[4],LayerInfoIn[3]
                    ,LayerInfoIn[2],LayerInfoIn[1],LayerInfoIn[0]}), .CLK (clk)
                    , .RST (rst), .EN (LayerInfEN), .Q ({LayerInfoOut[15],
                    LayerInfoOut[14],LayerInfoOut[13],LayerInfoOut[12],
                    LayerInfoOut[11],LayerInfoOut[10],LayerInfoOut[9],
                    LayerInfoOut[8],LayerInfoOut[7],LayerInfoOut[6],
                    LayerInfoOut[5],LayerInfoOut[4],LayerInfoOut[3],
                    LayerInfoOut[2],LayerInfoOut[1],LayerInfoOut[0]})) ;
    nBitRegister_16 ImgWidth (.D ({ImgWidthIn[15],ImgWidthIn[14],ImgWidthIn[13],
                    ImgWidthIn[12],ImgWidthIn[11],ImgWidthIn[10],ImgWidthIn[9],
                    ImgWidthIn[8],ImgWidthIn[7],ImgWidthIn[6],ImgWidthIn[5],
                    ImgWidthIn[4],ImgWidthIn[3],ImgWidthIn[2],ImgWidthIn[1],
                    ImgWidthIn[0]}), .CLK (clk), .RST (rst), .EN (ImgWidthEN), .Q (
                    {ImgWidthOut[15],ImgWidthOut[14],ImgWidthOut[13],
                    ImgWidthOut[12],ImgWidthOut[11],ImgWidthOut[10],
                    ImgWidthOut[9],ImgWidthOut[8],ImgWidthOut[7],ImgWidthOut[6],
                    ImgWidthOut[5],ImgWidthOut[4],ImgWidthOut[3],ImgWidthOut[2],
                    ImgWidthOut[1],ImgWidthOut[0]})) ;
    triStateBuffer_13 FilterAddTriDMA (.D ({FilterAdd[12],FilterAdd[11],
                      FilterAdd[10],FilterAdd[9],FilterAdd[8],FilterAdd[7],
                      FilterAdd[6],FilterAdd[5],FilterAdd[4],FilterAdd[3],
                      FilterAdd[2],FilterAdd[1],FilterAdd[0]}), .EN (
                      current_state[1]), .F ({FilterAddToDMA[12],
                      FilterAddToDMA[11],FilterAddToDMA[10],FilterAddToDMA[9],
                      FilterAddToDMA[8],FilterAddToDMA[7],FilterAddToDMA[6],
                      FilterAddToDMA[5],FilterAddToDMA[4],FilterAddToDMA[3],
                      FilterAddToDMA[2],FilterAddToDMA[1],FilterAddToDMA[0]})) ;
    triStateBuffer_13 ImgAddTriDMA (.D ({ImgAdd[12],ImgAdd[11],ImgAdd[10],
                      ImgAdd[9],ImgAdd[8],ImgAdd[7],ImgAdd[6],ImgAdd[5],
                      ImgAdd[4],ImgAdd[3],ImgAdd[2],ImgAdd[1],ImgAdd[0]}), .EN (
                      current_state[1]), .F ({ImgAddToDMA[12],ImgAddToDMA[11],
                      ImgAddToDMA[10],ImgAddToDMA[9],ImgAddToDMA[8],
                      ImgAddToDMA[7],ImgAddToDMA[6],ImgAddToDMA[5],
                      ImgAddToDMA[4],ImgAddToDMA[3],ImgAddToDMA[2],
                      ImgAddToDMA[1],ImgAddToDMA[0]})) ;
    and02 ix1 (.Y (ImgWidthEN), .A0 (ACKI), .A1 (current_state[1])) ;
    and02 ix3 (.Y (LayerInfEN), .A0 (ACKF), .A1 (current_state[1])) ;
endmodule


module my_nadder_13 ( a, b, cin, s, cout ) ;

    input [12:0]a ;
    input [12:0]b ;
    input cin ;
    output [12:0]s ;
    output cout ;

    wire temp_11, temp_10, temp_9, temp_8, temp_7, temp_6, temp_5, temp_4, 
         temp_3, temp_2, temp_1, temp_0;



    my_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (s[0]), .cout (temp_0)) ;
    my_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (s[1]), .cout (
             temp_1)) ;
    my_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (s[2]), .cout (
             temp_2)) ;
    my_adder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (s[3]), .cout (
             temp_3)) ;
    my_adder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (s[4]), .cout (
             temp_4)) ;
    my_adder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (s[5]), .cout (
             temp_5)) ;
    my_adder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (s[6]), .cout (
             temp_6)) ;
    my_adder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (s[7]), .cout (
             temp_7)) ;
    my_adder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (s[8]), .cout (
             temp_8)) ;
    my_adder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (s[9]), .cout (
             temp_9)) ;
    my_adder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (s[10]), .cout (
             temp_10)) ;
    my_adder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (s[11]), .cout (
             temp_11)) ;
    my_adder loop1_12_fx (.a (a[12]), .b (b[12]), .cin (temp_11), .s (s[12]), .cout (
             cout)) ;
endmodule


module my_adder ( a, b, cin, s, cout ) ;

    input a ;
    input b ;
    input cin ;
    output s ;
    output cout ;

    wire nx0, nx69;



    ao22 ix7 (.Y (cout), .A0 (b), .A1 (a), .B0 (cin), .B1 (nx0)) ;
    xnor2 ix9 (.Y (s), .A0 (nx69), .A1 (cin)) ;
    xnor2 ix70 (.Y (nx69), .A0 (a), .A1 (b)) ;
    inv01 ix1 (.Y (nx0), .A (nx69)) ;
endmodule


module ReadInfoState ( CLK, S, reset, MFC, filterAddressReg_out, filterRamData, 
                       noOfLayersReg_out, filterRamAddress ) ;

    input CLK ;
    input [14:0]S ;
    input reset ;
    input MFC ;
    input [12:0]filterAddressReg_out ;
    input [15:0]filterRamData ;
    output [15:0]noOfLayersReg_out ;
    output [12:0]filterRamAddress ;




    nBitRegister_16 noOfLayersReg (.D ({filterRamData[15],filterRamData[14],
                    filterRamData[13],filterRamData[12],filterRamData[11],
                    filterRamData[10],filterRamData[9],filterRamData[8],
                    filterRamData[7],filterRamData[6],filterRamData[5],
                    filterRamData[4],filterRamData[3],filterRamData[2],
                    filterRamData[1],filterRamData[0]}), .CLK (CLK), .RST (reset
                    ), .EN (S[0]), .Q ({noOfLayersReg_out[15],
                    noOfLayersReg_out[14],noOfLayersReg_out[13],
                    noOfLayersReg_out[12],noOfLayersReg_out[11],
                    noOfLayersReg_out[10],noOfLayersReg_out[9],
                    noOfLayersReg_out[8],noOfLayersReg_out[7],
                    noOfLayersReg_out[6],noOfLayersReg_out[5],
                    noOfLayersReg_out[4],noOfLayersReg_out[3],
                    noOfLayersReg_out[2],noOfLayersReg_out[1],
                    noOfLayersReg_out[0]})) ;
    triStateBuffer_13 dmaOut (.D ({filterAddressReg_out[12],
                      filterAddressReg_out[11],filterAddressReg_out[10],
                      filterAddressReg_out[9],filterAddressReg_out[8],
                      filterAddressReg_out[7],filterAddressReg_out[6],
                      filterAddressReg_out[5],filterAddressReg_out[4],
                      filterAddressReg_out[3],filterAddressReg_out[2],
                      filterAddressReg_out[1],filterAddressReg_out[0]}), .EN (
                      S[0]), .F ({filterRamAddress[12],filterRamAddress[11],
                      filterRamAddress[10],filterRamAddress[9],
                      filterRamAddress[8],filterRamAddress[7],
                      filterRamAddress[6],filterRamAddress[5],
                      filterRamAddress[4],filterRamAddress[3],
                      filterRamAddress[2],filterRamAddress[1],
                      filterRamAddress[0]})) ;
endmodule


module nBitRegister_16 ( D, CLK, RST, EN, Q ) ;

    input [15:0]D ;
    input CLK ;
    input RST ;
    input EN ;
    output [15:0]Q ;

    wire nx230, nx240, nx250, nx260, nx270, nx280, nx290, nx300, nx310, nx320, 
         nx330, nx340, nx350, nx360, nx370, nx380, nx445, nx447, nx449, nx455, 
         nx457, nx459, nx461;
    wire [15:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx230), .CLK (nx445), .R (
         RST)) ;
    mux21_ni ix231 (.Y (nx230), .A0 (Q[0]), .A1 (D[0]), .S0 (nx457)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx240), .CLK (nx445), .R (
         RST)) ;
    mux21_ni ix241 (.Y (nx240), .A0 (Q[1]), .A1 (D[1]), .S0 (nx457)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx250), .CLK (nx445), .R (
         RST)) ;
    mux21_ni ix251 (.Y (nx250), .A0 (Q[2]), .A1 (D[2]), .S0 (nx457)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx260), .CLK (nx445), .R (
         RST)) ;
    mux21_ni ix261 (.Y (nx260), .A0 (Q[3]), .A1 (D[3]), .S0 (nx457)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx270), .CLK (nx445), .R (
         RST)) ;
    mux21_ni ix271 (.Y (nx270), .A0 (Q[4]), .A1 (D[4]), .S0 (nx457)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx280), .CLK (nx445), .R (
         RST)) ;
    mux21_ni ix281 (.Y (nx280), .A0 (Q[5]), .A1 (D[5]), .S0 (nx457)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx290), .CLK (nx445), .R (
         RST)) ;
    mux21_ni ix291 (.Y (nx290), .A0 (Q[6]), .A1 (D[6]), .S0 (nx457)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx300), .CLK (nx447), .R (
         RST)) ;
    mux21_ni ix301 (.Y (nx300), .A0 (Q[7]), .A1 (D[7]), .S0 (nx459)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx310), .CLK (nx447), .R (
         RST)) ;
    mux21_ni ix311 (.Y (nx310), .A0 (Q[8]), .A1 (D[8]), .S0 (nx459)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx320), .CLK (nx447), .R (
         RST)) ;
    mux21_ni ix321 (.Y (nx320), .A0 (Q[9]), .A1 (D[9]), .S0 (nx459)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx330), .CLK (nx447), .R (
         RST)) ;
    mux21_ni ix331 (.Y (nx330), .A0 (Q[10]), .A1 (D[10]), .S0 (nx459)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx340), .CLK (nx447), .R (
         RST)) ;
    mux21_ni ix341 (.Y (nx340), .A0 (Q[11]), .A1 (D[11]), .S0 (nx459)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx350), .CLK (nx447), .R (
         RST)) ;
    mux21_ni ix351 (.Y (nx350), .A0 (Q[12]), .A1 (D[12]), .S0 (nx459)) ;
    dffr reg_Q_13 (.Q (Q[13]), .QB (\$dummy [13]), .D (nx360), .CLK (nx447), .R (
         RST)) ;
    mux21_ni ix361 (.Y (nx360), .A0 (Q[13]), .A1 (D[13]), .S0 (nx459)) ;
    dffr reg_Q_14 (.Q (Q[14]), .QB (\$dummy [14]), .D (nx370), .CLK (nx449), .R (
         RST)) ;
    mux21_ni ix371 (.Y (nx370), .A0 (Q[14]), .A1 (D[14]), .S0 (nx461)) ;
    dffr reg_Q_15 (.Q (Q[15]), .QB (\$dummy [15]), .D (nx380), .CLK (nx449), .R (
         RST)) ;
    mux21_ni ix381 (.Y (nx380), .A0 (Q[15]), .A1 (D[15]), .S0 (nx461)) ;
    inv02 ix444 (.Y (nx445), .A (CLK)) ;
    inv02 ix446 (.Y (nx447), .A (CLK)) ;
    inv02 ix448 (.Y (nx449), .A (CLK)) ;
    inv01 ix454 (.Y (nx455), .A (EN)) ;
    inv02 ix456 (.Y (nx457), .A (nx455)) ;
    inv02 ix458 (.Y (nx459), .A (nx455)) ;
    inv02 ix460 (.Y (nx461), .A (nx455)) ;
endmodule


module memoryDMA ( resetEN, AddressIn, dataIn, switcherEN, ramSelector, readEn, 
                   writeEn, CLK, Normal, MFC, counterOut, dataOut ) ;

    input resetEN ;
    input [12:0]AddressIn ;
    input [15:0]dataIn ;
    input switcherEN ;
    input ramSelector ;
    input readEn ;
    input writeEn ;
    input CLK ;
    input Normal ;
    output MFC ;
    output [3:0]counterOut ;
    output [447:0]dataOut ;

    wire dataFromRam1_447, dataFromRam2_447, dataToRam1_15, dataToRam1_14, 
         dataToRam1_13, dataToRam1_12, dataToRam1_11, dataToRam1_10, 
         dataToRam1_9, dataToRam1_8, dataToRam1_7, dataToRam1_6, dataToRam1_5, 
         dataToRam1_4, dataToRam1_3, dataToRam1_2, dataToRam1_1, dataToRam1_0, 
         dataToRam2_15, dataToRam2_14, dataToRam2_13, dataToRam2_12, 
         dataToRam2_11, dataToRam2_10, dataToRam2_9, dataToRam2_8, dataToRam2_7, 
         dataToRam2_6, dataToRam2_5, dataToRam2_4, dataToRam2_3, dataToRam2_2, 
         dataToRam2_1, dataToRam2_0, mfcOfRam1, mfcOfRam2, DInput, ram2Read, 
         ram1Read, ram2Write, ram1Write, GND, test, nx5632, nx5653, nx5655, 
         nx5657, nx5659, nx5661, nx5663, nx5665, nx5667, nx5669, nx5671, nx5673, 
         nx5675, nx5677, nx5679, nx5681, nx5683, nx5685, nx5687, nx5689, nx5691, 
         nx5693, nx5695, nx5697, nx5699, nx5701, nx5703, nx5705, nx5707, nx5709, 
         nx5711, nx5713, nx5715, nx5717, nx5719, nx5721, nx5723, nx5725, nx5727, 
         nx5729, nx5731, nx5733, nx5735, nx5737, nx5739, nx5741, nx5743, nx5745, 
         nx5747, nx5749, nx5751, nx5753, nx5755, nx5757, nx5759, nx5761, nx5763, 
         nx5765, nx5767, nx5769, nx5771, nx5773, nx5775, nx5777, nx5779, nx5781, 
         nx5783, nx5785, nx5787, nx5789, nx5791, nx5793, nx5795, nx5797, nx5799, 
         nx5801, nx5803, nx5805, nx5807, nx5809, nx5811, nx5813, nx5815, nx5817, 
         nx5819, nx5821, nx5823, nx5825, nx5827, nx5829, nx5831, nx5833, nx5835, 
         nx5837, nx5839, nx5841, nx5843, nx5845, nx5847, nx5849, nx5851, nx5853, 
         nx5855, nx5857, nx5859, nx5861, nx5863, nx5865, nx5867, nx5869, nx5871, 
         nx5873, nx5875, nx5877, nx5879, nx5881, nx5883, nx5885, nx5887, nx5889, 
         nx5891, nx5893, nx5895, nx5897, nx5899, nx5901, nx5903, nx5905, nx5907, 
         nx5909, nx5911, nx5913, nx5915, nx5917, nx5919, nx5921, nx5923, nx5925, 
         nx5927, nx5929, nx5931, nx5933, nx5935, nx5937, nx5939, nx5941, nx5943, 
         nx5945, nx5947, nx5953, nx5955, nx5957, nx5959;
    wire [901:0] \$dummy ;




    triStateBuffer_448 Ram1Rd (.D ({nx5655,nx5655,nx5655,nx5655,nx5655,nx5655,
                       nx5655,nx5657,nx5657,nx5657,nx5657,nx5657,nx5657,nx5657,
                       nx5659,nx5659,nx5659,nx5659,nx5659,nx5659,nx5659,nx5661,
                       nx5661,nx5661,nx5661,nx5661,nx5661,nx5661,nx5663,nx5663,
                       nx5663,nx5663,nx5663,nx5663,nx5663,nx5665,nx5665,nx5665,
                       nx5665,nx5665,nx5665,nx5665,nx5667,nx5667,nx5667,nx5667,
                       nx5667,nx5667,nx5667,nx5669,nx5669,nx5669,nx5669,nx5669,
                       nx5669,nx5669,nx5671,nx5671,nx5671,nx5671,nx5671,nx5671,
                       nx5671,nx5673,nx5673,nx5673,nx5673,nx5673,nx5673,nx5673,
                       nx5675,nx5675,nx5675,nx5675,nx5675,nx5675,nx5675,nx5677,
                       nx5677,nx5677,nx5677,nx5677,nx5677,nx5677,nx5679,nx5679,
                       nx5679,nx5679,nx5679,nx5679,nx5679,nx5681,nx5681,nx5681,
                       nx5681,nx5681,nx5681,nx5681,nx5683,nx5683,nx5683,nx5683,
                       nx5683,nx5683,nx5683,nx5685,nx5685,nx5685,nx5685,nx5685,
                       nx5685,nx5685,nx5687,nx5687,nx5687,nx5687,nx5687,nx5687,
                       nx5687,nx5689,nx5689,nx5689,nx5689,nx5689,nx5689,nx5689,
                       nx5691,nx5691,nx5691,nx5691,nx5691,nx5691,nx5691,nx5693,
                       nx5693,nx5693,nx5693,nx5693,nx5693,nx5693,nx5695,nx5695,
                       nx5695,nx5695,nx5695,nx5695,nx5695,nx5697,nx5697,nx5697,
                       nx5697,nx5697,nx5697,nx5697,nx5699,nx5699,nx5699,nx5699,
                       nx5699,nx5699,nx5699,nx5701,nx5701,nx5701,nx5701,nx5701,
                       nx5701,nx5701,nx5703,nx5703,nx5703,nx5703,nx5703,nx5703,
                       nx5703,nx5705,nx5705,nx5705,nx5705,nx5705,nx5705,nx5705,
                       nx5707,nx5707,nx5707,nx5707,nx5707,nx5707,nx5707,nx5709,
                       nx5709,nx5709,nx5709,nx5709,nx5709,nx5709,nx5711,nx5711,
                       nx5711,nx5711,nx5711,nx5711,nx5711,nx5713,nx5713,nx5713,
                       nx5713,nx5713,nx5713,nx5713,nx5715,nx5715,nx5715,nx5715,
                       nx5715,nx5715,nx5715,nx5717,nx5717,nx5717,nx5717,nx5717,
                       nx5717,nx5717,nx5719,nx5719,nx5719,nx5719,nx5719,nx5719,
                       nx5719,nx5721,nx5721,nx5721,nx5721,nx5721,nx5721,nx5721,
                       nx5723,nx5723,nx5723,nx5723,nx5723,nx5723,nx5723,nx5725,
                       nx5725,nx5725,nx5725,nx5725,nx5725,nx5725,nx5727,nx5727,
                       nx5727,nx5727,nx5727,nx5727,nx5727,nx5729,nx5729,nx5729,
                       nx5729,nx5729,nx5729,nx5729,nx5731,nx5731,nx5731,nx5731,
                       nx5731,nx5731,nx5731,nx5733,nx5733,nx5733,nx5733,nx5733,
                       nx5733,nx5733,nx5735,nx5735,nx5735,nx5735,nx5735,nx5735,
                       nx5735,nx5737,nx5737,nx5737,nx5737,nx5737,nx5737,nx5737,
                       nx5739,nx5739,nx5739,nx5739,nx5739,nx5739,nx5739,nx5741,
                       nx5741,nx5741,nx5741,nx5741,nx5741,nx5741,nx5743,nx5743,
                       nx5743,nx5743,nx5743,nx5743,nx5743,nx5745,nx5745,nx5745,
                       nx5745,nx5745,nx5745,nx5745,nx5747,nx5747,nx5747,nx5747,
                       nx5747,nx5747,nx5747,nx5749,nx5749,nx5749,nx5749,nx5749,
                       nx5749,nx5749,nx5751,nx5751,nx5751,nx5751,nx5751,nx5751,
                       nx5751,nx5753,nx5753,nx5753,nx5753,nx5753,nx5753,nx5753,
                       nx5755,nx5755,nx5755,nx5755,nx5755,nx5755,nx5755,nx5757,
                       nx5757,nx5757,nx5757,nx5757,nx5757,nx5757,nx5759,nx5759,
                       nx5759,nx5759,nx5759,nx5759,nx5759,nx5761,nx5761,nx5761,
                       nx5761,nx5761,nx5761,nx5761,nx5763,nx5763,nx5763,nx5763,
                       nx5763,nx5763,nx5763,nx5765,nx5765,nx5765,nx5765,nx5765,
                       nx5765,nx5765,nx5767,nx5767,nx5767,nx5767,nx5767,nx5767,
                       nx5767,nx5769,nx5769,nx5769,nx5769,nx5769,nx5769,nx5769,
                       nx5771,nx5771,nx5771,nx5771,nx5771,nx5771,nx5771,nx5773,
                       nx5773,nx5773,nx5773,nx5773,nx5773,nx5773,nx5775,nx5775,
                       nx5775,nx5775,nx5775,nx5775,nx5775,nx5777,nx5777,nx5777,
                       nx5777,nx5777,nx5777,nx5777,nx5779,nx5779,nx5779,nx5779,
                       nx5779,nx5779,nx5779,nx5781,nx5781,nx5781,nx5781,nx5781,
                       nx5781,nx5781}), .EN (test), .F ({dataOut[447],
                       dataOut[446],dataOut[445],dataOut[444],dataOut[443],
                       dataOut[442],dataOut[441],dataOut[440],dataOut[439],
                       dataOut[438],dataOut[437],dataOut[436],dataOut[435],
                       dataOut[434],dataOut[433],dataOut[432],dataOut[431],
                       dataOut[430],dataOut[429],dataOut[428],dataOut[427],
                       dataOut[426],dataOut[425],dataOut[424],dataOut[423],
                       dataOut[422],dataOut[421],dataOut[420],dataOut[419],
                       dataOut[418],dataOut[417],dataOut[416],dataOut[415],
                       dataOut[414],dataOut[413],dataOut[412],dataOut[411],
                       dataOut[410],dataOut[409],dataOut[408],dataOut[407],
                       dataOut[406],dataOut[405],dataOut[404],dataOut[403],
                       dataOut[402],dataOut[401],dataOut[400],dataOut[399],
                       dataOut[398],dataOut[397],dataOut[396],dataOut[395],
                       dataOut[394],dataOut[393],dataOut[392],dataOut[391],
                       dataOut[390],dataOut[389],dataOut[388],dataOut[387],
                       dataOut[386],dataOut[385],dataOut[384],dataOut[383],
                       dataOut[382],dataOut[381],dataOut[380],dataOut[379],
                       dataOut[378],dataOut[377],dataOut[376],dataOut[375],
                       dataOut[374],dataOut[373],dataOut[372],dataOut[371],
                       dataOut[370],dataOut[369],dataOut[368],dataOut[367],
                       dataOut[366],dataOut[365],dataOut[364],dataOut[363],
                       dataOut[362],dataOut[361],dataOut[360],dataOut[359],
                       dataOut[358],dataOut[357],dataOut[356],dataOut[355],
                       dataOut[354],dataOut[353],dataOut[352],dataOut[351],
                       dataOut[350],dataOut[349],dataOut[348],dataOut[347],
                       dataOut[346],dataOut[345],dataOut[344],dataOut[343],
                       dataOut[342],dataOut[341],dataOut[340],dataOut[339],
                       dataOut[338],dataOut[337],dataOut[336],dataOut[335],
                       dataOut[334],dataOut[333],dataOut[332],dataOut[331],
                       dataOut[330],dataOut[329],dataOut[328],dataOut[327],
                       dataOut[326],dataOut[325],dataOut[324],dataOut[323],
                       dataOut[322],dataOut[321],dataOut[320],dataOut[319],
                       dataOut[318],dataOut[317],dataOut[316],dataOut[315],
                       dataOut[314],dataOut[313],dataOut[312],dataOut[311],
                       dataOut[310],dataOut[309],dataOut[308],dataOut[307],
                       dataOut[306],dataOut[305],dataOut[304],dataOut[303],
                       dataOut[302],dataOut[301],dataOut[300],dataOut[299],
                       dataOut[298],dataOut[297],dataOut[296],dataOut[295],
                       dataOut[294],dataOut[293],dataOut[292],dataOut[291],
                       dataOut[290],dataOut[289],dataOut[288],dataOut[287],
                       dataOut[286],dataOut[285],dataOut[284],dataOut[283],
                       dataOut[282],dataOut[281],dataOut[280],dataOut[279],
                       dataOut[278],dataOut[277],dataOut[276],dataOut[275],
                       dataOut[274],dataOut[273],dataOut[272],dataOut[271],
                       dataOut[270],dataOut[269],dataOut[268],dataOut[267],
                       dataOut[266],dataOut[265],dataOut[264],dataOut[263],
                       dataOut[262],dataOut[261],dataOut[260],dataOut[259],
                       dataOut[258],dataOut[257],dataOut[256],dataOut[255],
                       dataOut[254],dataOut[253],dataOut[252],dataOut[251],
                       dataOut[250],dataOut[249],dataOut[248],dataOut[247],
                       dataOut[246],dataOut[245],dataOut[244],dataOut[243],
                       dataOut[242],dataOut[241],dataOut[240],dataOut[239],
                       dataOut[238],dataOut[237],dataOut[236],dataOut[235],
                       dataOut[234],dataOut[233],dataOut[232],dataOut[231],
                       dataOut[230],dataOut[229],dataOut[228],dataOut[227],
                       dataOut[226],dataOut[225],dataOut[224],dataOut[223],
                       dataOut[222],dataOut[221],dataOut[220],dataOut[219],
                       dataOut[218],dataOut[217],dataOut[216],dataOut[215],
                       dataOut[214],dataOut[213],dataOut[212],dataOut[211],
                       dataOut[210],dataOut[209],dataOut[208],dataOut[207],
                       dataOut[206],dataOut[205],dataOut[204],dataOut[203],
                       dataOut[202],dataOut[201],dataOut[200],dataOut[199],
                       dataOut[198],dataOut[197],dataOut[196],dataOut[195],
                       dataOut[194],dataOut[193],dataOut[192],dataOut[191],
                       dataOut[190],dataOut[189],dataOut[188],dataOut[187],
                       dataOut[186],dataOut[185],dataOut[184],dataOut[183],
                       dataOut[182],dataOut[181],dataOut[180],dataOut[179],
                       dataOut[178],dataOut[177],dataOut[176],dataOut[175],
                       dataOut[174],dataOut[173],dataOut[172],dataOut[171],
                       dataOut[170],dataOut[169],dataOut[168],dataOut[167],
                       dataOut[166],dataOut[165],dataOut[164],dataOut[163],
                       dataOut[162],dataOut[161],dataOut[160],dataOut[159],
                       dataOut[158],dataOut[157],dataOut[156],dataOut[155],
                       dataOut[154],dataOut[153],dataOut[152],dataOut[151],
                       dataOut[150],dataOut[149],dataOut[148],dataOut[147],
                       dataOut[146],dataOut[145],dataOut[144],dataOut[143],
                       dataOut[142],dataOut[141],dataOut[140],dataOut[139],
                       dataOut[138],dataOut[137],dataOut[136],dataOut[135],
                       dataOut[134],dataOut[133],dataOut[132],dataOut[131],
                       dataOut[130],dataOut[129],dataOut[128],dataOut[127],
                       dataOut[126],dataOut[125],dataOut[124],dataOut[123],
                       dataOut[122],dataOut[121],dataOut[120],dataOut[119],
                       dataOut[118],dataOut[117],dataOut[116],dataOut[115],
                       dataOut[114],dataOut[113],dataOut[112],dataOut[111],
                       dataOut[110],dataOut[109],dataOut[108],dataOut[107],
                       dataOut[106],dataOut[105],dataOut[104],dataOut[103],
                       dataOut[102],dataOut[101],dataOut[100],dataOut[99],
                       dataOut[98],dataOut[97],dataOut[96],dataOut[95],
                       dataOut[94],dataOut[93],dataOut[92],dataOut[91],
                       dataOut[90],dataOut[89],dataOut[88],dataOut[87],
                       dataOut[86],dataOut[85],dataOut[84],dataOut[83],
                       dataOut[82],dataOut[81],dataOut[80],dataOut[79],
                       dataOut[78],dataOut[77],dataOut[76],dataOut[75],
                       dataOut[74],dataOut[73],dataOut[72],dataOut[71],
                       dataOut[70],dataOut[69],dataOut[68],dataOut[67],
                       dataOut[66],dataOut[65],dataOut[64],dataOut[63],
                       dataOut[62],dataOut[61],dataOut[60],dataOut[59],
                       dataOut[58],dataOut[57],dataOut[56],dataOut[55],
                       dataOut[54],dataOut[53],dataOut[52],dataOut[51],
                       dataOut[50],dataOut[49],dataOut[48],dataOut[47],
                       dataOut[46],dataOut[45],dataOut[44],dataOut[43],
                       dataOut[42],dataOut[41],dataOut[40],dataOut[39],
                       dataOut[38],dataOut[37],dataOut[36],dataOut[35],
                       dataOut[34],dataOut[33],dataOut[32],dataOut[31],
                       dataOut[30],dataOut[29],dataOut[28],dataOut[27],
                       dataOut[26],dataOut[25],dataOut[24],dataOut[23],
                       dataOut[22],dataOut[21],dataOut[20],dataOut[19],
                       dataOut[18],dataOut[17],dataOut[16],dataOut[15],
                       dataOut[14],dataOut[13],dataOut[12],dataOut[11],
                       dataOut[10],dataOut[9],dataOut[8],dataOut[7],dataOut[6],
                       dataOut[5],dataOut[4],dataOut[3],dataOut[2],dataOut[1],
                       dataOut[0]})) ;
    triStateBuffer_16 Ram1Wr (.D ({dataIn[15],dataIn[14],dataIn[13],dataIn[12],
                      dataIn[11],dataIn[10],dataIn[9],dataIn[8],dataIn[7],
                      dataIn[6],dataIn[5],dataIn[4],dataIn[3],dataIn[2],
                      dataIn[1],dataIn[0]}), .EN (ram1Write), .F ({dataToRam1_15
                      ,dataToRam1_14,dataToRam1_13,dataToRam1_12,dataToRam1_11,
                      dataToRam1_10,dataToRam1_9,dataToRam1_8,dataToRam1_7,
                      dataToRam1_6,dataToRam1_5,dataToRam1_4,dataToRam1_3,
                      dataToRam1_2,dataToRam1_1,dataToRam1_0})) ;
    triStateBuffer_448 Ram2Rd (.D ({nx5785,nx5785,nx5785,nx5785,nx5785,nx5785,
                       nx5785,nx5787,nx5787,nx5787,nx5787,nx5787,nx5787,nx5787,
                       nx5789,nx5789,nx5789,nx5789,nx5789,nx5789,nx5789,nx5791,
                       nx5791,nx5791,nx5791,nx5791,nx5791,nx5791,nx5793,nx5793,
                       nx5793,nx5793,nx5793,nx5793,nx5793,nx5795,nx5795,nx5795,
                       nx5795,nx5795,nx5795,nx5795,nx5797,nx5797,nx5797,nx5797,
                       nx5797,nx5797,nx5797,nx5799,nx5799,nx5799,nx5799,nx5799,
                       nx5799,nx5799,nx5801,nx5801,nx5801,nx5801,nx5801,nx5801,
                       nx5801,nx5803,nx5803,nx5803,nx5803,nx5803,nx5803,nx5803,
                       nx5805,nx5805,nx5805,nx5805,nx5805,nx5805,nx5805,nx5807,
                       nx5807,nx5807,nx5807,nx5807,nx5807,nx5807,nx5809,nx5809,
                       nx5809,nx5809,nx5809,nx5809,nx5809,nx5811,nx5811,nx5811,
                       nx5811,nx5811,nx5811,nx5811,nx5813,nx5813,nx5813,nx5813,
                       nx5813,nx5813,nx5813,nx5815,nx5815,nx5815,nx5815,nx5815,
                       nx5815,nx5815,nx5817,nx5817,nx5817,nx5817,nx5817,nx5817,
                       nx5817,nx5819,nx5819,nx5819,nx5819,nx5819,nx5819,nx5819,
                       nx5821,nx5821,nx5821,nx5821,nx5821,nx5821,nx5821,nx5823,
                       nx5823,nx5823,nx5823,nx5823,nx5823,nx5823,nx5825,nx5825,
                       nx5825,nx5825,nx5825,nx5825,nx5825,nx5827,nx5827,nx5827,
                       nx5827,nx5827,nx5827,nx5827,nx5829,nx5829,nx5829,nx5829,
                       nx5829,nx5829,nx5829,nx5831,nx5831,nx5831,nx5831,nx5831,
                       nx5831,nx5831,nx5833,nx5833,nx5833,nx5833,nx5833,nx5833,
                       nx5833,nx5835,nx5835,nx5835,nx5835,nx5835,nx5835,nx5835,
                       nx5837,nx5837,nx5837,nx5837,nx5837,nx5837,nx5837,nx5839,
                       nx5839,nx5839,nx5839,nx5839,nx5839,nx5839,nx5841,nx5841,
                       nx5841,nx5841,nx5841,nx5841,nx5841,nx5843,nx5843,nx5843,
                       nx5843,nx5843,nx5843,nx5843,nx5845,nx5845,nx5845,nx5845,
                       nx5845,nx5845,nx5845,nx5847,nx5847,nx5847,nx5847,nx5847,
                       nx5847,nx5847,nx5849,nx5849,nx5849,nx5849,nx5849,nx5849,
                       nx5849,nx5851,nx5851,nx5851,nx5851,nx5851,nx5851,nx5851,
                       nx5853,nx5853,nx5853,nx5853,nx5853,nx5853,nx5853,nx5855,
                       nx5855,nx5855,nx5855,nx5855,nx5855,nx5855,nx5857,nx5857,
                       nx5857,nx5857,nx5857,nx5857,nx5857,nx5859,nx5859,nx5859,
                       nx5859,nx5859,nx5859,nx5859,nx5861,nx5861,nx5861,nx5861,
                       nx5861,nx5861,nx5861,nx5863,nx5863,nx5863,nx5863,nx5863,
                       nx5863,nx5863,nx5865,nx5865,nx5865,nx5865,nx5865,nx5865,
                       nx5865,nx5867,nx5867,nx5867,nx5867,nx5867,nx5867,nx5867,
                       nx5869,nx5869,nx5869,nx5869,nx5869,nx5869,nx5869,nx5871,
                       nx5871,nx5871,nx5871,nx5871,nx5871,nx5871,nx5873,nx5873,
                       nx5873,nx5873,nx5873,nx5873,nx5873,nx5875,nx5875,nx5875,
                       nx5875,nx5875,nx5875,nx5875,nx5877,nx5877,nx5877,nx5877,
                       nx5877,nx5877,nx5877,nx5879,nx5879,nx5879,nx5879,nx5879,
                       nx5879,nx5879,nx5881,nx5881,nx5881,nx5881,nx5881,nx5881,
                       nx5881,nx5883,nx5883,nx5883,nx5883,nx5883,nx5883,nx5883,
                       nx5885,nx5885,nx5885,nx5885,nx5885,nx5885,nx5885,nx5887,
                       nx5887,nx5887,nx5887,nx5887,nx5887,nx5887,nx5889,nx5889,
                       nx5889,nx5889,nx5889,nx5889,nx5889,nx5891,nx5891,nx5891,
                       nx5891,nx5891,nx5891,nx5891,nx5893,nx5893,nx5893,nx5893,
                       nx5893,nx5893,nx5893,nx5895,nx5895,nx5895,nx5895,nx5895,
                       nx5895,nx5895,nx5897,nx5897,nx5897,nx5897,nx5897,nx5897,
                       nx5897,nx5899,nx5899,nx5899,nx5899,nx5899,nx5899,nx5899,
                       nx5901,nx5901,nx5901,nx5901,nx5901,nx5901,nx5901,nx5903,
                       nx5903,nx5903,nx5903,nx5903,nx5903,nx5903,nx5905,nx5905,
                       nx5905,nx5905,nx5905,nx5905,nx5905,nx5907,nx5907,nx5907,
                       nx5907,nx5907,nx5907,nx5907,nx5909,nx5909,nx5909,nx5909,
                       nx5909,nx5909,nx5909,nx5911,nx5911,nx5911,nx5911,nx5911,
                       nx5911,nx5911}), .EN (DInput), .F ({dataOut[447],
                       dataOut[446],dataOut[445],dataOut[444],dataOut[443],
                       dataOut[442],dataOut[441],dataOut[440],dataOut[439],
                       dataOut[438],dataOut[437],dataOut[436],dataOut[435],
                       dataOut[434],dataOut[433],dataOut[432],dataOut[431],
                       dataOut[430],dataOut[429],dataOut[428],dataOut[427],
                       dataOut[426],dataOut[425],dataOut[424],dataOut[423],
                       dataOut[422],dataOut[421],dataOut[420],dataOut[419],
                       dataOut[418],dataOut[417],dataOut[416],dataOut[415],
                       dataOut[414],dataOut[413],dataOut[412],dataOut[411],
                       dataOut[410],dataOut[409],dataOut[408],dataOut[407],
                       dataOut[406],dataOut[405],dataOut[404],dataOut[403],
                       dataOut[402],dataOut[401],dataOut[400],dataOut[399],
                       dataOut[398],dataOut[397],dataOut[396],dataOut[395],
                       dataOut[394],dataOut[393],dataOut[392],dataOut[391],
                       dataOut[390],dataOut[389],dataOut[388],dataOut[387],
                       dataOut[386],dataOut[385],dataOut[384],dataOut[383],
                       dataOut[382],dataOut[381],dataOut[380],dataOut[379],
                       dataOut[378],dataOut[377],dataOut[376],dataOut[375],
                       dataOut[374],dataOut[373],dataOut[372],dataOut[371],
                       dataOut[370],dataOut[369],dataOut[368],dataOut[367],
                       dataOut[366],dataOut[365],dataOut[364],dataOut[363],
                       dataOut[362],dataOut[361],dataOut[360],dataOut[359],
                       dataOut[358],dataOut[357],dataOut[356],dataOut[355],
                       dataOut[354],dataOut[353],dataOut[352],dataOut[351],
                       dataOut[350],dataOut[349],dataOut[348],dataOut[347],
                       dataOut[346],dataOut[345],dataOut[344],dataOut[343],
                       dataOut[342],dataOut[341],dataOut[340],dataOut[339],
                       dataOut[338],dataOut[337],dataOut[336],dataOut[335],
                       dataOut[334],dataOut[333],dataOut[332],dataOut[331],
                       dataOut[330],dataOut[329],dataOut[328],dataOut[327],
                       dataOut[326],dataOut[325],dataOut[324],dataOut[323],
                       dataOut[322],dataOut[321],dataOut[320],dataOut[319],
                       dataOut[318],dataOut[317],dataOut[316],dataOut[315],
                       dataOut[314],dataOut[313],dataOut[312],dataOut[311],
                       dataOut[310],dataOut[309],dataOut[308],dataOut[307],
                       dataOut[306],dataOut[305],dataOut[304],dataOut[303],
                       dataOut[302],dataOut[301],dataOut[300],dataOut[299],
                       dataOut[298],dataOut[297],dataOut[296],dataOut[295],
                       dataOut[294],dataOut[293],dataOut[292],dataOut[291],
                       dataOut[290],dataOut[289],dataOut[288],dataOut[287],
                       dataOut[286],dataOut[285],dataOut[284],dataOut[283],
                       dataOut[282],dataOut[281],dataOut[280],dataOut[279],
                       dataOut[278],dataOut[277],dataOut[276],dataOut[275],
                       dataOut[274],dataOut[273],dataOut[272],dataOut[271],
                       dataOut[270],dataOut[269],dataOut[268],dataOut[267],
                       dataOut[266],dataOut[265],dataOut[264],dataOut[263],
                       dataOut[262],dataOut[261],dataOut[260],dataOut[259],
                       dataOut[258],dataOut[257],dataOut[256],dataOut[255],
                       dataOut[254],dataOut[253],dataOut[252],dataOut[251],
                       dataOut[250],dataOut[249],dataOut[248],dataOut[247],
                       dataOut[246],dataOut[245],dataOut[244],dataOut[243],
                       dataOut[242],dataOut[241],dataOut[240],dataOut[239],
                       dataOut[238],dataOut[237],dataOut[236],dataOut[235],
                       dataOut[234],dataOut[233],dataOut[232],dataOut[231],
                       dataOut[230],dataOut[229],dataOut[228],dataOut[227],
                       dataOut[226],dataOut[225],dataOut[224],dataOut[223],
                       dataOut[222],dataOut[221],dataOut[220],dataOut[219],
                       dataOut[218],dataOut[217],dataOut[216],dataOut[215],
                       dataOut[214],dataOut[213],dataOut[212],dataOut[211],
                       dataOut[210],dataOut[209],dataOut[208],dataOut[207],
                       dataOut[206],dataOut[205],dataOut[204],dataOut[203],
                       dataOut[202],dataOut[201],dataOut[200],dataOut[199],
                       dataOut[198],dataOut[197],dataOut[196],dataOut[195],
                       dataOut[194],dataOut[193],dataOut[192],dataOut[191],
                       dataOut[190],dataOut[189],dataOut[188],dataOut[187],
                       dataOut[186],dataOut[185],dataOut[184],dataOut[183],
                       dataOut[182],dataOut[181],dataOut[180],dataOut[179],
                       dataOut[178],dataOut[177],dataOut[176],dataOut[175],
                       dataOut[174],dataOut[173],dataOut[172],dataOut[171],
                       dataOut[170],dataOut[169],dataOut[168],dataOut[167],
                       dataOut[166],dataOut[165],dataOut[164],dataOut[163],
                       dataOut[162],dataOut[161],dataOut[160],dataOut[159],
                       dataOut[158],dataOut[157],dataOut[156],dataOut[155],
                       dataOut[154],dataOut[153],dataOut[152],dataOut[151],
                       dataOut[150],dataOut[149],dataOut[148],dataOut[147],
                       dataOut[146],dataOut[145],dataOut[144],dataOut[143],
                       dataOut[142],dataOut[141],dataOut[140],dataOut[139],
                       dataOut[138],dataOut[137],dataOut[136],dataOut[135],
                       dataOut[134],dataOut[133],dataOut[132],dataOut[131],
                       dataOut[130],dataOut[129],dataOut[128],dataOut[127],
                       dataOut[126],dataOut[125],dataOut[124],dataOut[123],
                       dataOut[122],dataOut[121],dataOut[120],dataOut[119],
                       dataOut[118],dataOut[117],dataOut[116],dataOut[115],
                       dataOut[114],dataOut[113],dataOut[112],dataOut[111],
                       dataOut[110],dataOut[109],dataOut[108],dataOut[107],
                       dataOut[106],dataOut[105],dataOut[104],dataOut[103],
                       dataOut[102],dataOut[101],dataOut[100],dataOut[99],
                       dataOut[98],dataOut[97],dataOut[96],dataOut[95],
                       dataOut[94],dataOut[93],dataOut[92],dataOut[91],
                       dataOut[90],dataOut[89],dataOut[88],dataOut[87],
                       dataOut[86],dataOut[85],dataOut[84],dataOut[83],
                       dataOut[82],dataOut[81],dataOut[80],dataOut[79],
                       dataOut[78],dataOut[77],dataOut[76],dataOut[75],
                       dataOut[74],dataOut[73],dataOut[72],dataOut[71],
                       dataOut[70],dataOut[69],dataOut[68],dataOut[67],
                       dataOut[66],dataOut[65],dataOut[64],dataOut[63],
                       dataOut[62],dataOut[61],dataOut[60],dataOut[59],
                       dataOut[58],dataOut[57],dataOut[56],dataOut[55],
                       dataOut[54],dataOut[53],dataOut[52],dataOut[51],
                       dataOut[50],dataOut[49],dataOut[48],dataOut[47],
                       dataOut[46],dataOut[45],dataOut[44],dataOut[43],
                       dataOut[42],dataOut[41],dataOut[40],dataOut[39],
                       dataOut[38],dataOut[37],dataOut[36],dataOut[35],
                       dataOut[34],dataOut[33],dataOut[32],dataOut[31],
                       dataOut[30],dataOut[29],dataOut[28],dataOut[27],
                       dataOut[26],dataOut[25],dataOut[24],dataOut[23],
                       dataOut[22],dataOut[21],dataOut[20],dataOut[19],
                       dataOut[18],dataOut[17],dataOut[16],dataOut[15],
                       dataOut[14],dataOut[13],dataOut[12],dataOut[11],
                       dataOut[10],dataOut[9],dataOut[8],dataOut[7],dataOut[6],
                       dataOut[5],dataOut[4],dataOut[3],dataOut[2],dataOut[1],
                       dataOut[0]})) ;
    triStateBuffer_16 Ram2Wr (.D ({dataIn[15],dataIn[14],dataIn[13],dataIn[12],
                      dataIn[11],dataIn[10],dataIn[9],dataIn[8],dataIn[7],
                      dataIn[6],dataIn[5],dataIn[4],dataIn[3],dataIn[2],
                      dataIn[1],dataIn[0]}), .EN (ram2Write), .F ({dataToRam2_15
                      ,dataToRam2_14,dataToRam2_13,dataToRam2_12,dataToRam2_11,
                      dataToRam2_10,dataToRam2_9,dataToRam2_8,dataToRam2_7,
                      dataToRam2_6,dataToRam2_5,dataToRam2_4,dataToRam2_3,
                      dataToRam2_2,dataToRam2_1,dataToRam2_0})) ;
    RAM_28 Ram1 (.reset (resetEN), .CLK (CLK), .W (ram1Write), .R (ram1Read), .address (
           {AddressIn[12],AddressIn[11],AddressIn[10],AddressIn[9],AddressIn[8],
           AddressIn[7],AddressIn[6],AddressIn[5],AddressIn[4],AddressIn[3],
           AddressIn[2],AddressIn[1],AddressIn[0]}), .dataIn ({dataToRam1_15,
           dataToRam1_14,dataToRam1_13,dataToRam1_12,dataToRam1_11,dataToRam1_10
           ,dataToRam1_9,dataToRam1_8,dataToRam1_7,dataToRam1_6,dataToRam1_5,
           dataToRam1_4,dataToRam1_3,dataToRam1_2,dataToRam1_1,dataToRam1_0}), .dataOut (
           {dataFromRam1_447,\$dummy [0],\$dummy [1],\$dummy [2],\$dummy [3],
           \$dummy [4],\$dummy [5],\$dummy [6],\$dummy [7],\$dummy [8],
           \$dummy [9],\$dummy [10],\$dummy [11],\$dummy [12],\$dummy [13],
           \$dummy [14],\$dummy [15],\$dummy [16],\$dummy [17],\$dummy [18],
           \$dummy [19],\$dummy [20],\$dummy [21],\$dummy [22],\$dummy [23],
           \$dummy [24],\$dummy [25],\$dummy [26],\$dummy [27],\$dummy [28],
           \$dummy [29],\$dummy [30],\$dummy [31],\$dummy [32],\$dummy [33],
           \$dummy [34],\$dummy [35],\$dummy [36],\$dummy [37],\$dummy [38],
           \$dummy [39],\$dummy [40],\$dummy [41],\$dummy [42],\$dummy [43],
           \$dummy [44],\$dummy [45],\$dummy [46],\$dummy [47],\$dummy [48],
           \$dummy [49],\$dummy [50],\$dummy [51],\$dummy [52],\$dummy [53],
           \$dummy [54],\$dummy [55],\$dummy [56],\$dummy [57],\$dummy [58],
           \$dummy [59],\$dummy [60],\$dummy [61],\$dummy [62],\$dummy [63],
           \$dummy [64],\$dummy [65],\$dummy [66],\$dummy [67],\$dummy [68],
           \$dummy [69],\$dummy [70],\$dummy [71],\$dummy [72],\$dummy [73],
           \$dummy [74],\$dummy [75],\$dummy [76],\$dummy [77],\$dummy [78],
           \$dummy [79],\$dummy [80],\$dummy [81],\$dummy [82],\$dummy [83],
           \$dummy [84],\$dummy [85],\$dummy [86],\$dummy [87],\$dummy [88],
           \$dummy [89],\$dummy [90],\$dummy [91],\$dummy [92],\$dummy [93],
           \$dummy [94],\$dummy [95],\$dummy [96],\$dummy [97],\$dummy [98],
           \$dummy [99],\$dummy [100],\$dummy [101],\$dummy [102],\$dummy [103],
           \$dummy [104],\$dummy [105],\$dummy [106],\$dummy [107],\$dummy [108]
           ,\$dummy [109],\$dummy [110],\$dummy [111],\$dummy [112],
           \$dummy [113],\$dummy [114],\$dummy [115],\$dummy [116],\$dummy [117]
           ,\$dummy [118],\$dummy [119],\$dummy [120],\$dummy [121],
           \$dummy [122],\$dummy [123],\$dummy [124],\$dummy [125],\$dummy [126]
           ,\$dummy [127],\$dummy [128],\$dummy [129],\$dummy [130],
           \$dummy [131],\$dummy [132],\$dummy [133],\$dummy [134],\$dummy [135]
           ,\$dummy [136],\$dummy [137],\$dummy [138],\$dummy [139],
           \$dummy [140],\$dummy [141],\$dummy [142],\$dummy [143],\$dummy [144]
           ,\$dummy [145],\$dummy [146],\$dummy [147],\$dummy [148],
           \$dummy [149],\$dummy [150],\$dummy [151],\$dummy [152],\$dummy [153]
           ,\$dummy [154],\$dummy [155],\$dummy [156],\$dummy [157],
           \$dummy [158],\$dummy [159],\$dummy [160],\$dummy [161],\$dummy [162]
           ,\$dummy [163],\$dummy [164],\$dummy [165],\$dummy [166],
           \$dummy [167],\$dummy [168],\$dummy [169],\$dummy [170],\$dummy [171]
           ,\$dummy [172],\$dummy [173],\$dummy [174],\$dummy [175],
           \$dummy [176],\$dummy [177],\$dummy [178],\$dummy [179],\$dummy [180]
           ,\$dummy [181],\$dummy [182],\$dummy [183],\$dummy [184],
           \$dummy [185],\$dummy [186],\$dummy [187],\$dummy [188],\$dummy [189]
           ,\$dummy [190],\$dummy [191],\$dummy [192],\$dummy [193],
           \$dummy [194],\$dummy [195],\$dummy [196],\$dummy [197],\$dummy [198]
           ,\$dummy [199],\$dummy [200],\$dummy [201],\$dummy [202],
           \$dummy [203],\$dummy [204],\$dummy [205],\$dummy [206],\$dummy [207]
           ,\$dummy [208],\$dummy [209],\$dummy [210],\$dummy [211],
           \$dummy [212],\$dummy [213],\$dummy [214],\$dummy [215],\$dummy [216]
           ,\$dummy [217],\$dummy [218],\$dummy [219],\$dummy [220],
           \$dummy [221],\$dummy [222],\$dummy [223],\$dummy [224],\$dummy [225]
           ,\$dummy [226],\$dummy [227],\$dummy [228],\$dummy [229],
           \$dummy [230],\$dummy [231],\$dummy [232],\$dummy [233],\$dummy [234]
           ,\$dummy [235],\$dummy [236],\$dummy [237],\$dummy [238],
           \$dummy [239],\$dummy [240],\$dummy [241],\$dummy [242],\$dummy [243]
           ,\$dummy [244],\$dummy [245],\$dummy [246],\$dummy [247],
           \$dummy [248],\$dummy [249],\$dummy [250],\$dummy [251],\$dummy [252]
           ,\$dummy [253],\$dummy [254],\$dummy [255],\$dummy [256],
           \$dummy [257],\$dummy [258],\$dummy [259],\$dummy [260],\$dummy [261]
           ,\$dummy [262],\$dummy [263],\$dummy [264],\$dummy [265],
           \$dummy [266],\$dummy [267],\$dummy [268],\$dummy [269],\$dummy [270]
           ,\$dummy [271],\$dummy [272],\$dummy [273],\$dummy [274],
           \$dummy [275],\$dummy [276],\$dummy [277],\$dummy [278],\$dummy [279]
           ,\$dummy [280],\$dummy [281],\$dummy [282],\$dummy [283],
           \$dummy [284],\$dummy [285],\$dummy [286],\$dummy [287],\$dummy [288]
           ,\$dummy [289],\$dummy [290],\$dummy [291],\$dummy [292],
           \$dummy [293],\$dummy [294],\$dummy [295],\$dummy [296],\$dummy [297]
           ,\$dummy [298],\$dummy [299],\$dummy [300],\$dummy [301],
           \$dummy [302],\$dummy [303],\$dummy [304],\$dummy [305],\$dummy [306]
           ,\$dummy [307],\$dummy [308],\$dummy [309],\$dummy [310],
           \$dummy [311],\$dummy [312],\$dummy [313],\$dummy [314],\$dummy [315]
           ,\$dummy [316],\$dummy [317],\$dummy [318],\$dummy [319],
           \$dummy [320],\$dummy [321],\$dummy [322],\$dummy [323],\$dummy [324]
           ,\$dummy [325],\$dummy [326],\$dummy [327],\$dummy [328],
           \$dummy [329],\$dummy [330],\$dummy [331],\$dummy [332],\$dummy [333]
           ,\$dummy [334],\$dummy [335],\$dummy [336],\$dummy [337],
           \$dummy [338],\$dummy [339],\$dummy [340],\$dummy [341],\$dummy [342]
           ,\$dummy [343],\$dummy [344],\$dummy [345],\$dummy [346],
           \$dummy [347],\$dummy [348],\$dummy [349],\$dummy [350],\$dummy [351]
           ,\$dummy [352],\$dummy [353],\$dummy [354],\$dummy [355],
           \$dummy [356],\$dummy [357],\$dummy [358],\$dummy [359],\$dummy [360]
           ,\$dummy [361],\$dummy [362],\$dummy [363],\$dummy [364],
           \$dummy [365],\$dummy [366],\$dummy [367],\$dummy [368],\$dummy [369]
           ,\$dummy [370],\$dummy [371],\$dummy [372],\$dummy [373],
           \$dummy [374],\$dummy [375],\$dummy [376],\$dummy [377],\$dummy [378]
           ,\$dummy [379],\$dummy [380],\$dummy [381],\$dummy [382],
           \$dummy [383],\$dummy [384],\$dummy [385],\$dummy [386],\$dummy [387]
           ,\$dummy [388],\$dummy [389],\$dummy [390],\$dummy [391],
           \$dummy [392],\$dummy [393],\$dummy [394],\$dummy [395],\$dummy [396]
           ,\$dummy [397],\$dummy [398],\$dummy [399],\$dummy [400],
           \$dummy [401],\$dummy [402],\$dummy [403],\$dummy [404],\$dummy [405]
           ,\$dummy [406],\$dummy [407],\$dummy [408],\$dummy [409],
           \$dummy [410],\$dummy [411],\$dummy [412],\$dummy [413],\$dummy [414]
           ,\$dummy [415],\$dummy [416],\$dummy [417],\$dummy [418],
           \$dummy [419],\$dummy [420],\$dummy [421],\$dummy [422],\$dummy [423]
           ,\$dummy [424],\$dummy [425],\$dummy [426],\$dummy [427],
           \$dummy [428],\$dummy [429],\$dummy [430],\$dummy [431],\$dummy [432]
           ,\$dummy [433],\$dummy [434],\$dummy [435],\$dummy [436],
           \$dummy [437],\$dummy [438],\$dummy [439],\$dummy [440],\$dummy [441]
           ,\$dummy [442],\$dummy [443],\$dummy [444],\$dummy [445],
           \$dummy [446]}), .MFC (mfcOfRam1), .counterOut ({\$dummy [447],
           \$dummy [448],\$dummy [449],\$dummy [450]})) ;
    RAM_28 Ram2 (.reset (resetEN), .CLK (CLK), .W (ram2Write), .R (ram2Read), .address (
           {AddressIn[12],AddressIn[11],AddressIn[10],AddressIn[9],AddressIn[8],
           AddressIn[7],AddressIn[6],AddressIn[5],AddressIn[4],AddressIn[3],
           AddressIn[2],AddressIn[1],AddressIn[0]}), .dataIn ({dataToRam2_15,
           dataToRam2_14,dataToRam2_13,dataToRam2_12,dataToRam2_11,dataToRam2_10
           ,dataToRam2_9,dataToRam2_8,dataToRam2_7,dataToRam2_6,dataToRam2_5,
           dataToRam2_4,dataToRam2_3,dataToRam2_2,dataToRam2_1,dataToRam2_0}), .dataOut (
           {dataFromRam2_447,\$dummy [451],\$dummy [452],\$dummy [453],
           \$dummy [454],\$dummy [455],\$dummy [456],\$dummy [457],\$dummy [458]
           ,\$dummy [459],\$dummy [460],\$dummy [461],\$dummy [462],
           \$dummy [463],\$dummy [464],\$dummy [465],\$dummy [466],\$dummy [467]
           ,\$dummy [468],\$dummy [469],\$dummy [470],\$dummy [471],
           \$dummy [472],\$dummy [473],\$dummy [474],\$dummy [475],\$dummy [476]
           ,\$dummy [477],\$dummy [478],\$dummy [479],\$dummy [480],
           \$dummy [481],\$dummy [482],\$dummy [483],\$dummy [484],\$dummy [485]
           ,\$dummy [486],\$dummy [487],\$dummy [488],\$dummy [489],
           \$dummy [490],\$dummy [491],\$dummy [492],\$dummy [493],\$dummy [494]
           ,\$dummy [495],\$dummy [496],\$dummy [497],\$dummy [498],
           \$dummy [499],\$dummy [500],\$dummy [501],\$dummy [502],\$dummy [503]
           ,\$dummy [504],\$dummy [505],\$dummy [506],\$dummy [507],
           \$dummy [508],\$dummy [509],\$dummy [510],\$dummy [511],\$dummy [512]
           ,\$dummy [513],\$dummy [514],\$dummy [515],\$dummy [516],
           \$dummy [517],\$dummy [518],\$dummy [519],\$dummy [520],\$dummy [521]
           ,\$dummy [522],\$dummy [523],\$dummy [524],\$dummy [525],
           \$dummy [526],\$dummy [527],\$dummy [528],\$dummy [529],\$dummy [530]
           ,\$dummy [531],\$dummy [532],\$dummy [533],\$dummy [534],
           \$dummy [535],\$dummy [536],\$dummy [537],\$dummy [538],\$dummy [539]
           ,\$dummy [540],\$dummy [541],\$dummy [542],\$dummy [543],
           \$dummy [544],\$dummy [545],\$dummy [546],\$dummy [547],\$dummy [548]
           ,\$dummy [549],\$dummy [550],\$dummy [551],\$dummy [552],
           \$dummy [553],\$dummy [554],\$dummy [555],\$dummy [556],\$dummy [557]
           ,\$dummy [558],\$dummy [559],\$dummy [560],\$dummy [561],
           \$dummy [562],\$dummy [563],\$dummy [564],\$dummy [565],\$dummy [566]
           ,\$dummy [567],\$dummy [568],\$dummy [569],\$dummy [570],
           \$dummy [571],\$dummy [572],\$dummy [573],\$dummy [574],\$dummy [575]
           ,\$dummy [576],\$dummy [577],\$dummy [578],\$dummy [579],
           \$dummy [580],\$dummy [581],\$dummy [582],\$dummy [583],\$dummy [584]
           ,\$dummy [585],\$dummy [586],\$dummy [587],\$dummy [588],
           \$dummy [589],\$dummy [590],\$dummy [591],\$dummy [592],\$dummy [593]
           ,\$dummy [594],\$dummy [595],\$dummy [596],\$dummy [597],
           \$dummy [598],\$dummy [599],\$dummy [600],\$dummy [601],\$dummy [602]
           ,\$dummy [603],\$dummy [604],\$dummy [605],\$dummy [606],
           \$dummy [607],\$dummy [608],\$dummy [609],\$dummy [610],\$dummy [611]
           ,\$dummy [612],\$dummy [613],\$dummy [614],\$dummy [615],
           \$dummy [616],\$dummy [617],\$dummy [618],\$dummy [619],\$dummy [620]
           ,\$dummy [621],\$dummy [622],\$dummy [623],\$dummy [624],
           \$dummy [625],\$dummy [626],\$dummy [627],\$dummy [628],\$dummy [629]
           ,\$dummy [630],\$dummy [631],\$dummy [632],\$dummy [633],
           \$dummy [634],\$dummy [635],\$dummy [636],\$dummy [637],\$dummy [638]
           ,\$dummy [639],\$dummy [640],\$dummy [641],\$dummy [642],
           \$dummy [643],\$dummy [644],\$dummy [645],\$dummy [646],\$dummy [647]
           ,\$dummy [648],\$dummy [649],\$dummy [650],\$dummy [651],
           \$dummy [652],\$dummy [653],\$dummy [654],\$dummy [655],\$dummy [656]
           ,\$dummy [657],\$dummy [658],\$dummy [659],\$dummy [660],
           \$dummy [661],\$dummy [662],\$dummy [663],\$dummy [664],\$dummy [665]
           ,\$dummy [666],\$dummy [667],\$dummy [668],\$dummy [669],
           \$dummy [670],\$dummy [671],\$dummy [672],\$dummy [673],\$dummy [674]
           ,\$dummy [675],\$dummy [676],\$dummy [677],\$dummy [678],
           \$dummy [679],\$dummy [680],\$dummy [681],\$dummy [682],\$dummy [683]
           ,\$dummy [684],\$dummy [685],\$dummy [686],\$dummy [687],
           \$dummy [688],\$dummy [689],\$dummy [690],\$dummy [691],\$dummy [692]
           ,\$dummy [693],\$dummy [694],\$dummy [695],\$dummy [696],
           \$dummy [697],\$dummy [698],\$dummy [699],\$dummy [700],\$dummy [701]
           ,\$dummy [702],\$dummy [703],\$dummy [704],\$dummy [705],
           \$dummy [706],\$dummy [707],\$dummy [708],\$dummy [709],\$dummy [710]
           ,\$dummy [711],\$dummy [712],\$dummy [713],\$dummy [714],
           \$dummy [715],\$dummy [716],\$dummy [717],\$dummy [718],\$dummy [719]
           ,\$dummy [720],\$dummy [721],\$dummy [722],\$dummy [723],
           \$dummy [724],\$dummy [725],\$dummy [726],\$dummy [727],\$dummy [728]
           ,\$dummy [729],\$dummy [730],\$dummy [731],\$dummy [732],
           \$dummy [733],\$dummy [734],\$dummy [735],\$dummy [736],\$dummy [737]
           ,\$dummy [738],\$dummy [739],\$dummy [740],\$dummy [741],
           \$dummy [742],\$dummy [743],\$dummy [744],\$dummy [745],\$dummy [746]
           ,\$dummy [747],\$dummy [748],\$dummy [749],\$dummy [750],
           \$dummy [751],\$dummy [752],\$dummy [753],\$dummy [754],\$dummy [755]
           ,\$dummy [756],\$dummy [757],\$dummy [758],\$dummy [759],
           \$dummy [760],\$dummy [761],\$dummy [762],\$dummy [763],\$dummy [764]
           ,\$dummy [765],\$dummy [766],\$dummy [767],\$dummy [768],
           \$dummy [769],\$dummy [770],\$dummy [771],\$dummy [772],\$dummy [773]
           ,\$dummy [774],\$dummy [775],\$dummy [776],\$dummy [777],
           \$dummy [778],\$dummy [779],\$dummy [780],\$dummy [781],\$dummy [782]
           ,\$dummy [783],\$dummy [784],\$dummy [785],\$dummy [786],
           \$dummy [787],\$dummy [788],\$dummy [789],\$dummy [790],\$dummy [791]
           ,\$dummy [792],\$dummy [793],\$dummy [794],\$dummy [795],
           \$dummy [796],\$dummy [797],\$dummy [798],\$dummy [799],\$dummy [800]
           ,\$dummy [801],\$dummy [802],\$dummy [803],\$dummy [804],
           \$dummy [805],\$dummy [806],\$dummy [807],\$dummy [808],\$dummy [809]
           ,\$dummy [810],\$dummy [811],\$dummy [812],\$dummy [813],
           \$dummy [814],\$dummy [815],\$dummy [816],\$dummy [817],\$dummy [818]
           ,\$dummy [819],\$dummy [820],\$dummy [821],\$dummy [822],
           \$dummy [823],\$dummy [824],\$dummy [825],\$dummy [826],\$dummy [827]
           ,\$dummy [828],\$dummy [829],\$dummy [830],\$dummy [831],
           \$dummy [832],\$dummy [833],\$dummy [834],\$dummy [835],\$dummy [836]
           ,\$dummy [837],\$dummy [838],\$dummy [839],\$dummy [840],
           \$dummy [841],\$dummy [842],\$dummy [843],\$dummy [844],\$dummy [845]
           ,\$dummy [846],\$dummy [847],\$dummy [848],\$dummy [849],
           \$dummy [850],\$dummy [851],\$dummy [852],\$dummy [853],\$dummy [854]
           ,\$dummy [855],\$dummy [856],\$dummy [857],\$dummy [858],
           \$dummy [859],\$dummy [860],\$dummy [861],\$dummy [862],\$dummy [863]
           ,\$dummy [864],\$dummy [865],\$dummy [866],\$dummy [867],
           \$dummy [868],\$dummy [869],\$dummy [870],\$dummy [871],\$dummy [872]
           ,\$dummy [873],\$dummy [874],\$dummy [875],\$dummy [876],
           \$dummy [877],\$dummy [878],\$dummy [879],\$dummy [880],\$dummy [881]
           ,\$dummy [882],\$dummy [883],\$dummy [884],\$dummy [885],
           \$dummy [886],\$dummy [887],\$dummy [888],\$dummy [889],\$dummy [890]
           ,\$dummy [891],\$dummy [892],\$dummy [893],\$dummy [894],
           \$dummy [895],\$dummy [896],\$dummy [897]}), .MFC (mfcOfRam2), .counterOut (
           {\$dummy [898],\$dummy [899],\$dummy [900],\$dummy [901]})) ;
    fake_vcc ix5633 (.Y (nx5632)) ;
    xnor2 ix5636 (.Y (test), .A0 (switcherEN), .A1 (ramSelector)) ;
    fake_gnd ix5623 (.Y (GND)) ;
    tri01 tri_counterOut_0 (.Y (counterOut[0]), .A (nx5632), .E (GND)) ;
    tri01 tri_counterOut_1 (.Y (counterOut[1]), .A (nx5632), .E (GND)) ;
    tri01 tri_counterOut_2 (.Y (counterOut[2]), .A (nx5632), .E (GND)) ;
    tri01 tri_counterOut_3 (.Y (counterOut[3]), .A (nx5632), .E (GND)) ;
    inv01 ix1 (.Y (DInput), .A (test)) ;
    inv01 ix5652 (.Y (nx5653), .A (dataFromRam1_447)) ;
    inv01 ix5654 (.Y (nx5655), .A (nx5913)) ;
    inv01 ix5656 (.Y (nx5657), .A (nx5913)) ;
    inv01 ix5658 (.Y (nx5659), .A (nx5913)) ;
    inv01 ix5660 (.Y (nx5661), .A (nx5913)) ;
    inv01 ix5662 (.Y (nx5663), .A (nx5913)) ;
    inv01 ix5664 (.Y (nx5665), .A (nx5913)) ;
    inv01 ix5666 (.Y (nx5667), .A (nx5913)) ;
    inv01 ix5668 (.Y (nx5669), .A (nx5915)) ;
    inv01 ix5670 (.Y (nx5671), .A (nx5915)) ;
    inv01 ix5672 (.Y (nx5673), .A (nx5915)) ;
    inv01 ix5674 (.Y (nx5675), .A (nx5915)) ;
    inv01 ix5676 (.Y (nx5677), .A (nx5915)) ;
    inv01 ix5678 (.Y (nx5679), .A (nx5915)) ;
    inv01 ix5680 (.Y (nx5681), .A (nx5915)) ;
    inv01 ix5682 (.Y (nx5683), .A (nx5917)) ;
    inv01 ix5684 (.Y (nx5685), .A (nx5917)) ;
    inv01 ix5686 (.Y (nx5687), .A (nx5917)) ;
    inv01 ix5688 (.Y (nx5689), .A (nx5917)) ;
    inv01 ix5690 (.Y (nx5691), .A (nx5917)) ;
    inv01 ix5692 (.Y (nx5693), .A (nx5917)) ;
    inv01 ix5694 (.Y (nx5695), .A (nx5917)) ;
    inv01 ix5696 (.Y (nx5697), .A (nx5919)) ;
    inv01 ix5698 (.Y (nx5699), .A (nx5919)) ;
    inv01 ix5700 (.Y (nx5701), .A (nx5919)) ;
    inv01 ix5702 (.Y (nx5703), .A (nx5919)) ;
    inv01 ix5704 (.Y (nx5705), .A (nx5919)) ;
    inv01 ix5706 (.Y (nx5707), .A (nx5919)) ;
    inv01 ix5708 (.Y (nx5709), .A (nx5919)) ;
    inv01 ix5710 (.Y (nx5711), .A (nx5921)) ;
    inv01 ix5712 (.Y (nx5713), .A (nx5921)) ;
    inv01 ix5714 (.Y (nx5715), .A (nx5921)) ;
    inv01 ix5716 (.Y (nx5717), .A (nx5921)) ;
    inv01 ix5718 (.Y (nx5719), .A (nx5921)) ;
    inv01 ix5720 (.Y (nx5721), .A (nx5921)) ;
    inv01 ix5722 (.Y (nx5723), .A (nx5921)) ;
    inv01 ix5724 (.Y (nx5725), .A (nx5923)) ;
    inv01 ix5726 (.Y (nx5727), .A (nx5923)) ;
    inv01 ix5728 (.Y (nx5729), .A (nx5923)) ;
    inv01 ix5730 (.Y (nx5731), .A (nx5923)) ;
    inv01 ix5732 (.Y (nx5733), .A (nx5923)) ;
    inv01 ix5734 (.Y (nx5735), .A (nx5923)) ;
    inv01 ix5736 (.Y (nx5737), .A (nx5923)) ;
    inv01 ix5738 (.Y (nx5739), .A (nx5925)) ;
    inv01 ix5740 (.Y (nx5741), .A (nx5925)) ;
    inv01 ix5742 (.Y (nx5743), .A (nx5925)) ;
    inv01 ix5744 (.Y (nx5745), .A (nx5925)) ;
    inv01 ix5746 (.Y (nx5747), .A (nx5925)) ;
    inv01 ix5748 (.Y (nx5749), .A (nx5925)) ;
    inv01 ix5750 (.Y (nx5751), .A (nx5925)) ;
    inv01 ix5752 (.Y (nx5753), .A (nx5927)) ;
    inv01 ix5754 (.Y (nx5755), .A (nx5927)) ;
    inv01 ix5756 (.Y (nx5757), .A (nx5927)) ;
    inv01 ix5758 (.Y (nx5759), .A (nx5927)) ;
    inv01 ix5760 (.Y (nx5761), .A (nx5927)) ;
    inv01 ix5762 (.Y (nx5763), .A (nx5927)) ;
    inv01 ix5764 (.Y (nx5765), .A (nx5927)) ;
    inv01 ix5766 (.Y (nx5767), .A (nx5929)) ;
    inv01 ix5768 (.Y (nx5769), .A (nx5929)) ;
    inv01 ix5770 (.Y (nx5771), .A (nx5929)) ;
    inv01 ix5772 (.Y (nx5773), .A (nx5929)) ;
    inv01 ix5774 (.Y (nx5775), .A (nx5929)) ;
    inv01 ix5776 (.Y (nx5777), .A (nx5929)) ;
    inv01 ix5778 (.Y (nx5779), .A (nx5929)) ;
    inv01 ix5780 (.Y (nx5781), .A (nx5653)) ;
    inv01 ix5782 (.Y (nx5783), .A (dataFromRam2_447)) ;
    inv01 ix5784 (.Y (nx5785), .A (nx5931)) ;
    inv01 ix5786 (.Y (nx5787), .A (nx5931)) ;
    inv01 ix5788 (.Y (nx5789), .A (nx5931)) ;
    inv01 ix5790 (.Y (nx5791), .A (nx5931)) ;
    inv01 ix5792 (.Y (nx5793), .A (nx5931)) ;
    inv01 ix5794 (.Y (nx5795), .A (nx5931)) ;
    inv01 ix5796 (.Y (nx5797), .A (nx5931)) ;
    inv01 ix5798 (.Y (nx5799), .A (nx5933)) ;
    inv01 ix5800 (.Y (nx5801), .A (nx5933)) ;
    inv01 ix5802 (.Y (nx5803), .A (nx5933)) ;
    inv01 ix5804 (.Y (nx5805), .A (nx5933)) ;
    inv01 ix5806 (.Y (nx5807), .A (nx5933)) ;
    inv01 ix5808 (.Y (nx5809), .A (nx5933)) ;
    inv01 ix5810 (.Y (nx5811), .A (nx5933)) ;
    inv01 ix5812 (.Y (nx5813), .A (nx5935)) ;
    inv01 ix5814 (.Y (nx5815), .A (nx5935)) ;
    inv01 ix5816 (.Y (nx5817), .A (nx5935)) ;
    inv01 ix5818 (.Y (nx5819), .A (nx5935)) ;
    inv01 ix5820 (.Y (nx5821), .A (nx5935)) ;
    inv01 ix5822 (.Y (nx5823), .A (nx5935)) ;
    inv01 ix5824 (.Y (nx5825), .A (nx5935)) ;
    inv01 ix5826 (.Y (nx5827), .A (nx5937)) ;
    inv01 ix5828 (.Y (nx5829), .A (nx5937)) ;
    inv01 ix5830 (.Y (nx5831), .A (nx5937)) ;
    inv01 ix5832 (.Y (nx5833), .A (nx5937)) ;
    inv01 ix5834 (.Y (nx5835), .A (nx5937)) ;
    inv01 ix5836 (.Y (nx5837), .A (nx5937)) ;
    inv01 ix5838 (.Y (nx5839), .A (nx5937)) ;
    inv01 ix5840 (.Y (nx5841), .A (nx5939)) ;
    inv01 ix5842 (.Y (nx5843), .A (nx5939)) ;
    inv01 ix5844 (.Y (nx5845), .A (nx5939)) ;
    inv01 ix5846 (.Y (nx5847), .A (nx5939)) ;
    inv01 ix5848 (.Y (nx5849), .A (nx5939)) ;
    inv01 ix5850 (.Y (nx5851), .A (nx5939)) ;
    inv01 ix5852 (.Y (nx5853), .A (nx5939)) ;
    inv01 ix5854 (.Y (nx5855), .A (nx5941)) ;
    inv01 ix5856 (.Y (nx5857), .A (nx5941)) ;
    inv01 ix5858 (.Y (nx5859), .A (nx5941)) ;
    inv01 ix5860 (.Y (nx5861), .A (nx5941)) ;
    inv01 ix5862 (.Y (nx5863), .A (nx5941)) ;
    inv01 ix5864 (.Y (nx5865), .A (nx5941)) ;
    inv01 ix5866 (.Y (nx5867), .A (nx5941)) ;
    inv01 ix5868 (.Y (nx5869), .A (nx5943)) ;
    inv01 ix5870 (.Y (nx5871), .A (nx5943)) ;
    inv01 ix5872 (.Y (nx5873), .A (nx5943)) ;
    inv01 ix5874 (.Y (nx5875), .A (nx5943)) ;
    inv01 ix5876 (.Y (nx5877), .A (nx5943)) ;
    inv01 ix5878 (.Y (nx5879), .A (nx5943)) ;
    inv01 ix5880 (.Y (nx5881), .A (nx5943)) ;
    inv01 ix5882 (.Y (nx5883), .A (nx5945)) ;
    inv01 ix5884 (.Y (nx5885), .A (nx5945)) ;
    inv01 ix5886 (.Y (nx5887), .A (nx5945)) ;
    inv01 ix5888 (.Y (nx5889), .A (nx5945)) ;
    inv01 ix5890 (.Y (nx5891), .A (nx5945)) ;
    inv01 ix5892 (.Y (nx5893), .A (nx5945)) ;
    inv01 ix5894 (.Y (nx5895), .A (nx5945)) ;
    inv01 ix5896 (.Y (nx5897), .A (nx5947)) ;
    inv01 ix5898 (.Y (nx5899), .A (nx5947)) ;
    inv01 ix5900 (.Y (nx5901), .A (nx5947)) ;
    inv01 ix5902 (.Y (nx5903), .A (nx5947)) ;
    inv01 ix5904 (.Y (nx5905), .A (nx5947)) ;
    inv01 ix5906 (.Y (nx5907), .A (nx5947)) ;
    inv01 ix5908 (.Y (nx5909), .A (nx5947)) ;
    inv01 ix5910 (.Y (nx5911), .A (nx5783)) ;
    inv01 ix5912 (.Y (nx5913), .A (nx5953)) ;
    inv01 ix5914 (.Y (nx5915), .A (nx5953)) ;
    inv01 ix5916 (.Y (nx5917), .A (nx5953)) ;
    inv01 ix5918 (.Y (nx5919), .A (nx5953)) ;
    inv01 ix5920 (.Y (nx5921), .A (nx5953)) ;
    inv01 ix5922 (.Y (nx5923), .A (nx5953)) ;
    inv01 ix5924 (.Y (nx5925), .A (nx5953)) ;
    inv01 ix5926 (.Y (nx5927), .A (nx5955)) ;
    inv01 ix5928 (.Y (nx5929), .A (nx5955)) ;
    inv01 ix5930 (.Y (nx5931), .A (nx5957)) ;
    inv01 ix5932 (.Y (nx5933), .A (nx5957)) ;
    inv01 ix5934 (.Y (nx5935), .A (nx5957)) ;
    inv01 ix5936 (.Y (nx5937), .A (nx5957)) ;
    inv01 ix5938 (.Y (nx5939), .A (nx5957)) ;
    inv01 ix5940 (.Y (nx5941), .A (nx5957)) ;
    inv01 ix5942 (.Y (nx5943), .A (nx5957)) ;
    inv01 ix5944 (.Y (nx5945), .A (nx5959)) ;
    inv01 ix5946 (.Y (nx5947), .A (nx5959)) ;
    inv01 ix5952 (.Y (nx5953), .A (nx5653)) ;
    inv01 ix5954 (.Y (nx5955), .A (nx5653)) ;
    inv01 ix5956 (.Y (nx5957), .A (nx5783)) ;
    inv01 ix5958 (.Y (nx5959), .A (nx5783)) ;
    and02 ix13 (.Y (ram1Write), .A0 (test), .A1 (writeEn)) ;
    nor02ii ix15 (.Y (ram2Write), .A0 (test), .A1 (writeEn)) ;
    and02 ix19 (.Y (ram1Read), .A0 (test), .A1 (readEn)) ;
    nor02ii ix21 (.Y (ram2Read), .A0 (test), .A1 (readEn)) ;
    mux21_ni ix9 (.Y (MFC), .A0 (mfcOfRam2), .A1 (mfcOfRam1), .S0 (test)) ;
endmodule


module RAM_28 ( reset, CLK, W, R, address, dataIn, dataOut, MFC, counterOut ) ;

    input reset ;
    input CLK ;
    input W ;
    input R ;
    input [12:0]address ;
    input [15:0]dataIn ;
    output [447:0]dataOut ;
    output MFC ;
    output [3:0]counterOut ;

    wire nx12, nx30, nx34, nx42, nx46, nx52, nx98, nx104, nx114, nx116, nx118, 
         nx6871, nx6873, nx6876, nx6881, nx6888, nx6895, nx6897, nx6899, nx6901, 
         nx6903, nx6914, nx1, nx5;



    assign dataOut[447] = dataOut[0] ;
    assign dataOut[446] = dataOut[0] ;
    assign dataOut[445] = dataOut[0] ;
    assign dataOut[444] = dataOut[0] ;
    assign dataOut[443] = dataOut[0] ;
    assign dataOut[442] = dataOut[0] ;
    assign dataOut[441] = dataOut[0] ;
    assign dataOut[440] = dataOut[0] ;
    assign dataOut[439] = dataOut[0] ;
    assign dataOut[438] = dataOut[0] ;
    assign dataOut[437] = dataOut[0] ;
    assign dataOut[436] = dataOut[0] ;
    assign dataOut[435] = dataOut[0] ;
    assign dataOut[434] = dataOut[0] ;
    assign dataOut[433] = dataOut[0] ;
    assign dataOut[432] = dataOut[0] ;
    assign dataOut[431] = dataOut[0] ;
    assign dataOut[430] = dataOut[0] ;
    assign dataOut[429] = dataOut[0] ;
    assign dataOut[428] = dataOut[0] ;
    assign dataOut[427] = dataOut[0] ;
    assign dataOut[426] = dataOut[0] ;
    assign dataOut[425] = dataOut[0] ;
    assign dataOut[424] = dataOut[0] ;
    assign dataOut[423] = dataOut[0] ;
    assign dataOut[422] = dataOut[0] ;
    assign dataOut[421] = dataOut[0] ;
    assign dataOut[420] = dataOut[0] ;
    assign dataOut[419] = dataOut[0] ;
    assign dataOut[418] = dataOut[0] ;
    assign dataOut[417] = dataOut[0] ;
    assign dataOut[416] = dataOut[0] ;
    assign dataOut[415] = dataOut[0] ;
    assign dataOut[414] = dataOut[0] ;
    assign dataOut[413] = dataOut[0] ;
    assign dataOut[412] = dataOut[0] ;
    assign dataOut[411] = dataOut[0] ;
    assign dataOut[410] = dataOut[0] ;
    assign dataOut[409] = dataOut[0] ;
    assign dataOut[408] = dataOut[0] ;
    assign dataOut[407] = dataOut[0] ;
    assign dataOut[406] = dataOut[0] ;
    assign dataOut[405] = dataOut[0] ;
    assign dataOut[404] = dataOut[0] ;
    assign dataOut[403] = dataOut[0] ;
    assign dataOut[402] = dataOut[0] ;
    assign dataOut[401] = dataOut[0] ;
    assign dataOut[400] = dataOut[0] ;
    assign dataOut[399] = dataOut[0] ;
    assign dataOut[398] = dataOut[0] ;
    assign dataOut[397] = dataOut[0] ;
    assign dataOut[396] = dataOut[0] ;
    assign dataOut[395] = dataOut[0] ;
    assign dataOut[394] = dataOut[0] ;
    assign dataOut[393] = dataOut[0] ;
    assign dataOut[392] = dataOut[0] ;
    assign dataOut[391] = dataOut[0] ;
    assign dataOut[390] = dataOut[0] ;
    assign dataOut[389] = dataOut[0] ;
    assign dataOut[388] = dataOut[0] ;
    assign dataOut[387] = dataOut[0] ;
    assign dataOut[386] = dataOut[0] ;
    assign dataOut[385] = dataOut[0] ;
    assign dataOut[384] = dataOut[0] ;
    assign dataOut[383] = dataOut[0] ;
    assign dataOut[382] = dataOut[0] ;
    assign dataOut[381] = dataOut[0] ;
    assign dataOut[380] = dataOut[0] ;
    assign dataOut[379] = dataOut[0] ;
    assign dataOut[378] = dataOut[0] ;
    assign dataOut[377] = dataOut[0] ;
    assign dataOut[376] = dataOut[0] ;
    assign dataOut[375] = dataOut[0] ;
    assign dataOut[374] = dataOut[0] ;
    assign dataOut[373] = dataOut[0] ;
    assign dataOut[372] = dataOut[0] ;
    assign dataOut[371] = dataOut[0] ;
    assign dataOut[370] = dataOut[0] ;
    assign dataOut[369] = dataOut[0] ;
    assign dataOut[368] = dataOut[0] ;
    assign dataOut[367] = dataOut[0] ;
    assign dataOut[366] = dataOut[0] ;
    assign dataOut[365] = dataOut[0] ;
    assign dataOut[364] = dataOut[0] ;
    assign dataOut[363] = dataOut[0] ;
    assign dataOut[362] = dataOut[0] ;
    assign dataOut[361] = dataOut[0] ;
    assign dataOut[360] = dataOut[0] ;
    assign dataOut[359] = dataOut[0] ;
    assign dataOut[358] = dataOut[0] ;
    assign dataOut[357] = dataOut[0] ;
    assign dataOut[356] = dataOut[0] ;
    assign dataOut[355] = dataOut[0] ;
    assign dataOut[354] = dataOut[0] ;
    assign dataOut[353] = dataOut[0] ;
    assign dataOut[352] = dataOut[0] ;
    assign dataOut[351] = dataOut[0] ;
    assign dataOut[350] = dataOut[0] ;
    assign dataOut[349] = dataOut[0] ;
    assign dataOut[348] = dataOut[0] ;
    assign dataOut[347] = dataOut[0] ;
    assign dataOut[346] = dataOut[0] ;
    assign dataOut[345] = dataOut[0] ;
    assign dataOut[344] = dataOut[0] ;
    assign dataOut[343] = dataOut[0] ;
    assign dataOut[342] = dataOut[0] ;
    assign dataOut[341] = dataOut[0] ;
    assign dataOut[340] = dataOut[0] ;
    assign dataOut[339] = dataOut[0] ;
    assign dataOut[338] = dataOut[0] ;
    assign dataOut[337] = dataOut[0] ;
    assign dataOut[336] = dataOut[0] ;
    assign dataOut[335] = dataOut[0] ;
    assign dataOut[334] = dataOut[0] ;
    assign dataOut[333] = dataOut[0] ;
    assign dataOut[332] = dataOut[0] ;
    assign dataOut[331] = dataOut[0] ;
    assign dataOut[330] = dataOut[0] ;
    assign dataOut[329] = dataOut[0] ;
    assign dataOut[328] = dataOut[0] ;
    assign dataOut[327] = dataOut[0] ;
    assign dataOut[326] = dataOut[0] ;
    assign dataOut[325] = dataOut[0] ;
    assign dataOut[324] = dataOut[0] ;
    assign dataOut[323] = dataOut[0] ;
    assign dataOut[322] = dataOut[0] ;
    assign dataOut[321] = dataOut[0] ;
    assign dataOut[320] = dataOut[0] ;
    assign dataOut[319] = dataOut[0] ;
    assign dataOut[318] = dataOut[0] ;
    assign dataOut[317] = dataOut[0] ;
    assign dataOut[316] = dataOut[0] ;
    assign dataOut[315] = dataOut[0] ;
    assign dataOut[314] = dataOut[0] ;
    assign dataOut[313] = dataOut[0] ;
    assign dataOut[312] = dataOut[0] ;
    assign dataOut[311] = dataOut[0] ;
    assign dataOut[310] = dataOut[0] ;
    assign dataOut[309] = dataOut[0] ;
    assign dataOut[308] = dataOut[0] ;
    assign dataOut[307] = dataOut[0] ;
    assign dataOut[306] = dataOut[0] ;
    assign dataOut[305] = dataOut[0] ;
    assign dataOut[304] = dataOut[0] ;
    assign dataOut[303] = dataOut[0] ;
    assign dataOut[302] = dataOut[0] ;
    assign dataOut[301] = dataOut[0] ;
    assign dataOut[300] = dataOut[0] ;
    assign dataOut[299] = dataOut[0] ;
    assign dataOut[298] = dataOut[0] ;
    assign dataOut[297] = dataOut[0] ;
    assign dataOut[296] = dataOut[0] ;
    assign dataOut[295] = dataOut[0] ;
    assign dataOut[294] = dataOut[0] ;
    assign dataOut[293] = dataOut[0] ;
    assign dataOut[292] = dataOut[0] ;
    assign dataOut[291] = dataOut[0] ;
    assign dataOut[290] = dataOut[0] ;
    assign dataOut[289] = dataOut[0] ;
    assign dataOut[288] = dataOut[0] ;
    assign dataOut[287] = dataOut[0] ;
    assign dataOut[286] = dataOut[0] ;
    assign dataOut[285] = dataOut[0] ;
    assign dataOut[284] = dataOut[0] ;
    assign dataOut[283] = dataOut[0] ;
    assign dataOut[282] = dataOut[0] ;
    assign dataOut[281] = dataOut[0] ;
    assign dataOut[280] = dataOut[0] ;
    assign dataOut[279] = dataOut[0] ;
    assign dataOut[278] = dataOut[0] ;
    assign dataOut[277] = dataOut[0] ;
    assign dataOut[276] = dataOut[0] ;
    assign dataOut[275] = dataOut[0] ;
    assign dataOut[274] = dataOut[0] ;
    assign dataOut[273] = dataOut[0] ;
    assign dataOut[272] = dataOut[0] ;
    assign dataOut[271] = dataOut[0] ;
    assign dataOut[270] = dataOut[0] ;
    assign dataOut[269] = dataOut[0] ;
    assign dataOut[268] = dataOut[0] ;
    assign dataOut[267] = dataOut[0] ;
    assign dataOut[266] = dataOut[0] ;
    assign dataOut[265] = dataOut[0] ;
    assign dataOut[264] = dataOut[0] ;
    assign dataOut[263] = dataOut[0] ;
    assign dataOut[262] = dataOut[0] ;
    assign dataOut[261] = dataOut[0] ;
    assign dataOut[260] = dataOut[0] ;
    assign dataOut[259] = dataOut[0] ;
    assign dataOut[258] = dataOut[0] ;
    assign dataOut[257] = dataOut[0] ;
    assign dataOut[256] = dataOut[0] ;
    assign dataOut[255] = dataOut[0] ;
    assign dataOut[254] = dataOut[0] ;
    assign dataOut[253] = dataOut[0] ;
    assign dataOut[252] = dataOut[0] ;
    assign dataOut[251] = dataOut[0] ;
    assign dataOut[250] = dataOut[0] ;
    assign dataOut[249] = dataOut[0] ;
    assign dataOut[248] = dataOut[0] ;
    assign dataOut[247] = dataOut[0] ;
    assign dataOut[246] = dataOut[0] ;
    assign dataOut[245] = dataOut[0] ;
    assign dataOut[244] = dataOut[0] ;
    assign dataOut[243] = dataOut[0] ;
    assign dataOut[242] = dataOut[0] ;
    assign dataOut[241] = dataOut[0] ;
    assign dataOut[240] = dataOut[0] ;
    assign dataOut[239] = dataOut[0] ;
    assign dataOut[238] = dataOut[0] ;
    assign dataOut[237] = dataOut[0] ;
    assign dataOut[236] = dataOut[0] ;
    assign dataOut[235] = dataOut[0] ;
    assign dataOut[234] = dataOut[0] ;
    assign dataOut[233] = dataOut[0] ;
    assign dataOut[232] = dataOut[0] ;
    assign dataOut[231] = dataOut[0] ;
    assign dataOut[230] = dataOut[0] ;
    assign dataOut[229] = dataOut[0] ;
    assign dataOut[228] = dataOut[0] ;
    assign dataOut[227] = dataOut[0] ;
    assign dataOut[226] = dataOut[0] ;
    assign dataOut[225] = dataOut[0] ;
    assign dataOut[224] = dataOut[0] ;
    assign dataOut[223] = dataOut[0] ;
    assign dataOut[222] = dataOut[0] ;
    assign dataOut[221] = dataOut[0] ;
    assign dataOut[220] = dataOut[0] ;
    assign dataOut[219] = dataOut[0] ;
    assign dataOut[218] = dataOut[0] ;
    assign dataOut[217] = dataOut[0] ;
    assign dataOut[216] = dataOut[0] ;
    assign dataOut[215] = dataOut[0] ;
    assign dataOut[214] = dataOut[0] ;
    assign dataOut[213] = dataOut[0] ;
    assign dataOut[212] = dataOut[0] ;
    assign dataOut[211] = dataOut[0] ;
    assign dataOut[210] = dataOut[0] ;
    assign dataOut[209] = dataOut[0] ;
    assign dataOut[208] = dataOut[0] ;
    assign dataOut[207] = dataOut[0] ;
    assign dataOut[206] = dataOut[0] ;
    assign dataOut[205] = dataOut[0] ;
    assign dataOut[204] = dataOut[0] ;
    assign dataOut[203] = dataOut[0] ;
    assign dataOut[202] = dataOut[0] ;
    assign dataOut[201] = dataOut[0] ;
    assign dataOut[200] = dataOut[0] ;
    assign dataOut[199] = dataOut[0] ;
    assign dataOut[198] = dataOut[0] ;
    assign dataOut[197] = dataOut[0] ;
    assign dataOut[196] = dataOut[0] ;
    assign dataOut[195] = dataOut[0] ;
    assign dataOut[194] = dataOut[0] ;
    assign dataOut[193] = dataOut[0] ;
    assign dataOut[192] = dataOut[0] ;
    assign dataOut[191] = dataOut[0] ;
    assign dataOut[190] = dataOut[0] ;
    assign dataOut[189] = dataOut[0] ;
    assign dataOut[188] = dataOut[0] ;
    assign dataOut[187] = dataOut[0] ;
    assign dataOut[186] = dataOut[0] ;
    assign dataOut[185] = dataOut[0] ;
    assign dataOut[184] = dataOut[0] ;
    assign dataOut[183] = dataOut[0] ;
    assign dataOut[182] = dataOut[0] ;
    assign dataOut[181] = dataOut[0] ;
    assign dataOut[180] = dataOut[0] ;
    assign dataOut[179] = dataOut[0] ;
    assign dataOut[178] = dataOut[0] ;
    assign dataOut[177] = dataOut[0] ;
    assign dataOut[176] = dataOut[0] ;
    assign dataOut[175] = dataOut[0] ;
    assign dataOut[174] = dataOut[0] ;
    assign dataOut[173] = dataOut[0] ;
    assign dataOut[172] = dataOut[0] ;
    assign dataOut[171] = dataOut[0] ;
    assign dataOut[170] = dataOut[0] ;
    assign dataOut[169] = dataOut[0] ;
    assign dataOut[168] = dataOut[0] ;
    assign dataOut[167] = dataOut[0] ;
    assign dataOut[166] = dataOut[0] ;
    assign dataOut[165] = dataOut[0] ;
    assign dataOut[164] = dataOut[0] ;
    assign dataOut[163] = dataOut[0] ;
    assign dataOut[162] = dataOut[0] ;
    assign dataOut[161] = dataOut[0] ;
    assign dataOut[160] = dataOut[0] ;
    assign dataOut[159] = dataOut[0] ;
    assign dataOut[158] = dataOut[0] ;
    assign dataOut[157] = dataOut[0] ;
    assign dataOut[156] = dataOut[0] ;
    assign dataOut[155] = dataOut[0] ;
    assign dataOut[154] = dataOut[0] ;
    assign dataOut[153] = dataOut[0] ;
    assign dataOut[152] = dataOut[0] ;
    assign dataOut[151] = dataOut[0] ;
    assign dataOut[150] = dataOut[0] ;
    assign dataOut[149] = dataOut[0] ;
    assign dataOut[148] = dataOut[0] ;
    assign dataOut[147] = dataOut[0] ;
    assign dataOut[146] = dataOut[0] ;
    assign dataOut[145] = dataOut[0] ;
    assign dataOut[144] = dataOut[0] ;
    assign dataOut[143] = dataOut[0] ;
    assign dataOut[142] = dataOut[0] ;
    assign dataOut[141] = dataOut[0] ;
    assign dataOut[140] = dataOut[0] ;
    assign dataOut[139] = dataOut[0] ;
    assign dataOut[138] = dataOut[0] ;
    assign dataOut[137] = dataOut[0] ;
    assign dataOut[136] = dataOut[0] ;
    assign dataOut[135] = dataOut[0] ;
    assign dataOut[134] = dataOut[0] ;
    assign dataOut[133] = dataOut[0] ;
    assign dataOut[132] = dataOut[0] ;
    assign dataOut[131] = dataOut[0] ;
    assign dataOut[130] = dataOut[0] ;
    assign dataOut[129] = dataOut[0] ;
    assign dataOut[128] = dataOut[0] ;
    assign dataOut[127] = dataOut[0] ;
    assign dataOut[126] = dataOut[0] ;
    assign dataOut[125] = dataOut[0] ;
    assign dataOut[124] = dataOut[0] ;
    assign dataOut[123] = dataOut[0] ;
    assign dataOut[122] = dataOut[0] ;
    assign dataOut[121] = dataOut[0] ;
    assign dataOut[120] = dataOut[0] ;
    assign dataOut[119] = dataOut[0] ;
    assign dataOut[118] = dataOut[0] ;
    assign dataOut[117] = dataOut[0] ;
    assign dataOut[116] = dataOut[0] ;
    assign dataOut[115] = dataOut[0] ;
    assign dataOut[114] = dataOut[0] ;
    assign dataOut[113] = dataOut[0] ;
    assign dataOut[112] = dataOut[0] ;
    assign dataOut[111] = dataOut[0] ;
    assign dataOut[110] = dataOut[0] ;
    assign dataOut[109] = dataOut[0] ;
    assign dataOut[108] = dataOut[0] ;
    assign dataOut[107] = dataOut[0] ;
    assign dataOut[106] = dataOut[0] ;
    assign dataOut[105] = dataOut[0] ;
    assign dataOut[104] = dataOut[0] ;
    assign dataOut[103] = dataOut[0] ;
    assign dataOut[102] = dataOut[0] ;
    assign dataOut[101] = dataOut[0] ;
    assign dataOut[100] = dataOut[0] ;
    assign dataOut[99] = dataOut[0] ;
    assign dataOut[98] = dataOut[0] ;
    assign dataOut[97] = dataOut[0] ;
    assign dataOut[96] = dataOut[0] ;
    assign dataOut[95] = dataOut[0] ;
    assign dataOut[94] = dataOut[0] ;
    assign dataOut[93] = dataOut[0] ;
    assign dataOut[92] = dataOut[0] ;
    assign dataOut[91] = dataOut[0] ;
    assign dataOut[90] = dataOut[0] ;
    assign dataOut[89] = dataOut[0] ;
    assign dataOut[88] = dataOut[0] ;
    assign dataOut[87] = dataOut[0] ;
    assign dataOut[86] = dataOut[0] ;
    assign dataOut[85] = dataOut[0] ;
    assign dataOut[84] = dataOut[0] ;
    assign dataOut[83] = dataOut[0] ;
    assign dataOut[82] = dataOut[0] ;
    assign dataOut[81] = dataOut[0] ;
    assign dataOut[80] = dataOut[0] ;
    assign dataOut[79] = dataOut[0] ;
    assign dataOut[78] = dataOut[0] ;
    assign dataOut[77] = dataOut[0] ;
    assign dataOut[76] = dataOut[0] ;
    assign dataOut[75] = dataOut[0] ;
    assign dataOut[74] = dataOut[0] ;
    assign dataOut[73] = dataOut[0] ;
    assign dataOut[72] = dataOut[0] ;
    assign dataOut[71] = dataOut[0] ;
    assign dataOut[70] = dataOut[0] ;
    assign dataOut[69] = dataOut[0] ;
    assign dataOut[68] = dataOut[0] ;
    assign dataOut[67] = dataOut[0] ;
    assign dataOut[66] = dataOut[0] ;
    assign dataOut[65] = dataOut[0] ;
    assign dataOut[64] = dataOut[0] ;
    assign dataOut[63] = dataOut[0] ;
    assign dataOut[62] = dataOut[0] ;
    assign dataOut[61] = dataOut[0] ;
    assign dataOut[60] = dataOut[0] ;
    assign dataOut[59] = dataOut[0] ;
    assign dataOut[58] = dataOut[0] ;
    assign dataOut[57] = dataOut[0] ;
    assign dataOut[56] = dataOut[0] ;
    assign dataOut[55] = dataOut[0] ;
    assign dataOut[54] = dataOut[0] ;
    assign dataOut[53] = dataOut[0] ;
    assign dataOut[52] = dataOut[0] ;
    assign dataOut[51] = dataOut[0] ;
    assign dataOut[50] = dataOut[0] ;
    assign dataOut[49] = dataOut[0] ;
    assign dataOut[48] = dataOut[0] ;
    assign dataOut[47] = dataOut[0] ;
    assign dataOut[46] = dataOut[0] ;
    assign dataOut[45] = dataOut[0] ;
    assign dataOut[44] = dataOut[0] ;
    assign dataOut[43] = dataOut[0] ;
    assign dataOut[42] = dataOut[0] ;
    assign dataOut[41] = dataOut[0] ;
    assign dataOut[40] = dataOut[0] ;
    assign dataOut[39] = dataOut[0] ;
    assign dataOut[38] = dataOut[0] ;
    assign dataOut[37] = dataOut[0] ;
    assign dataOut[36] = dataOut[0] ;
    assign dataOut[35] = dataOut[0] ;
    assign dataOut[34] = dataOut[0] ;
    assign dataOut[33] = dataOut[0] ;
    assign dataOut[32] = dataOut[0] ;
    assign dataOut[31] = dataOut[0] ;
    assign dataOut[30] = dataOut[0] ;
    assign dataOut[29] = dataOut[0] ;
    assign dataOut[28] = dataOut[0] ;
    assign dataOut[27] = dataOut[0] ;
    assign dataOut[26] = dataOut[0] ;
    assign dataOut[25] = dataOut[0] ;
    assign dataOut[24] = dataOut[0] ;
    assign dataOut[23] = dataOut[0] ;
    assign dataOut[22] = dataOut[0] ;
    assign dataOut[21] = dataOut[0] ;
    assign dataOut[20] = dataOut[0] ;
    assign dataOut[19] = dataOut[0] ;
    assign dataOut[18] = dataOut[0] ;
    assign dataOut[17] = dataOut[0] ;
    assign dataOut[16] = dataOut[0] ;
    assign dataOut[15] = dataOut[0] ;
    assign dataOut[14] = dataOut[0] ;
    assign dataOut[13] = dataOut[0] ;
    assign dataOut[12] = dataOut[0] ;
    assign dataOut[11] = dataOut[0] ;
    assign dataOut[10] = dataOut[0] ;
    assign dataOut[9] = dataOut[0] ;
    assign dataOut[8] = dataOut[0] ;
    assign dataOut[7] = dataOut[0] ;
    assign dataOut[6] = dataOut[0] ;
    assign dataOut[5] = dataOut[0] ;
    assign dataOut[4] = dataOut[0] ;
    assign dataOut[3] = dataOut[0] ;
    assign dataOut[2] = dataOut[0] ;
    assign dataOut[1] = dataOut[0] ;
    fake_vcc ix117 (.Y (nx116)) ;
    ao21 ix61 (.Y (counterOut[1]), .A0 (dataIn[1]), .A1 (nx52), .B0 (nx46)) ;
    nor02_2x ix53 (.Y (nx52), .A0 (nx42), .A1 (nx46)) ;
    nor03_2x ix43 (.Y (nx42), .A0 (nx6871), .A1 (nx6873), .A2 (nx6876)) ;
    nand04 ix6872 (.Y (nx6871), .A0 (address[1]), .A1 (address[2]), .A2 (
           address[3]), .A3 (address[4])) ;
    nand03 ix6874 (.Y (nx6873), .A0 (address[5]), .A1 (address[6]), .A2 (nx12)
           ) ;
    nor02_2x ix13 (.Y (nx12), .A0 (address[12]), .A1 (address[11])) ;
    nand04 ix6877 (.Y (nx6876), .A0 (nx30), .A1 (nx34), .A2 (reset), .A3 (CLK)
           ) ;
    nor04 ix31 (.Y (nx30), .A0 (address[10]), .A1 (address[9]), .A2 (address[8])
          , .A3 (address[7])) ;
    nor02ii ix35 (.Y (nx34), .A0 (address[0]), .A1 (W)) ;
    inv01 ix6882 (.Y (nx6881), .A (R)) ;
    ao21 ix65 (.Y (counterOut[2]), .A0 (dataIn[2]), .A1 (nx52), .B0 (nx46)) ;
    ao21 ix57 (.Y (counterOut[0]), .A0 (dataIn[0]), .A1 (nx6888), .B0 (nx42)) ;
    and02 ix67 (.Y (counterOut[3]), .A0 (dataIn[3]), .A1 (nx52)) ;
    nor04 ix115 (.Y (nx114), .A0 (nx6895), .A1 (nx6897), .A2 (nx6899), .A3 (
          nx6903)) ;
    nand03 ix6896 (.Y (nx6895), .A0 (dataIn[7]), .A1 (dataIn[4]), .A2 (dataIn[5]
           )) ;
    nand02 ix6898 (.Y (nx6897), .A0 (dataIn[9]), .A1 (dataIn[12])) ;
    nand04 ix6900 (.Y (nx6899), .A0 (dataIn[0]), .A1 (dataIn[1]), .A2 (dataIn[2]
           ), .A3 (nx6901)) ;
    inv01 ix6902 (.Y (nx6901), .A (dataIn[15])) ;
    nand04 ix6904 (.Y (nx6903), .A0 (nx98), .A1 (nx104), .A2 (dataIn[3]), .A3 (
           nx6881)) ;
    nor04 ix99 (.Y (nx98), .A0 (dataIn[14]), .A1 (dataIn[13]), .A2 (dataIn[11])
          , .A3 (dataIn[10])) ;
    nor02_2x ix105 (.Y (nx104), .A0 (dataIn[8]), .A1 (dataIn[6])) ;
    and02 ix119 (.Y (nx118), .A0 (R), .A1 (CLK)) ;
    inv01 ix6889 (.Y (nx6888), .A (nx46)) ;
    nor02ii ix47 (.Y (nx46), .A0 (CLK), .A1 (R)) ;
    and03 ix129 (.Y (MFC), .A0 (reset), .A1 (R), .A2 (nx6914)) ;
    inv01 ix6913 (.Y (nx6914), .A (W)) ;
    latchr lat_dataOut_0__u1 (.QB (nx5), .D (nx116), .CLK (nx114), .R (nx118)) ;
    inv01 lat_dataOut_0__u2 (.Y (dataOut[0]), .A (nx5)) ;
    buf02 lat_dataOut_0__u3 (.Y (nx1), .A (nx5)) ;
endmodule


module triStateBuffer_16 ( D, EN, F ) ;

    input [15:0]D ;
    input EN ;
    output [15:0]F ;

    wire nx215, nx218, nx221, nx224, nx227, nx230, nx233, nx236, nx239, nx242, 
         nx245, nx248, nx251, nx254, nx257, nx260, nx267, nx269, nx271, nx273;



    tri01 tri_F_0 (.Y (F[0]), .A (nx215), .E (nx269)) ;
    inv01 ix216 (.Y (nx215), .A (D[0])) ;
    tri01 tri_F_1 (.Y (F[1]), .A (nx218), .E (nx269)) ;
    inv01 ix219 (.Y (nx218), .A (D[1])) ;
    tri01 tri_F_2 (.Y (F[2]), .A (nx221), .E (nx269)) ;
    inv01 ix222 (.Y (nx221), .A (D[2])) ;
    tri01 tri_F_3 (.Y (F[3]), .A (nx224), .E (nx269)) ;
    inv01 ix225 (.Y (nx224), .A (D[3])) ;
    tri01 tri_F_4 (.Y (F[4]), .A (nx227), .E (nx269)) ;
    inv01 ix228 (.Y (nx227), .A (D[4])) ;
    tri01 tri_F_5 (.Y (F[5]), .A (nx230), .E (nx269)) ;
    inv01 ix231 (.Y (nx230), .A (D[5])) ;
    tri01 tri_F_6 (.Y (F[6]), .A (nx233), .E (nx269)) ;
    inv01 ix234 (.Y (nx233), .A (D[6])) ;
    tri01 tri_F_7 (.Y (F[7]), .A (nx236), .E (nx271)) ;
    inv01 ix237 (.Y (nx236), .A (D[7])) ;
    tri01 tri_F_8 (.Y (F[8]), .A (nx239), .E (nx271)) ;
    inv01 ix240 (.Y (nx239), .A (D[8])) ;
    tri01 tri_F_9 (.Y (F[9]), .A (nx242), .E (nx271)) ;
    inv01 ix243 (.Y (nx242), .A (D[9])) ;
    tri01 tri_F_10 (.Y (F[10]), .A (nx245), .E (nx271)) ;
    inv01 ix246 (.Y (nx245), .A (D[10])) ;
    tri01 tri_F_11 (.Y (F[11]), .A (nx248), .E (nx271)) ;
    inv01 ix249 (.Y (nx248), .A (D[11])) ;
    tri01 tri_F_12 (.Y (F[12]), .A (nx251), .E (nx271)) ;
    inv01 ix252 (.Y (nx251), .A (D[12])) ;
    tri01 tri_F_13 (.Y (F[13]), .A (nx254), .E (nx271)) ;
    inv01 ix255 (.Y (nx254), .A (D[13])) ;
    tri01 tri_F_14 (.Y (F[14]), .A (nx257), .E (nx273)) ;
    inv01 ix258 (.Y (nx257), .A (D[14])) ;
    tri01 tri_F_15 (.Y (F[15]), .A (nx260), .E (nx273)) ;
    inv01 ix261 (.Y (nx260), .A (D[15])) ;
    inv01 ix266 (.Y (nx267), .A (EN)) ;
    inv01 ix268 (.Y (nx269), .A (nx267)) ;
    inv01 ix270 (.Y (nx271), .A (nx267)) ;
    inv01 ix272 (.Y (nx273), .A (nx267)) ;
endmodule


module triStateBuffer_448 ( D, EN, F ) ;

    input [447:0]D ;
    input EN ;
    output [447:0]F ;

    wire nx4535, nx4538, nx4541, nx4544, nx4547, nx4550, nx4553, nx4556, nx4559, 
         nx4562, nx4565, nx4568, nx4571, nx4574, nx4577, nx4580, nx4583, nx4586, 
         nx4589, nx4592, nx4595, nx4598, nx4601, nx4604, nx4607, nx4610, nx4613, 
         nx4616, nx4619, nx4622, nx4625, nx4628, nx4631, nx4634, nx4637, nx4640, 
         nx4643, nx4646, nx4649, nx4652, nx4655, nx4658, nx4661, nx4664, nx4667, 
         nx4670, nx4673, nx4676, nx4679, nx4682, nx4685, nx4688, nx4691, nx4694, 
         nx4697, nx4700, nx4703, nx4706, nx4709, nx4712, nx4715, nx4718, nx4721, 
         nx4724, nx4727, nx4730, nx4733, nx4736, nx4739, nx4742, nx4745, nx4748, 
         nx4751, nx4754, nx4757, nx4760, nx4763, nx4766, nx4769, nx4772, nx4775, 
         nx4778, nx4781, nx4784, nx4787, nx4790, nx4793, nx4796, nx4799, nx4802, 
         nx4805, nx4808, nx4811, nx4814, nx4817, nx4820, nx4823, nx4826, nx4829, 
         nx4832, nx4835, nx4838, nx4841, nx4844, nx4847, nx4850, nx4853, nx4856, 
         nx4859, nx4862, nx4865, nx4868, nx4871, nx4874, nx4877, nx4880, nx4883, 
         nx4886, nx4889, nx4892, nx4895, nx4898, nx4901, nx4904, nx4907, nx4910, 
         nx4913, nx4916, nx4919, nx4922, nx4925, nx4928, nx4931, nx4934, nx4937, 
         nx4940, nx4943, nx4946, nx4949, nx4952, nx4955, nx4958, nx4961, nx4964, 
         nx4967, nx4970, nx4973, nx4976, nx4979, nx4982, nx4985, nx4988, nx4991, 
         nx4994, nx4997, nx5000, nx5003, nx5006, nx5009, nx5012, nx5015, nx5018, 
         nx5021, nx5024, nx5027, nx5030, nx5033, nx5036, nx5039, nx5042, nx5045, 
         nx5048, nx5051, nx5054, nx5057, nx5060, nx5063, nx5066, nx5069, nx5072, 
         nx5075, nx5078, nx5081, nx5084, nx5087, nx5090, nx5093, nx5096, nx5099, 
         nx5102, nx5105, nx5108, nx5111, nx5114, nx5117, nx5120, nx5123, nx5126, 
         nx5129, nx5132, nx5135, nx5138, nx5141, nx5144, nx5147, nx5150, nx5153, 
         nx5156, nx5159, nx5162, nx5165, nx5168, nx5171, nx5174, nx5177, nx5180, 
         nx5183, nx5186, nx5189, nx5192, nx5195, nx5198, nx5201, nx5204, nx5207, 
         nx5210, nx5213, nx5216, nx5219, nx5222, nx5225, nx5228, nx5231, nx5234, 
         nx5237, nx5240, nx5243, nx5246, nx5249, nx5252, nx5255, nx5258, nx5261, 
         nx5264, nx5267, nx5270, nx5273, nx5276, nx5279, nx5282, nx5285, nx5288, 
         nx5291, nx5294, nx5297, nx5300, nx5303, nx5306, nx5309, nx5312, nx5315, 
         nx5318, nx5321, nx5324, nx5327, nx5330, nx5333, nx5336, nx5339, nx5342, 
         nx5345, nx5348, nx5351, nx5354, nx5357, nx5360, nx5363, nx5366, nx5369, 
         nx5372, nx5375, nx5378, nx5381, nx5384, nx5387, nx5390, nx5393, nx5396, 
         nx5399, nx5402, nx5405, nx5408, nx5411, nx5414, nx5417, nx5420, nx5423, 
         nx5426, nx5429, nx5432, nx5435, nx5438, nx5441, nx5444, nx5447, nx5450, 
         nx5453, nx5456, nx5459, nx5462, nx5465, nx5468, nx5471, nx5474, nx5477, 
         nx5480, nx5483, nx5486, nx5489, nx5492, nx5495, nx5498, nx5501, nx5504, 
         nx5507, nx5510, nx5513, nx5516, nx5519, nx5522, nx5525, nx5528, nx5531, 
         nx5534, nx5537, nx5540, nx5543, nx5546, nx5549, nx5552, nx5555, nx5558, 
         nx5561, nx5564, nx5567, nx5570, nx5573, nx5576, nx5579, nx5582, nx5585, 
         nx5588, nx5591, nx5594, nx5597, nx5600, nx5603, nx5606, nx5609, nx5612, 
         nx5615, nx5618, nx5621, nx5624, nx5627, nx5630, nx5633, nx5636, nx5639, 
         nx5642, nx5645, nx5648, nx5651, nx5654, nx5657, nx5660, nx5663, nx5666, 
         nx5669, nx5672, nx5675, nx5678, nx5681, nx5684, nx5687, nx5690, nx5693, 
         nx5696, nx5699, nx5702, nx5705, nx5708, nx5711, nx5714, nx5717, nx5720, 
         nx5723, nx5726, nx5729, nx5732, nx5735, nx5738, nx5741, nx5744, nx5747, 
         nx5750, nx5753, nx5756, nx5759, nx5762, nx5765, nx5768, nx5771, nx5774, 
         nx5777, nx5780, nx5783, nx5786, nx5789, nx5792, nx5795, nx5798, nx5801, 
         nx5804, nx5807, nx5810, nx5813, nx5816, nx5819, nx5822, nx5825, nx5828, 
         nx5831, nx5834, nx5837, nx5840, nx5843, nx5846, nx5849, nx5852, nx5855, 
         nx5858, nx5861, nx5864, nx5867, nx5870, nx5873, nx5876, nx5883, nx5885, 
         nx5887, nx5889, nx5891, nx5893, nx5895, nx5897, nx5899, nx5901, nx5903, 
         nx5905, nx5907, nx5909, nx5911, nx5913, nx5915, nx5917, nx5919, nx5921, 
         nx5923, nx5925, nx5927, nx5929, nx5931, nx5933, nx5935, nx5937, nx5939, 
         nx5941, nx5943, nx5945, nx5947, nx5949, nx5951, nx5953, nx5955, nx5957, 
         nx5959, nx5961, nx5963, nx5965, nx5967, nx5969, nx5971, nx5973, nx5975, 
         nx5977, nx5979, nx5981, nx5983, nx5985, nx5987, nx5989, nx5991, nx5993, 
         nx5995, nx5997, nx5999, nx6001, nx6003, nx6005, nx6007, nx6009, nx6011, 
         nx6013, nx6015, nx6017, nx6019, nx6021, nx6023, nx6025, nx6027, nx6029, 
         nx6035, nx6037;



    tri01 tri_F_0 (.Y (F[0]), .A (nx4535), .E (nx5885)) ;
    inv01 ix4536 (.Y (nx4535), .A (D[0])) ;
    tri01 tri_F_1 (.Y (F[1]), .A (nx4538), .E (nx5885)) ;
    inv01 ix4539 (.Y (nx4538), .A (D[1])) ;
    tri01 tri_F_2 (.Y (F[2]), .A (nx4541), .E (nx5885)) ;
    inv01 ix4542 (.Y (nx4541), .A (D[2])) ;
    tri01 tri_F_3 (.Y (F[3]), .A (nx4544), .E (nx5885)) ;
    inv01 ix4545 (.Y (nx4544), .A (D[3])) ;
    tri01 tri_F_4 (.Y (F[4]), .A (nx4547), .E (nx5885)) ;
    inv01 ix4548 (.Y (nx4547), .A (D[4])) ;
    tri01 tri_F_5 (.Y (F[5]), .A (nx4550), .E (nx5885)) ;
    inv01 ix4551 (.Y (nx4550), .A (D[5])) ;
    tri01 tri_F_6 (.Y (F[6]), .A (nx4553), .E (nx5885)) ;
    inv01 ix4554 (.Y (nx4553), .A (D[6])) ;
    tri01 tri_F_7 (.Y (F[7]), .A (nx4556), .E (nx5887)) ;
    inv01 ix4557 (.Y (nx4556), .A (D[7])) ;
    tri01 tri_F_8 (.Y (F[8]), .A (nx4559), .E (nx5887)) ;
    inv01 ix4560 (.Y (nx4559), .A (D[8])) ;
    tri01 tri_F_9 (.Y (F[9]), .A (nx4562), .E (nx5887)) ;
    inv01 ix4563 (.Y (nx4562), .A (D[9])) ;
    tri01 tri_F_10 (.Y (F[10]), .A (nx4565), .E (nx5887)) ;
    inv01 ix4566 (.Y (nx4565), .A (D[10])) ;
    tri01 tri_F_11 (.Y (F[11]), .A (nx4568), .E (nx5887)) ;
    inv01 ix4569 (.Y (nx4568), .A (D[11])) ;
    tri01 tri_F_12 (.Y (F[12]), .A (nx4571), .E (nx5887)) ;
    inv01 ix4572 (.Y (nx4571), .A (D[12])) ;
    tri01 tri_F_13 (.Y (F[13]), .A (nx4574), .E (nx5887)) ;
    inv01 ix4575 (.Y (nx4574), .A (D[13])) ;
    tri01 tri_F_14 (.Y (F[14]), .A (nx4577), .E (nx5889)) ;
    inv01 ix4578 (.Y (nx4577), .A (D[14])) ;
    tri01 tri_F_15 (.Y (F[15]), .A (nx4580), .E (nx5889)) ;
    inv01 ix4581 (.Y (nx4580), .A (D[15])) ;
    tri01 tri_F_16 (.Y (F[16]), .A (nx4583), .E (nx5889)) ;
    inv01 ix4584 (.Y (nx4583), .A (D[16])) ;
    tri01 tri_F_17 (.Y (F[17]), .A (nx4586), .E (nx5889)) ;
    inv01 ix4587 (.Y (nx4586), .A (D[17])) ;
    tri01 tri_F_18 (.Y (F[18]), .A (nx4589), .E (nx5889)) ;
    inv01 ix4590 (.Y (nx4589), .A (D[18])) ;
    tri01 tri_F_19 (.Y (F[19]), .A (nx4592), .E (nx5889)) ;
    inv01 ix4593 (.Y (nx4592), .A (D[19])) ;
    tri01 tri_F_20 (.Y (F[20]), .A (nx4595), .E (nx5889)) ;
    inv01 ix4596 (.Y (nx4595), .A (D[20])) ;
    tri01 tri_F_21 (.Y (F[21]), .A (nx4598), .E (nx5891)) ;
    inv01 ix4599 (.Y (nx4598), .A (D[21])) ;
    tri01 tri_F_22 (.Y (F[22]), .A (nx4601), .E (nx5891)) ;
    inv01 ix4602 (.Y (nx4601), .A (D[22])) ;
    tri01 tri_F_23 (.Y (F[23]), .A (nx4604), .E (nx5891)) ;
    inv01 ix4605 (.Y (nx4604), .A (D[23])) ;
    tri01 tri_F_24 (.Y (F[24]), .A (nx4607), .E (nx5891)) ;
    inv01 ix4608 (.Y (nx4607), .A (D[24])) ;
    tri01 tri_F_25 (.Y (F[25]), .A (nx4610), .E (nx5891)) ;
    inv01 ix4611 (.Y (nx4610), .A (D[25])) ;
    tri01 tri_F_26 (.Y (F[26]), .A (nx4613), .E (nx5891)) ;
    inv01 ix4614 (.Y (nx4613), .A (D[26])) ;
    tri01 tri_F_27 (.Y (F[27]), .A (nx4616), .E (nx5891)) ;
    inv01 ix4617 (.Y (nx4616), .A (D[27])) ;
    tri01 tri_F_28 (.Y (F[28]), .A (nx4619), .E (nx5893)) ;
    inv01 ix4620 (.Y (nx4619), .A (D[28])) ;
    tri01 tri_F_29 (.Y (F[29]), .A (nx4622), .E (nx5893)) ;
    inv01 ix4623 (.Y (nx4622), .A (D[29])) ;
    tri01 tri_F_30 (.Y (F[30]), .A (nx4625), .E (nx5893)) ;
    inv01 ix4626 (.Y (nx4625), .A (D[30])) ;
    tri01 tri_F_31 (.Y (F[31]), .A (nx4628), .E (nx5893)) ;
    inv01 ix4629 (.Y (nx4628), .A (D[31])) ;
    tri01 tri_F_32 (.Y (F[32]), .A (nx4631), .E (nx5893)) ;
    inv01 ix4632 (.Y (nx4631), .A (D[32])) ;
    tri01 tri_F_33 (.Y (F[33]), .A (nx4634), .E (nx5893)) ;
    inv01 ix4635 (.Y (nx4634), .A (D[33])) ;
    tri01 tri_F_34 (.Y (F[34]), .A (nx4637), .E (nx5893)) ;
    inv01 ix4638 (.Y (nx4637), .A (D[34])) ;
    tri01 tri_F_35 (.Y (F[35]), .A (nx4640), .E (nx5895)) ;
    inv01 ix4641 (.Y (nx4640), .A (D[35])) ;
    tri01 tri_F_36 (.Y (F[36]), .A (nx4643), .E (nx5895)) ;
    inv01 ix4644 (.Y (nx4643), .A (D[36])) ;
    tri01 tri_F_37 (.Y (F[37]), .A (nx4646), .E (nx5895)) ;
    inv01 ix4647 (.Y (nx4646), .A (D[37])) ;
    tri01 tri_F_38 (.Y (F[38]), .A (nx4649), .E (nx5895)) ;
    inv01 ix4650 (.Y (nx4649), .A (D[38])) ;
    tri01 tri_F_39 (.Y (F[39]), .A (nx4652), .E (nx5895)) ;
    inv01 ix4653 (.Y (nx4652), .A (D[39])) ;
    tri01 tri_F_40 (.Y (F[40]), .A (nx4655), .E (nx5895)) ;
    inv01 ix4656 (.Y (nx4655), .A (D[40])) ;
    tri01 tri_F_41 (.Y (F[41]), .A (nx4658), .E (nx5895)) ;
    inv01 ix4659 (.Y (nx4658), .A (D[41])) ;
    tri01 tri_F_42 (.Y (F[42]), .A (nx4661), .E (nx5897)) ;
    inv01 ix4662 (.Y (nx4661), .A (D[42])) ;
    tri01 tri_F_43 (.Y (F[43]), .A (nx4664), .E (nx5897)) ;
    inv01 ix4665 (.Y (nx4664), .A (D[43])) ;
    tri01 tri_F_44 (.Y (F[44]), .A (nx4667), .E (nx5897)) ;
    inv01 ix4668 (.Y (nx4667), .A (D[44])) ;
    tri01 tri_F_45 (.Y (F[45]), .A (nx4670), .E (nx5897)) ;
    inv01 ix4671 (.Y (nx4670), .A (D[45])) ;
    tri01 tri_F_46 (.Y (F[46]), .A (nx4673), .E (nx5897)) ;
    inv01 ix4674 (.Y (nx4673), .A (D[46])) ;
    tri01 tri_F_47 (.Y (F[47]), .A (nx4676), .E (nx5897)) ;
    inv01 ix4677 (.Y (nx4676), .A (D[47])) ;
    tri01 tri_F_48 (.Y (F[48]), .A (nx4679), .E (nx5897)) ;
    inv01 ix4680 (.Y (nx4679), .A (D[48])) ;
    tri01 tri_F_49 (.Y (F[49]), .A (nx4682), .E (nx5899)) ;
    inv01 ix4683 (.Y (nx4682), .A (D[49])) ;
    tri01 tri_F_50 (.Y (F[50]), .A (nx4685), .E (nx5899)) ;
    inv01 ix4686 (.Y (nx4685), .A (D[50])) ;
    tri01 tri_F_51 (.Y (F[51]), .A (nx4688), .E (nx5899)) ;
    inv01 ix4689 (.Y (nx4688), .A (D[51])) ;
    tri01 tri_F_52 (.Y (F[52]), .A (nx4691), .E (nx5899)) ;
    inv01 ix4692 (.Y (nx4691), .A (D[52])) ;
    tri01 tri_F_53 (.Y (F[53]), .A (nx4694), .E (nx5899)) ;
    inv01 ix4695 (.Y (nx4694), .A (D[53])) ;
    tri01 tri_F_54 (.Y (F[54]), .A (nx4697), .E (nx5899)) ;
    inv01 ix4698 (.Y (nx4697), .A (D[54])) ;
    tri01 tri_F_55 (.Y (F[55]), .A (nx4700), .E (nx5899)) ;
    inv01 ix4701 (.Y (nx4700), .A (D[55])) ;
    tri01 tri_F_56 (.Y (F[56]), .A (nx4703), .E (nx5901)) ;
    inv01 ix4704 (.Y (nx4703), .A (D[56])) ;
    tri01 tri_F_57 (.Y (F[57]), .A (nx4706), .E (nx5901)) ;
    inv01 ix4707 (.Y (nx4706), .A (D[57])) ;
    tri01 tri_F_58 (.Y (F[58]), .A (nx4709), .E (nx5901)) ;
    inv01 ix4710 (.Y (nx4709), .A (D[58])) ;
    tri01 tri_F_59 (.Y (F[59]), .A (nx4712), .E (nx5901)) ;
    inv01 ix4713 (.Y (nx4712), .A (D[59])) ;
    tri01 tri_F_60 (.Y (F[60]), .A (nx4715), .E (nx5901)) ;
    inv01 ix4716 (.Y (nx4715), .A (D[60])) ;
    tri01 tri_F_61 (.Y (F[61]), .A (nx4718), .E (nx5901)) ;
    inv01 ix4719 (.Y (nx4718), .A (D[61])) ;
    tri01 tri_F_62 (.Y (F[62]), .A (nx4721), .E (nx5901)) ;
    inv01 ix4722 (.Y (nx4721), .A (D[62])) ;
    tri01 tri_F_63 (.Y (F[63]), .A (nx4724), .E (nx5903)) ;
    inv01 ix4725 (.Y (nx4724), .A (D[63])) ;
    tri01 tri_F_64 (.Y (F[64]), .A (nx4727), .E (nx5903)) ;
    inv01 ix4728 (.Y (nx4727), .A (D[64])) ;
    tri01 tri_F_65 (.Y (F[65]), .A (nx4730), .E (nx5903)) ;
    inv01 ix4731 (.Y (nx4730), .A (D[65])) ;
    tri01 tri_F_66 (.Y (F[66]), .A (nx4733), .E (nx5903)) ;
    inv01 ix4734 (.Y (nx4733), .A (D[66])) ;
    tri01 tri_F_67 (.Y (F[67]), .A (nx4736), .E (nx5903)) ;
    inv01 ix4737 (.Y (nx4736), .A (D[67])) ;
    tri01 tri_F_68 (.Y (F[68]), .A (nx4739), .E (nx5903)) ;
    inv01 ix4740 (.Y (nx4739), .A (D[68])) ;
    tri01 tri_F_69 (.Y (F[69]), .A (nx4742), .E (nx5903)) ;
    inv01 ix4743 (.Y (nx4742), .A (D[69])) ;
    tri01 tri_F_70 (.Y (F[70]), .A (nx4745), .E (nx5905)) ;
    inv01 ix4746 (.Y (nx4745), .A (D[70])) ;
    tri01 tri_F_71 (.Y (F[71]), .A (nx4748), .E (nx5905)) ;
    inv01 ix4749 (.Y (nx4748), .A (D[71])) ;
    tri01 tri_F_72 (.Y (F[72]), .A (nx4751), .E (nx5905)) ;
    inv01 ix4752 (.Y (nx4751), .A (D[72])) ;
    tri01 tri_F_73 (.Y (F[73]), .A (nx4754), .E (nx5905)) ;
    inv01 ix4755 (.Y (nx4754), .A (D[73])) ;
    tri01 tri_F_74 (.Y (F[74]), .A (nx4757), .E (nx5905)) ;
    inv01 ix4758 (.Y (nx4757), .A (D[74])) ;
    tri01 tri_F_75 (.Y (F[75]), .A (nx4760), .E (nx5905)) ;
    inv01 ix4761 (.Y (nx4760), .A (D[75])) ;
    tri01 tri_F_76 (.Y (F[76]), .A (nx4763), .E (nx5905)) ;
    inv01 ix4764 (.Y (nx4763), .A (D[76])) ;
    tri01 tri_F_77 (.Y (F[77]), .A (nx4766), .E (nx5907)) ;
    inv01 ix4767 (.Y (nx4766), .A (D[77])) ;
    tri01 tri_F_78 (.Y (F[78]), .A (nx4769), .E (nx5907)) ;
    inv01 ix4770 (.Y (nx4769), .A (D[78])) ;
    tri01 tri_F_79 (.Y (F[79]), .A (nx4772), .E (nx5907)) ;
    inv01 ix4773 (.Y (nx4772), .A (D[79])) ;
    tri01 tri_F_80 (.Y (F[80]), .A (nx4775), .E (nx5907)) ;
    inv01 ix4776 (.Y (nx4775), .A (D[80])) ;
    tri01 tri_F_81 (.Y (F[81]), .A (nx4778), .E (nx5907)) ;
    inv01 ix4779 (.Y (nx4778), .A (D[81])) ;
    tri01 tri_F_82 (.Y (F[82]), .A (nx4781), .E (nx5907)) ;
    inv01 ix4782 (.Y (nx4781), .A (D[82])) ;
    tri01 tri_F_83 (.Y (F[83]), .A (nx4784), .E (nx5907)) ;
    inv01 ix4785 (.Y (nx4784), .A (D[83])) ;
    tri01 tri_F_84 (.Y (F[84]), .A (nx4787), .E (nx5909)) ;
    inv01 ix4788 (.Y (nx4787), .A (D[84])) ;
    tri01 tri_F_85 (.Y (F[85]), .A (nx4790), .E (nx5909)) ;
    inv01 ix4791 (.Y (nx4790), .A (D[85])) ;
    tri01 tri_F_86 (.Y (F[86]), .A (nx4793), .E (nx5909)) ;
    inv01 ix4794 (.Y (nx4793), .A (D[86])) ;
    tri01 tri_F_87 (.Y (F[87]), .A (nx4796), .E (nx5909)) ;
    inv01 ix4797 (.Y (nx4796), .A (D[87])) ;
    tri01 tri_F_88 (.Y (F[88]), .A (nx4799), .E (nx5909)) ;
    inv01 ix4800 (.Y (nx4799), .A (D[88])) ;
    tri01 tri_F_89 (.Y (F[89]), .A (nx4802), .E (nx5909)) ;
    inv01 ix4803 (.Y (nx4802), .A (D[89])) ;
    tri01 tri_F_90 (.Y (F[90]), .A (nx4805), .E (nx5909)) ;
    inv01 ix4806 (.Y (nx4805), .A (D[90])) ;
    tri01 tri_F_91 (.Y (F[91]), .A (nx4808), .E (nx5911)) ;
    inv01 ix4809 (.Y (nx4808), .A (D[91])) ;
    tri01 tri_F_92 (.Y (F[92]), .A (nx4811), .E (nx5911)) ;
    inv01 ix4812 (.Y (nx4811), .A (D[92])) ;
    tri01 tri_F_93 (.Y (F[93]), .A (nx4814), .E (nx5911)) ;
    inv01 ix4815 (.Y (nx4814), .A (D[93])) ;
    tri01 tri_F_94 (.Y (F[94]), .A (nx4817), .E (nx5911)) ;
    inv01 ix4818 (.Y (nx4817), .A (D[94])) ;
    tri01 tri_F_95 (.Y (F[95]), .A (nx4820), .E (nx5911)) ;
    inv01 ix4821 (.Y (nx4820), .A (D[95])) ;
    tri01 tri_F_96 (.Y (F[96]), .A (nx4823), .E (nx5911)) ;
    inv01 ix4824 (.Y (nx4823), .A (D[96])) ;
    tri01 tri_F_97 (.Y (F[97]), .A (nx4826), .E (nx5911)) ;
    inv01 ix4827 (.Y (nx4826), .A (D[97])) ;
    tri01 tri_F_98 (.Y (F[98]), .A (nx4829), .E (nx5913)) ;
    inv01 ix4830 (.Y (nx4829), .A (D[98])) ;
    tri01 tri_F_99 (.Y (F[99]), .A (nx4832), .E (nx5913)) ;
    inv01 ix4833 (.Y (nx4832), .A (D[99])) ;
    tri01 tri_F_100 (.Y (F[100]), .A (nx4835), .E (nx5913)) ;
    inv01 ix4836 (.Y (nx4835), .A (D[100])) ;
    tri01 tri_F_101 (.Y (F[101]), .A (nx4838), .E (nx5913)) ;
    inv01 ix4839 (.Y (nx4838), .A (D[101])) ;
    tri01 tri_F_102 (.Y (F[102]), .A (nx4841), .E (nx5913)) ;
    inv01 ix4842 (.Y (nx4841), .A (D[102])) ;
    tri01 tri_F_103 (.Y (F[103]), .A (nx4844), .E (nx5913)) ;
    inv01 ix4845 (.Y (nx4844), .A (D[103])) ;
    tri01 tri_F_104 (.Y (F[104]), .A (nx4847), .E (nx5913)) ;
    inv01 ix4848 (.Y (nx4847), .A (D[104])) ;
    tri01 tri_F_105 (.Y (F[105]), .A (nx4850), .E (nx5915)) ;
    inv01 ix4851 (.Y (nx4850), .A (D[105])) ;
    tri01 tri_F_106 (.Y (F[106]), .A (nx4853), .E (nx5915)) ;
    inv01 ix4854 (.Y (nx4853), .A (D[106])) ;
    tri01 tri_F_107 (.Y (F[107]), .A (nx4856), .E (nx5915)) ;
    inv01 ix4857 (.Y (nx4856), .A (D[107])) ;
    tri01 tri_F_108 (.Y (F[108]), .A (nx4859), .E (nx5915)) ;
    inv01 ix4860 (.Y (nx4859), .A (D[108])) ;
    tri01 tri_F_109 (.Y (F[109]), .A (nx4862), .E (nx5915)) ;
    inv01 ix4863 (.Y (nx4862), .A (D[109])) ;
    tri01 tri_F_110 (.Y (F[110]), .A (nx4865), .E (nx5915)) ;
    inv01 ix4866 (.Y (nx4865), .A (D[110])) ;
    tri01 tri_F_111 (.Y (F[111]), .A (nx4868), .E (nx5915)) ;
    inv01 ix4869 (.Y (nx4868), .A (D[111])) ;
    tri01 tri_F_112 (.Y (F[112]), .A (nx4871), .E (nx5917)) ;
    inv01 ix4872 (.Y (nx4871), .A (D[112])) ;
    tri01 tri_F_113 (.Y (F[113]), .A (nx4874), .E (nx5917)) ;
    inv01 ix4875 (.Y (nx4874), .A (D[113])) ;
    tri01 tri_F_114 (.Y (F[114]), .A (nx4877), .E (nx5917)) ;
    inv01 ix4878 (.Y (nx4877), .A (D[114])) ;
    tri01 tri_F_115 (.Y (F[115]), .A (nx4880), .E (nx5917)) ;
    inv01 ix4881 (.Y (nx4880), .A (D[115])) ;
    tri01 tri_F_116 (.Y (F[116]), .A (nx4883), .E (nx5917)) ;
    inv01 ix4884 (.Y (nx4883), .A (D[116])) ;
    tri01 tri_F_117 (.Y (F[117]), .A (nx4886), .E (nx5917)) ;
    inv01 ix4887 (.Y (nx4886), .A (D[117])) ;
    tri01 tri_F_118 (.Y (F[118]), .A (nx4889), .E (nx5917)) ;
    inv01 ix4890 (.Y (nx4889), .A (D[118])) ;
    tri01 tri_F_119 (.Y (F[119]), .A (nx4892), .E (nx5919)) ;
    inv01 ix4893 (.Y (nx4892), .A (D[119])) ;
    tri01 tri_F_120 (.Y (F[120]), .A (nx4895), .E (nx5919)) ;
    inv01 ix4896 (.Y (nx4895), .A (D[120])) ;
    tri01 tri_F_121 (.Y (F[121]), .A (nx4898), .E (nx5919)) ;
    inv01 ix4899 (.Y (nx4898), .A (D[121])) ;
    tri01 tri_F_122 (.Y (F[122]), .A (nx4901), .E (nx5919)) ;
    inv01 ix4902 (.Y (nx4901), .A (D[122])) ;
    tri01 tri_F_123 (.Y (F[123]), .A (nx4904), .E (nx5919)) ;
    inv01 ix4905 (.Y (nx4904), .A (D[123])) ;
    tri01 tri_F_124 (.Y (F[124]), .A (nx4907), .E (nx5919)) ;
    inv01 ix4908 (.Y (nx4907), .A (D[124])) ;
    tri01 tri_F_125 (.Y (F[125]), .A (nx4910), .E (nx5919)) ;
    inv01 ix4911 (.Y (nx4910), .A (D[125])) ;
    tri01 tri_F_126 (.Y (F[126]), .A (nx4913), .E (nx5921)) ;
    inv01 ix4914 (.Y (nx4913), .A (D[126])) ;
    tri01 tri_F_127 (.Y (F[127]), .A (nx4916), .E (nx5921)) ;
    inv01 ix4917 (.Y (nx4916), .A (D[127])) ;
    tri01 tri_F_128 (.Y (F[128]), .A (nx4919), .E (nx5921)) ;
    inv01 ix4920 (.Y (nx4919), .A (D[128])) ;
    tri01 tri_F_129 (.Y (F[129]), .A (nx4922), .E (nx5921)) ;
    inv01 ix4923 (.Y (nx4922), .A (D[129])) ;
    tri01 tri_F_130 (.Y (F[130]), .A (nx4925), .E (nx5921)) ;
    inv01 ix4926 (.Y (nx4925), .A (D[130])) ;
    tri01 tri_F_131 (.Y (F[131]), .A (nx4928), .E (nx5921)) ;
    inv01 ix4929 (.Y (nx4928), .A (D[131])) ;
    tri01 tri_F_132 (.Y (F[132]), .A (nx4931), .E (nx5921)) ;
    inv01 ix4932 (.Y (nx4931), .A (D[132])) ;
    tri01 tri_F_133 (.Y (F[133]), .A (nx4934), .E (nx5923)) ;
    inv01 ix4935 (.Y (nx4934), .A (D[133])) ;
    tri01 tri_F_134 (.Y (F[134]), .A (nx4937), .E (nx5923)) ;
    inv01 ix4938 (.Y (nx4937), .A (D[134])) ;
    tri01 tri_F_135 (.Y (F[135]), .A (nx4940), .E (nx5923)) ;
    inv01 ix4941 (.Y (nx4940), .A (D[135])) ;
    tri01 tri_F_136 (.Y (F[136]), .A (nx4943), .E (nx5923)) ;
    inv01 ix4944 (.Y (nx4943), .A (D[136])) ;
    tri01 tri_F_137 (.Y (F[137]), .A (nx4946), .E (nx5923)) ;
    inv01 ix4947 (.Y (nx4946), .A (D[137])) ;
    tri01 tri_F_138 (.Y (F[138]), .A (nx4949), .E (nx5923)) ;
    inv01 ix4950 (.Y (nx4949), .A (D[138])) ;
    tri01 tri_F_139 (.Y (F[139]), .A (nx4952), .E (nx5923)) ;
    inv01 ix4953 (.Y (nx4952), .A (D[139])) ;
    tri01 tri_F_140 (.Y (F[140]), .A (nx4955), .E (nx5925)) ;
    inv01 ix4956 (.Y (nx4955), .A (D[140])) ;
    tri01 tri_F_141 (.Y (F[141]), .A (nx4958), .E (nx5925)) ;
    inv01 ix4959 (.Y (nx4958), .A (D[141])) ;
    tri01 tri_F_142 (.Y (F[142]), .A (nx4961), .E (nx5925)) ;
    inv01 ix4962 (.Y (nx4961), .A (D[142])) ;
    tri01 tri_F_143 (.Y (F[143]), .A (nx4964), .E (nx5925)) ;
    inv01 ix4965 (.Y (nx4964), .A (D[143])) ;
    tri01 tri_F_144 (.Y (F[144]), .A (nx4967), .E (nx5925)) ;
    inv01 ix4968 (.Y (nx4967), .A (D[144])) ;
    tri01 tri_F_145 (.Y (F[145]), .A (nx4970), .E (nx5925)) ;
    inv01 ix4971 (.Y (nx4970), .A (D[145])) ;
    tri01 tri_F_146 (.Y (F[146]), .A (nx4973), .E (nx5925)) ;
    inv01 ix4974 (.Y (nx4973), .A (D[146])) ;
    tri01 tri_F_147 (.Y (F[147]), .A (nx4976), .E (nx5927)) ;
    inv01 ix4977 (.Y (nx4976), .A (D[147])) ;
    tri01 tri_F_148 (.Y (F[148]), .A (nx4979), .E (nx5927)) ;
    inv01 ix4980 (.Y (nx4979), .A (D[148])) ;
    tri01 tri_F_149 (.Y (F[149]), .A (nx4982), .E (nx5927)) ;
    inv01 ix4983 (.Y (nx4982), .A (D[149])) ;
    tri01 tri_F_150 (.Y (F[150]), .A (nx4985), .E (nx5927)) ;
    inv01 ix4986 (.Y (nx4985), .A (D[150])) ;
    tri01 tri_F_151 (.Y (F[151]), .A (nx4988), .E (nx5927)) ;
    inv01 ix4989 (.Y (nx4988), .A (D[151])) ;
    tri01 tri_F_152 (.Y (F[152]), .A (nx4991), .E (nx5927)) ;
    inv01 ix4992 (.Y (nx4991), .A (D[152])) ;
    tri01 tri_F_153 (.Y (F[153]), .A (nx4994), .E (nx5927)) ;
    inv01 ix4995 (.Y (nx4994), .A (D[153])) ;
    tri01 tri_F_154 (.Y (F[154]), .A (nx4997), .E (nx5929)) ;
    inv01 ix4998 (.Y (nx4997), .A (D[154])) ;
    tri01 tri_F_155 (.Y (F[155]), .A (nx5000), .E (nx5929)) ;
    inv01 ix5001 (.Y (nx5000), .A (D[155])) ;
    tri01 tri_F_156 (.Y (F[156]), .A (nx5003), .E (nx5929)) ;
    inv01 ix5004 (.Y (nx5003), .A (D[156])) ;
    tri01 tri_F_157 (.Y (F[157]), .A (nx5006), .E (nx5929)) ;
    inv01 ix5007 (.Y (nx5006), .A (D[157])) ;
    tri01 tri_F_158 (.Y (F[158]), .A (nx5009), .E (nx5929)) ;
    inv01 ix5010 (.Y (nx5009), .A (D[158])) ;
    tri01 tri_F_159 (.Y (F[159]), .A (nx5012), .E (nx5929)) ;
    inv01 ix5013 (.Y (nx5012), .A (D[159])) ;
    tri01 tri_F_160 (.Y (F[160]), .A (nx5015), .E (nx5929)) ;
    inv01 ix5016 (.Y (nx5015), .A (D[160])) ;
    tri01 tri_F_161 (.Y (F[161]), .A (nx5018), .E (nx5931)) ;
    inv01 ix5019 (.Y (nx5018), .A (D[161])) ;
    tri01 tri_F_162 (.Y (F[162]), .A (nx5021), .E (nx5931)) ;
    inv01 ix5022 (.Y (nx5021), .A (D[162])) ;
    tri01 tri_F_163 (.Y (F[163]), .A (nx5024), .E (nx5931)) ;
    inv01 ix5025 (.Y (nx5024), .A (D[163])) ;
    tri01 tri_F_164 (.Y (F[164]), .A (nx5027), .E (nx5931)) ;
    inv01 ix5028 (.Y (nx5027), .A (D[164])) ;
    tri01 tri_F_165 (.Y (F[165]), .A (nx5030), .E (nx5931)) ;
    inv01 ix5031 (.Y (nx5030), .A (D[165])) ;
    tri01 tri_F_166 (.Y (F[166]), .A (nx5033), .E (nx5931)) ;
    inv01 ix5034 (.Y (nx5033), .A (D[166])) ;
    tri01 tri_F_167 (.Y (F[167]), .A (nx5036), .E (nx5931)) ;
    inv01 ix5037 (.Y (nx5036), .A (D[167])) ;
    tri01 tri_F_168 (.Y (F[168]), .A (nx5039), .E (nx5933)) ;
    inv01 ix5040 (.Y (nx5039), .A (D[168])) ;
    tri01 tri_F_169 (.Y (F[169]), .A (nx5042), .E (nx5933)) ;
    inv01 ix5043 (.Y (nx5042), .A (D[169])) ;
    tri01 tri_F_170 (.Y (F[170]), .A (nx5045), .E (nx5933)) ;
    inv01 ix5046 (.Y (nx5045), .A (D[170])) ;
    tri01 tri_F_171 (.Y (F[171]), .A (nx5048), .E (nx5933)) ;
    inv01 ix5049 (.Y (nx5048), .A (D[171])) ;
    tri01 tri_F_172 (.Y (F[172]), .A (nx5051), .E (nx5933)) ;
    inv01 ix5052 (.Y (nx5051), .A (D[172])) ;
    tri01 tri_F_173 (.Y (F[173]), .A (nx5054), .E (nx5933)) ;
    inv01 ix5055 (.Y (nx5054), .A (D[173])) ;
    tri01 tri_F_174 (.Y (F[174]), .A (nx5057), .E (nx5933)) ;
    inv01 ix5058 (.Y (nx5057), .A (D[174])) ;
    tri01 tri_F_175 (.Y (F[175]), .A (nx5060), .E (nx5935)) ;
    inv01 ix5061 (.Y (nx5060), .A (D[175])) ;
    tri01 tri_F_176 (.Y (F[176]), .A (nx5063), .E (nx5935)) ;
    inv01 ix5064 (.Y (nx5063), .A (D[176])) ;
    tri01 tri_F_177 (.Y (F[177]), .A (nx5066), .E (nx5935)) ;
    inv01 ix5067 (.Y (nx5066), .A (D[177])) ;
    tri01 tri_F_178 (.Y (F[178]), .A (nx5069), .E (nx5935)) ;
    inv01 ix5070 (.Y (nx5069), .A (D[178])) ;
    tri01 tri_F_179 (.Y (F[179]), .A (nx5072), .E (nx5935)) ;
    inv01 ix5073 (.Y (nx5072), .A (D[179])) ;
    tri01 tri_F_180 (.Y (F[180]), .A (nx5075), .E (nx5935)) ;
    inv01 ix5076 (.Y (nx5075), .A (D[180])) ;
    tri01 tri_F_181 (.Y (F[181]), .A (nx5078), .E (nx5935)) ;
    inv01 ix5079 (.Y (nx5078), .A (D[181])) ;
    tri01 tri_F_182 (.Y (F[182]), .A (nx5081), .E (nx5937)) ;
    inv01 ix5082 (.Y (nx5081), .A (D[182])) ;
    tri01 tri_F_183 (.Y (F[183]), .A (nx5084), .E (nx5937)) ;
    inv01 ix5085 (.Y (nx5084), .A (D[183])) ;
    tri01 tri_F_184 (.Y (F[184]), .A (nx5087), .E (nx5937)) ;
    inv01 ix5088 (.Y (nx5087), .A (D[184])) ;
    tri01 tri_F_185 (.Y (F[185]), .A (nx5090), .E (nx5937)) ;
    inv01 ix5091 (.Y (nx5090), .A (D[185])) ;
    tri01 tri_F_186 (.Y (F[186]), .A (nx5093), .E (nx5937)) ;
    inv01 ix5094 (.Y (nx5093), .A (D[186])) ;
    tri01 tri_F_187 (.Y (F[187]), .A (nx5096), .E (nx5937)) ;
    inv01 ix5097 (.Y (nx5096), .A (D[187])) ;
    tri01 tri_F_188 (.Y (F[188]), .A (nx5099), .E (nx5937)) ;
    inv01 ix5100 (.Y (nx5099), .A (D[188])) ;
    tri01 tri_F_189 (.Y (F[189]), .A (nx5102), .E (nx5939)) ;
    inv01 ix5103 (.Y (nx5102), .A (D[189])) ;
    tri01 tri_F_190 (.Y (F[190]), .A (nx5105), .E (nx5939)) ;
    inv01 ix5106 (.Y (nx5105), .A (D[190])) ;
    tri01 tri_F_191 (.Y (F[191]), .A (nx5108), .E (nx5939)) ;
    inv01 ix5109 (.Y (nx5108), .A (D[191])) ;
    tri01 tri_F_192 (.Y (F[192]), .A (nx5111), .E (nx5939)) ;
    inv01 ix5112 (.Y (nx5111), .A (D[192])) ;
    tri01 tri_F_193 (.Y (F[193]), .A (nx5114), .E (nx5939)) ;
    inv01 ix5115 (.Y (nx5114), .A (D[193])) ;
    tri01 tri_F_194 (.Y (F[194]), .A (nx5117), .E (nx5939)) ;
    inv01 ix5118 (.Y (nx5117), .A (D[194])) ;
    tri01 tri_F_195 (.Y (F[195]), .A (nx5120), .E (nx5939)) ;
    inv01 ix5121 (.Y (nx5120), .A (D[195])) ;
    tri01 tri_F_196 (.Y (F[196]), .A (nx5123), .E (nx5941)) ;
    inv01 ix5124 (.Y (nx5123), .A (D[196])) ;
    tri01 tri_F_197 (.Y (F[197]), .A (nx5126), .E (nx5941)) ;
    inv01 ix5127 (.Y (nx5126), .A (D[197])) ;
    tri01 tri_F_198 (.Y (F[198]), .A (nx5129), .E (nx5941)) ;
    inv01 ix5130 (.Y (nx5129), .A (D[198])) ;
    tri01 tri_F_199 (.Y (F[199]), .A (nx5132), .E (nx5941)) ;
    inv01 ix5133 (.Y (nx5132), .A (D[199])) ;
    tri01 tri_F_200 (.Y (F[200]), .A (nx5135), .E (nx5941)) ;
    inv01 ix5136 (.Y (nx5135), .A (D[200])) ;
    tri01 tri_F_201 (.Y (F[201]), .A (nx5138), .E (nx5941)) ;
    inv01 ix5139 (.Y (nx5138), .A (D[201])) ;
    tri01 tri_F_202 (.Y (F[202]), .A (nx5141), .E (nx5941)) ;
    inv01 ix5142 (.Y (nx5141), .A (D[202])) ;
    tri01 tri_F_203 (.Y (F[203]), .A (nx5144), .E (nx5943)) ;
    inv01 ix5145 (.Y (nx5144), .A (D[203])) ;
    tri01 tri_F_204 (.Y (F[204]), .A (nx5147), .E (nx5943)) ;
    inv01 ix5148 (.Y (nx5147), .A (D[204])) ;
    tri01 tri_F_205 (.Y (F[205]), .A (nx5150), .E (nx5943)) ;
    inv01 ix5151 (.Y (nx5150), .A (D[205])) ;
    tri01 tri_F_206 (.Y (F[206]), .A (nx5153), .E (nx5943)) ;
    inv01 ix5154 (.Y (nx5153), .A (D[206])) ;
    tri01 tri_F_207 (.Y (F[207]), .A (nx5156), .E (nx5943)) ;
    inv01 ix5157 (.Y (nx5156), .A (D[207])) ;
    tri01 tri_F_208 (.Y (F[208]), .A (nx5159), .E (nx5943)) ;
    inv01 ix5160 (.Y (nx5159), .A (D[208])) ;
    tri01 tri_F_209 (.Y (F[209]), .A (nx5162), .E (nx5943)) ;
    inv01 ix5163 (.Y (nx5162), .A (D[209])) ;
    tri01 tri_F_210 (.Y (F[210]), .A (nx5165), .E (nx5945)) ;
    inv01 ix5166 (.Y (nx5165), .A (D[210])) ;
    tri01 tri_F_211 (.Y (F[211]), .A (nx5168), .E (nx5945)) ;
    inv01 ix5169 (.Y (nx5168), .A (D[211])) ;
    tri01 tri_F_212 (.Y (F[212]), .A (nx5171), .E (nx5945)) ;
    inv01 ix5172 (.Y (nx5171), .A (D[212])) ;
    tri01 tri_F_213 (.Y (F[213]), .A (nx5174), .E (nx5945)) ;
    inv01 ix5175 (.Y (nx5174), .A (D[213])) ;
    tri01 tri_F_214 (.Y (F[214]), .A (nx5177), .E (nx5945)) ;
    inv01 ix5178 (.Y (nx5177), .A (D[214])) ;
    tri01 tri_F_215 (.Y (F[215]), .A (nx5180), .E (nx5945)) ;
    inv01 ix5181 (.Y (nx5180), .A (D[215])) ;
    tri01 tri_F_216 (.Y (F[216]), .A (nx5183), .E (nx5945)) ;
    inv01 ix5184 (.Y (nx5183), .A (D[216])) ;
    tri01 tri_F_217 (.Y (F[217]), .A (nx5186), .E (nx5947)) ;
    inv01 ix5187 (.Y (nx5186), .A (D[217])) ;
    tri01 tri_F_218 (.Y (F[218]), .A (nx5189), .E (nx5947)) ;
    inv01 ix5190 (.Y (nx5189), .A (D[218])) ;
    tri01 tri_F_219 (.Y (F[219]), .A (nx5192), .E (nx5947)) ;
    inv01 ix5193 (.Y (nx5192), .A (D[219])) ;
    tri01 tri_F_220 (.Y (F[220]), .A (nx5195), .E (nx5947)) ;
    inv01 ix5196 (.Y (nx5195), .A (D[220])) ;
    tri01 tri_F_221 (.Y (F[221]), .A (nx5198), .E (nx5947)) ;
    inv01 ix5199 (.Y (nx5198), .A (D[221])) ;
    tri01 tri_F_222 (.Y (F[222]), .A (nx5201), .E (nx5947)) ;
    inv01 ix5202 (.Y (nx5201), .A (D[222])) ;
    tri01 tri_F_223 (.Y (F[223]), .A (nx5204), .E (nx5947)) ;
    inv01 ix5205 (.Y (nx5204), .A (D[223])) ;
    tri01 tri_F_224 (.Y (F[224]), .A (nx5207), .E (nx5949)) ;
    inv01 ix5208 (.Y (nx5207), .A (D[224])) ;
    tri01 tri_F_225 (.Y (F[225]), .A (nx5210), .E (nx5949)) ;
    inv01 ix5211 (.Y (nx5210), .A (D[225])) ;
    tri01 tri_F_226 (.Y (F[226]), .A (nx5213), .E (nx5949)) ;
    inv01 ix5214 (.Y (nx5213), .A (D[226])) ;
    tri01 tri_F_227 (.Y (F[227]), .A (nx5216), .E (nx5949)) ;
    inv01 ix5217 (.Y (nx5216), .A (D[227])) ;
    tri01 tri_F_228 (.Y (F[228]), .A (nx5219), .E (nx5949)) ;
    inv01 ix5220 (.Y (nx5219), .A (D[228])) ;
    tri01 tri_F_229 (.Y (F[229]), .A (nx5222), .E (nx5949)) ;
    inv01 ix5223 (.Y (nx5222), .A (D[229])) ;
    tri01 tri_F_230 (.Y (F[230]), .A (nx5225), .E (nx5949)) ;
    inv01 ix5226 (.Y (nx5225), .A (D[230])) ;
    tri01 tri_F_231 (.Y (F[231]), .A (nx5228), .E (nx5951)) ;
    inv01 ix5229 (.Y (nx5228), .A (D[231])) ;
    tri01 tri_F_232 (.Y (F[232]), .A (nx5231), .E (nx5951)) ;
    inv01 ix5232 (.Y (nx5231), .A (D[232])) ;
    tri01 tri_F_233 (.Y (F[233]), .A (nx5234), .E (nx5951)) ;
    inv01 ix5235 (.Y (nx5234), .A (D[233])) ;
    tri01 tri_F_234 (.Y (F[234]), .A (nx5237), .E (nx5951)) ;
    inv01 ix5238 (.Y (nx5237), .A (D[234])) ;
    tri01 tri_F_235 (.Y (F[235]), .A (nx5240), .E (nx5951)) ;
    inv01 ix5241 (.Y (nx5240), .A (D[235])) ;
    tri01 tri_F_236 (.Y (F[236]), .A (nx5243), .E (nx5951)) ;
    inv01 ix5244 (.Y (nx5243), .A (D[236])) ;
    tri01 tri_F_237 (.Y (F[237]), .A (nx5246), .E (nx5951)) ;
    inv01 ix5247 (.Y (nx5246), .A (D[237])) ;
    tri01 tri_F_238 (.Y (F[238]), .A (nx5249), .E (nx5953)) ;
    inv01 ix5250 (.Y (nx5249), .A (D[238])) ;
    tri01 tri_F_239 (.Y (F[239]), .A (nx5252), .E (nx5953)) ;
    inv01 ix5253 (.Y (nx5252), .A (D[239])) ;
    tri01 tri_F_240 (.Y (F[240]), .A (nx5255), .E (nx5953)) ;
    inv01 ix5256 (.Y (nx5255), .A (D[240])) ;
    tri01 tri_F_241 (.Y (F[241]), .A (nx5258), .E (nx5953)) ;
    inv01 ix5259 (.Y (nx5258), .A (D[241])) ;
    tri01 tri_F_242 (.Y (F[242]), .A (nx5261), .E (nx5953)) ;
    inv01 ix5262 (.Y (nx5261), .A (D[242])) ;
    tri01 tri_F_243 (.Y (F[243]), .A (nx5264), .E (nx5953)) ;
    inv01 ix5265 (.Y (nx5264), .A (D[243])) ;
    tri01 tri_F_244 (.Y (F[244]), .A (nx5267), .E (nx5953)) ;
    inv01 ix5268 (.Y (nx5267), .A (D[244])) ;
    tri01 tri_F_245 (.Y (F[245]), .A (nx5270), .E (nx5955)) ;
    inv01 ix5271 (.Y (nx5270), .A (D[245])) ;
    tri01 tri_F_246 (.Y (F[246]), .A (nx5273), .E (nx5955)) ;
    inv01 ix5274 (.Y (nx5273), .A (D[246])) ;
    tri01 tri_F_247 (.Y (F[247]), .A (nx5276), .E (nx5955)) ;
    inv01 ix5277 (.Y (nx5276), .A (D[247])) ;
    tri01 tri_F_248 (.Y (F[248]), .A (nx5279), .E (nx5955)) ;
    inv01 ix5280 (.Y (nx5279), .A (D[248])) ;
    tri01 tri_F_249 (.Y (F[249]), .A (nx5282), .E (nx5955)) ;
    inv01 ix5283 (.Y (nx5282), .A (D[249])) ;
    tri01 tri_F_250 (.Y (F[250]), .A (nx5285), .E (nx5955)) ;
    inv01 ix5286 (.Y (nx5285), .A (D[250])) ;
    tri01 tri_F_251 (.Y (F[251]), .A (nx5288), .E (nx5955)) ;
    inv01 ix5289 (.Y (nx5288), .A (D[251])) ;
    tri01 tri_F_252 (.Y (F[252]), .A (nx5291), .E (nx5957)) ;
    inv01 ix5292 (.Y (nx5291), .A (D[252])) ;
    tri01 tri_F_253 (.Y (F[253]), .A (nx5294), .E (nx5957)) ;
    inv01 ix5295 (.Y (nx5294), .A (D[253])) ;
    tri01 tri_F_254 (.Y (F[254]), .A (nx5297), .E (nx5957)) ;
    inv01 ix5298 (.Y (nx5297), .A (D[254])) ;
    tri01 tri_F_255 (.Y (F[255]), .A (nx5300), .E (nx5957)) ;
    inv01 ix5301 (.Y (nx5300), .A (D[255])) ;
    tri01 tri_F_256 (.Y (F[256]), .A (nx5303), .E (nx5957)) ;
    inv01 ix5304 (.Y (nx5303), .A (D[256])) ;
    tri01 tri_F_257 (.Y (F[257]), .A (nx5306), .E (nx5957)) ;
    inv01 ix5307 (.Y (nx5306), .A (D[257])) ;
    tri01 tri_F_258 (.Y (F[258]), .A (nx5309), .E (nx5957)) ;
    inv01 ix5310 (.Y (nx5309), .A (D[258])) ;
    tri01 tri_F_259 (.Y (F[259]), .A (nx5312), .E (nx5959)) ;
    inv01 ix5313 (.Y (nx5312), .A (D[259])) ;
    tri01 tri_F_260 (.Y (F[260]), .A (nx5315), .E (nx5959)) ;
    inv01 ix5316 (.Y (nx5315), .A (D[260])) ;
    tri01 tri_F_261 (.Y (F[261]), .A (nx5318), .E (nx5959)) ;
    inv01 ix5319 (.Y (nx5318), .A (D[261])) ;
    tri01 tri_F_262 (.Y (F[262]), .A (nx5321), .E (nx5959)) ;
    inv01 ix5322 (.Y (nx5321), .A (D[262])) ;
    tri01 tri_F_263 (.Y (F[263]), .A (nx5324), .E (nx5959)) ;
    inv01 ix5325 (.Y (nx5324), .A (D[263])) ;
    tri01 tri_F_264 (.Y (F[264]), .A (nx5327), .E (nx5959)) ;
    inv01 ix5328 (.Y (nx5327), .A (D[264])) ;
    tri01 tri_F_265 (.Y (F[265]), .A (nx5330), .E (nx5959)) ;
    inv01 ix5331 (.Y (nx5330), .A (D[265])) ;
    tri01 tri_F_266 (.Y (F[266]), .A (nx5333), .E (nx5961)) ;
    inv01 ix5334 (.Y (nx5333), .A (D[266])) ;
    tri01 tri_F_267 (.Y (F[267]), .A (nx5336), .E (nx5961)) ;
    inv01 ix5337 (.Y (nx5336), .A (D[267])) ;
    tri01 tri_F_268 (.Y (F[268]), .A (nx5339), .E (nx5961)) ;
    inv01 ix5340 (.Y (nx5339), .A (D[268])) ;
    tri01 tri_F_269 (.Y (F[269]), .A (nx5342), .E (nx5961)) ;
    inv01 ix5343 (.Y (nx5342), .A (D[269])) ;
    tri01 tri_F_270 (.Y (F[270]), .A (nx5345), .E (nx5961)) ;
    inv01 ix5346 (.Y (nx5345), .A (D[270])) ;
    tri01 tri_F_271 (.Y (F[271]), .A (nx5348), .E (nx5961)) ;
    inv01 ix5349 (.Y (nx5348), .A (D[271])) ;
    tri01 tri_F_272 (.Y (F[272]), .A (nx5351), .E (nx5961)) ;
    inv01 ix5352 (.Y (nx5351), .A (D[272])) ;
    tri01 tri_F_273 (.Y (F[273]), .A (nx5354), .E (nx5963)) ;
    inv01 ix5355 (.Y (nx5354), .A (D[273])) ;
    tri01 tri_F_274 (.Y (F[274]), .A (nx5357), .E (nx5963)) ;
    inv01 ix5358 (.Y (nx5357), .A (D[274])) ;
    tri01 tri_F_275 (.Y (F[275]), .A (nx5360), .E (nx5963)) ;
    inv01 ix5361 (.Y (nx5360), .A (D[275])) ;
    tri01 tri_F_276 (.Y (F[276]), .A (nx5363), .E (nx5963)) ;
    inv01 ix5364 (.Y (nx5363), .A (D[276])) ;
    tri01 tri_F_277 (.Y (F[277]), .A (nx5366), .E (nx5963)) ;
    inv01 ix5367 (.Y (nx5366), .A (D[277])) ;
    tri01 tri_F_278 (.Y (F[278]), .A (nx5369), .E (nx5963)) ;
    inv01 ix5370 (.Y (nx5369), .A (D[278])) ;
    tri01 tri_F_279 (.Y (F[279]), .A (nx5372), .E (nx5963)) ;
    inv01 ix5373 (.Y (nx5372), .A (D[279])) ;
    tri01 tri_F_280 (.Y (F[280]), .A (nx5375), .E (nx5965)) ;
    inv01 ix5376 (.Y (nx5375), .A (D[280])) ;
    tri01 tri_F_281 (.Y (F[281]), .A (nx5378), .E (nx5965)) ;
    inv01 ix5379 (.Y (nx5378), .A (D[281])) ;
    tri01 tri_F_282 (.Y (F[282]), .A (nx5381), .E (nx5965)) ;
    inv01 ix5382 (.Y (nx5381), .A (D[282])) ;
    tri01 tri_F_283 (.Y (F[283]), .A (nx5384), .E (nx5965)) ;
    inv01 ix5385 (.Y (nx5384), .A (D[283])) ;
    tri01 tri_F_284 (.Y (F[284]), .A (nx5387), .E (nx5965)) ;
    inv01 ix5388 (.Y (nx5387), .A (D[284])) ;
    tri01 tri_F_285 (.Y (F[285]), .A (nx5390), .E (nx5965)) ;
    inv01 ix5391 (.Y (nx5390), .A (D[285])) ;
    tri01 tri_F_286 (.Y (F[286]), .A (nx5393), .E (nx5965)) ;
    inv01 ix5394 (.Y (nx5393), .A (D[286])) ;
    tri01 tri_F_287 (.Y (F[287]), .A (nx5396), .E (nx5967)) ;
    inv01 ix5397 (.Y (nx5396), .A (D[287])) ;
    tri01 tri_F_288 (.Y (F[288]), .A (nx5399), .E (nx5967)) ;
    inv01 ix5400 (.Y (nx5399), .A (D[288])) ;
    tri01 tri_F_289 (.Y (F[289]), .A (nx5402), .E (nx5967)) ;
    inv01 ix5403 (.Y (nx5402), .A (D[289])) ;
    tri01 tri_F_290 (.Y (F[290]), .A (nx5405), .E (nx5967)) ;
    inv01 ix5406 (.Y (nx5405), .A (D[290])) ;
    tri01 tri_F_291 (.Y (F[291]), .A (nx5408), .E (nx5967)) ;
    inv01 ix5409 (.Y (nx5408), .A (D[291])) ;
    tri01 tri_F_292 (.Y (F[292]), .A (nx5411), .E (nx5967)) ;
    inv01 ix5412 (.Y (nx5411), .A (D[292])) ;
    tri01 tri_F_293 (.Y (F[293]), .A (nx5414), .E (nx5967)) ;
    inv01 ix5415 (.Y (nx5414), .A (D[293])) ;
    tri01 tri_F_294 (.Y (F[294]), .A (nx5417), .E (nx5969)) ;
    inv01 ix5418 (.Y (nx5417), .A (D[294])) ;
    tri01 tri_F_295 (.Y (F[295]), .A (nx5420), .E (nx5969)) ;
    inv01 ix5421 (.Y (nx5420), .A (D[295])) ;
    tri01 tri_F_296 (.Y (F[296]), .A (nx5423), .E (nx5969)) ;
    inv01 ix5424 (.Y (nx5423), .A (D[296])) ;
    tri01 tri_F_297 (.Y (F[297]), .A (nx5426), .E (nx5969)) ;
    inv01 ix5427 (.Y (nx5426), .A (D[297])) ;
    tri01 tri_F_298 (.Y (F[298]), .A (nx5429), .E (nx5969)) ;
    inv01 ix5430 (.Y (nx5429), .A (D[298])) ;
    tri01 tri_F_299 (.Y (F[299]), .A (nx5432), .E (nx5969)) ;
    inv01 ix5433 (.Y (nx5432), .A (D[299])) ;
    tri01 tri_F_300 (.Y (F[300]), .A (nx5435), .E (nx5969)) ;
    inv01 ix5436 (.Y (nx5435), .A (D[300])) ;
    tri01 tri_F_301 (.Y (F[301]), .A (nx5438), .E (nx5971)) ;
    inv01 ix5439 (.Y (nx5438), .A (D[301])) ;
    tri01 tri_F_302 (.Y (F[302]), .A (nx5441), .E (nx5971)) ;
    inv01 ix5442 (.Y (nx5441), .A (D[302])) ;
    tri01 tri_F_303 (.Y (F[303]), .A (nx5444), .E (nx5971)) ;
    inv01 ix5445 (.Y (nx5444), .A (D[303])) ;
    tri01 tri_F_304 (.Y (F[304]), .A (nx5447), .E (nx5971)) ;
    inv01 ix5448 (.Y (nx5447), .A (D[304])) ;
    tri01 tri_F_305 (.Y (F[305]), .A (nx5450), .E (nx5971)) ;
    inv01 ix5451 (.Y (nx5450), .A (D[305])) ;
    tri01 tri_F_306 (.Y (F[306]), .A (nx5453), .E (nx5971)) ;
    inv01 ix5454 (.Y (nx5453), .A (D[306])) ;
    tri01 tri_F_307 (.Y (F[307]), .A (nx5456), .E (nx5971)) ;
    inv01 ix5457 (.Y (nx5456), .A (D[307])) ;
    tri01 tri_F_308 (.Y (F[308]), .A (nx5459), .E (nx5973)) ;
    inv01 ix5460 (.Y (nx5459), .A (D[308])) ;
    tri01 tri_F_309 (.Y (F[309]), .A (nx5462), .E (nx5973)) ;
    inv01 ix5463 (.Y (nx5462), .A (D[309])) ;
    tri01 tri_F_310 (.Y (F[310]), .A (nx5465), .E (nx5973)) ;
    inv01 ix5466 (.Y (nx5465), .A (D[310])) ;
    tri01 tri_F_311 (.Y (F[311]), .A (nx5468), .E (nx5973)) ;
    inv01 ix5469 (.Y (nx5468), .A (D[311])) ;
    tri01 tri_F_312 (.Y (F[312]), .A (nx5471), .E (nx5973)) ;
    inv01 ix5472 (.Y (nx5471), .A (D[312])) ;
    tri01 tri_F_313 (.Y (F[313]), .A (nx5474), .E (nx5973)) ;
    inv01 ix5475 (.Y (nx5474), .A (D[313])) ;
    tri01 tri_F_314 (.Y (F[314]), .A (nx5477), .E (nx5973)) ;
    inv01 ix5478 (.Y (nx5477), .A (D[314])) ;
    tri01 tri_F_315 (.Y (F[315]), .A (nx5480), .E (nx5975)) ;
    inv01 ix5481 (.Y (nx5480), .A (D[315])) ;
    tri01 tri_F_316 (.Y (F[316]), .A (nx5483), .E (nx5975)) ;
    inv01 ix5484 (.Y (nx5483), .A (D[316])) ;
    tri01 tri_F_317 (.Y (F[317]), .A (nx5486), .E (nx5975)) ;
    inv01 ix5487 (.Y (nx5486), .A (D[317])) ;
    tri01 tri_F_318 (.Y (F[318]), .A (nx5489), .E (nx5975)) ;
    inv01 ix5490 (.Y (nx5489), .A (D[318])) ;
    tri01 tri_F_319 (.Y (F[319]), .A (nx5492), .E (nx5975)) ;
    inv01 ix5493 (.Y (nx5492), .A (D[319])) ;
    tri01 tri_F_320 (.Y (F[320]), .A (nx5495), .E (nx5975)) ;
    inv01 ix5496 (.Y (nx5495), .A (D[320])) ;
    tri01 tri_F_321 (.Y (F[321]), .A (nx5498), .E (nx5975)) ;
    inv01 ix5499 (.Y (nx5498), .A (D[321])) ;
    tri01 tri_F_322 (.Y (F[322]), .A (nx5501), .E (nx5977)) ;
    inv01 ix5502 (.Y (nx5501), .A (D[322])) ;
    tri01 tri_F_323 (.Y (F[323]), .A (nx5504), .E (nx5977)) ;
    inv01 ix5505 (.Y (nx5504), .A (D[323])) ;
    tri01 tri_F_324 (.Y (F[324]), .A (nx5507), .E (nx5977)) ;
    inv01 ix5508 (.Y (nx5507), .A (D[324])) ;
    tri01 tri_F_325 (.Y (F[325]), .A (nx5510), .E (nx5977)) ;
    inv01 ix5511 (.Y (nx5510), .A (D[325])) ;
    tri01 tri_F_326 (.Y (F[326]), .A (nx5513), .E (nx5977)) ;
    inv01 ix5514 (.Y (nx5513), .A (D[326])) ;
    tri01 tri_F_327 (.Y (F[327]), .A (nx5516), .E (nx5977)) ;
    inv01 ix5517 (.Y (nx5516), .A (D[327])) ;
    tri01 tri_F_328 (.Y (F[328]), .A (nx5519), .E (nx5977)) ;
    inv01 ix5520 (.Y (nx5519), .A (D[328])) ;
    tri01 tri_F_329 (.Y (F[329]), .A (nx5522), .E (nx5979)) ;
    inv01 ix5523 (.Y (nx5522), .A (D[329])) ;
    tri01 tri_F_330 (.Y (F[330]), .A (nx5525), .E (nx5979)) ;
    inv01 ix5526 (.Y (nx5525), .A (D[330])) ;
    tri01 tri_F_331 (.Y (F[331]), .A (nx5528), .E (nx5979)) ;
    inv01 ix5529 (.Y (nx5528), .A (D[331])) ;
    tri01 tri_F_332 (.Y (F[332]), .A (nx5531), .E (nx5979)) ;
    inv01 ix5532 (.Y (nx5531), .A (D[332])) ;
    tri01 tri_F_333 (.Y (F[333]), .A (nx5534), .E (nx5979)) ;
    inv01 ix5535 (.Y (nx5534), .A (D[333])) ;
    tri01 tri_F_334 (.Y (F[334]), .A (nx5537), .E (nx5979)) ;
    inv01 ix5538 (.Y (nx5537), .A (D[334])) ;
    tri01 tri_F_335 (.Y (F[335]), .A (nx5540), .E (nx5979)) ;
    inv01 ix5541 (.Y (nx5540), .A (D[335])) ;
    tri01 tri_F_336 (.Y (F[336]), .A (nx5543), .E (nx5981)) ;
    inv01 ix5544 (.Y (nx5543), .A (D[336])) ;
    tri01 tri_F_337 (.Y (F[337]), .A (nx5546), .E (nx5981)) ;
    inv01 ix5547 (.Y (nx5546), .A (D[337])) ;
    tri01 tri_F_338 (.Y (F[338]), .A (nx5549), .E (nx5981)) ;
    inv01 ix5550 (.Y (nx5549), .A (D[338])) ;
    tri01 tri_F_339 (.Y (F[339]), .A (nx5552), .E (nx5981)) ;
    inv01 ix5553 (.Y (nx5552), .A (D[339])) ;
    tri01 tri_F_340 (.Y (F[340]), .A (nx5555), .E (nx5981)) ;
    inv01 ix5556 (.Y (nx5555), .A (D[340])) ;
    tri01 tri_F_341 (.Y (F[341]), .A (nx5558), .E (nx5981)) ;
    inv01 ix5559 (.Y (nx5558), .A (D[341])) ;
    tri01 tri_F_342 (.Y (F[342]), .A (nx5561), .E (nx5981)) ;
    inv01 ix5562 (.Y (nx5561), .A (D[342])) ;
    tri01 tri_F_343 (.Y (F[343]), .A (nx5564), .E (nx5983)) ;
    inv01 ix5565 (.Y (nx5564), .A (D[343])) ;
    tri01 tri_F_344 (.Y (F[344]), .A (nx5567), .E (nx5983)) ;
    inv01 ix5568 (.Y (nx5567), .A (D[344])) ;
    tri01 tri_F_345 (.Y (F[345]), .A (nx5570), .E (nx5983)) ;
    inv01 ix5571 (.Y (nx5570), .A (D[345])) ;
    tri01 tri_F_346 (.Y (F[346]), .A (nx5573), .E (nx5983)) ;
    inv01 ix5574 (.Y (nx5573), .A (D[346])) ;
    tri01 tri_F_347 (.Y (F[347]), .A (nx5576), .E (nx5983)) ;
    inv01 ix5577 (.Y (nx5576), .A (D[347])) ;
    tri01 tri_F_348 (.Y (F[348]), .A (nx5579), .E (nx5983)) ;
    inv01 ix5580 (.Y (nx5579), .A (D[348])) ;
    tri01 tri_F_349 (.Y (F[349]), .A (nx5582), .E (nx5983)) ;
    inv01 ix5583 (.Y (nx5582), .A (D[349])) ;
    tri01 tri_F_350 (.Y (F[350]), .A (nx5585), .E (nx5985)) ;
    inv01 ix5586 (.Y (nx5585), .A (D[350])) ;
    tri01 tri_F_351 (.Y (F[351]), .A (nx5588), .E (nx5985)) ;
    inv01 ix5589 (.Y (nx5588), .A (D[351])) ;
    tri01 tri_F_352 (.Y (F[352]), .A (nx5591), .E (nx5985)) ;
    inv01 ix5592 (.Y (nx5591), .A (D[352])) ;
    tri01 tri_F_353 (.Y (F[353]), .A (nx5594), .E (nx5985)) ;
    inv01 ix5595 (.Y (nx5594), .A (D[353])) ;
    tri01 tri_F_354 (.Y (F[354]), .A (nx5597), .E (nx5985)) ;
    inv01 ix5598 (.Y (nx5597), .A (D[354])) ;
    tri01 tri_F_355 (.Y (F[355]), .A (nx5600), .E (nx5985)) ;
    inv01 ix5601 (.Y (nx5600), .A (D[355])) ;
    tri01 tri_F_356 (.Y (F[356]), .A (nx5603), .E (nx5985)) ;
    inv01 ix5604 (.Y (nx5603), .A (D[356])) ;
    tri01 tri_F_357 (.Y (F[357]), .A (nx5606), .E (nx5987)) ;
    inv01 ix5607 (.Y (nx5606), .A (D[357])) ;
    tri01 tri_F_358 (.Y (F[358]), .A (nx5609), .E (nx5987)) ;
    inv01 ix5610 (.Y (nx5609), .A (D[358])) ;
    tri01 tri_F_359 (.Y (F[359]), .A (nx5612), .E (nx5987)) ;
    inv01 ix5613 (.Y (nx5612), .A (D[359])) ;
    tri01 tri_F_360 (.Y (F[360]), .A (nx5615), .E (nx5987)) ;
    inv01 ix5616 (.Y (nx5615), .A (D[360])) ;
    tri01 tri_F_361 (.Y (F[361]), .A (nx5618), .E (nx5987)) ;
    inv01 ix5619 (.Y (nx5618), .A (D[361])) ;
    tri01 tri_F_362 (.Y (F[362]), .A (nx5621), .E (nx5987)) ;
    inv01 ix5622 (.Y (nx5621), .A (D[362])) ;
    tri01 tri_F_363 (.Y (F[363]), .A (nx5624), .E (nx5987)) ;
    inv01 ix5625 (.Y (nx5624), .A (D[363])) ;
    tri01 tri_F_364 (.Y (F[364]), .A (nx5627), .E (nx5989)) ;
    inv01 ix5628 (.Y (nx5627), .A (D[364])) ;
    tri01 tri_F_365 (.Y (F[365]), .A (nx5630), .E (nx5989)) ;
    inv01 ix5631 (.Y (nx5630), .A (D[365])) ;
    tri01 tri_F_366 (.Y (F[366]), .A (nx5633), .E (nx5989)) ;
    inv01 ix5634 (.Y (nx5633), .A (D[366])) ;
    tri01 tri_F_367 (.Y (F[367]), .A (nx5636), .E (nx5989)) ;
    inv01 ix5637 (.Y (nx5636), .A (D[367])) ;
    tri01 tri_F_368 (.Y (F[368]), .A (nx5639), .E (nx5989)) ;
    inv01 ix5640 (.Y (nx5639), .A (D[368])) ;
    tri01 tri_F_369 (.Y (F[369]), .A (nx5642), .E (nx5989)) ;
    inv01 ix5643 (.Y (nx5642), .A (D[369])) ;
    tri01 tri_F_370 (.Y (F[370]), .A (nx5645), .E (nx5989)) ;
    inv01 ix5646 (.Y (nx5645), .A (D[370])) ;
    tri01 tri_F_371 (.Y (F[371]), .A (nx5648), .E (nx5991)) ;
    inv01 ix5649 (.Y (nx5648), .A (D[371])) ;
    tri01 tri_F_372 (.Y (F[372]), .A (nx5651), .E (nx5991)) ;
    inv01 ix5652 (.Y (nx5651), .A (D[372])) ;
    tri01 tri_F_373 (.Y (F[373]), .A (nx5654), .E (nx5991)) ;
    inv01 ix5655 (.Y (nx5654), .A (D[373])) ;
    tri01 tri_F_374 (.Y (F[374]), .A (nx5657), .E (nx5991)) ;
    inv01 ix5658 (.Y (nx5657), .A (D[374])) ;
    tri01 tri_F_375 (.Y (F[375]), .A (nx5660), .E (nx5991)) ;
    inv01 ix5661 (.Y (nx5660), .A (D[375])) ;
    tri01 tri_F_376 (.Y (F[376]), .A (nx5663), .E (nx5991)) ;
    inv01 ix5664 (.Y (nx5663), .A (D[376])) ;
    tri01 tri_F_377 (.Y (F[377]), .A (nx5666), .E (nx5991)) ;
    inv01 ix5667 (.Y (nx5666), .A (D[377])) ;
    tri01 tri_F_378 (.Y (F[378]), .A (nx5669), .E (nx5993)) ;
    inv01 ix5670 (.Y (nx5669), .A (D[378])) ;
    tri01 tri_F_379 (.Y (F[379]), .A (nx5672), .E (nx5993)) ;
    inv01 ix5673 (.Y (nx5672), .A (D[379])) ;
    tri01 tri_F_380 (.Y (F[380]), .A (nx5675), .E (nx5993)) ;
    inv01 ix5676 (.Y (nx5675), .A (D[380])) ;
    tri01 tri_F_381 (.Y (F[381]), .A (nx5678), .E (nx5993)) ;
    inv01 ix5679 (.Y (nx5678), .A (D[381])) ;
    tri01 tri_F_382 (.Y (F[382]), .A (nx5681), .E (nx5993)) ;
    inv01 ix5682 (.Y (nx5681), .A (D[382])) ;
    tri01 tri_F_383 (.Y (F[383]), .A (nx5684), .E (nx5993)) ;
    inv01 ix5685 (.Y (nx5684), .A (D[383])) ;
    tri01 tri_F_384 (.Y (F[384]), .A (nx5687), .E (nx5993)) ;
    inv01 ix5688 (.Y (nx5687), .A (D[384])) ;
    tri01 tri_F_385 (.Y (F[385]), .A (nx5690), .E (nx5995)) ;
    inv01 ix5691 (.Y (nx5690), .A (D[385])) ;
    tri01 tri_F_386 (.Y (F[386]), .A (nx5693), .E (nx5995)) ;
    inv01 ix5694 (.Y (nx5693), .A (D[386])) ;
    tri01 tri_F_387 (.Y (F[387]), .A (nx5696), .E (nx5995)) ;
    inv01 ix5697 (.Y (nx5696), .A (D[387])) ;
    tri01 tri_F_388 (.Y (F[388]), .A (nx5699), .E (nx5995)) ;
    inv01 ix5700 (.Y (nx5699), .A (D[388])) ;
    tri01 tri_F_389 (.Y (F[389]), .A (nx5702), .E (nx5995)) ;
    inv01 ix5703 (.Y (nx5702), .A (D[389])) ;
    tri01 tri_F_390 (.Y (F[390]), .A (nx5705), .E (nx5995)) ;
    inv01 ix5706 (.Y (nx5705), .A (D[390])) ;
    tri01 tri_F_391 (.Y (F[391]), .A (nx5708), .E (nx5995)) ;
    inv01 ix5709 (.Y (nx5708), .A (D[391])) ;
    tri01 tri_F_392 (.Y (F[392]), .A (nx5711), .E (nx5997)) ;
    inv01 ix5712 (.Y (nx5711), .A (D[392])) ;
    tri01 tri_F_393 (.Y (F[393]), .A (nx5714), .E (nx5997)) ;
    inv01 ix5715 (.Y (nx5714), .A (D[393])) ;
    tri01 tri_F_394 (.Y (F[394]), .A (nx5717), .E (nx5997)) ;
    inv01 ix5718 (.Y (nx5717), .A (D[394])) ;
    tri01 tri_F_395 (.Y (F[395]), .A (nx5720), .E (nx5997)) ;
    inv01 ix5721 (.Y (nx5720), .A (D[395])) ;
    tri01 tri_F_396 (.Y (F[396]), .A (nx5723), .E (nx5997)) ;
    inv01 ix5724 (.Y (nx5723), .A (D[396])) ;
    tri01 tri_F_397 (.Y (F[397]), .A (nx5726), .E (nx5997)) ;
    inv01 ix5727 (.Y (nx5726), .A (D[397])) ;
    tri01 tri_F_398 (.Y (F[398]), .A (nx5729), .E (nx5997)) ;
    inv01 ix5730 (.Y (nx5729), .A (D[398])) ;
    tri01 tri_F_399 (.Y (F[399]), .A (nx5732), .E (nx5999)) ;
    inv01 ix5733 (.Y (nx5732), .A (D[399])) ;
    tri01 tri_F_400 (.Y (F[400]), .A (nx5735), .E (nx5999)) ;
    inv01 ix5736 (.Y (nx5735), .A (D[400])) ;
    tri01 tri_F_401 (.Y (F[401]), .A (nx5738), .E (nx5999)) ;
    inv01 ix5739 (.Y (nx5738), .A (D[401])) ;
    tri01 tri_F_402 (.Y (F[402]), .A (nx5741), .E (nx5999)) ;
    inv01 ix5742 (.Y (nx5741), .A (D[402])) ;
    tri01 tri_F_403 (.Y (F[403]), .A (nx5744), .E (nx5999)) ;
    inv01 ix5745 (.Y (nx5744), .A (D[403])) ;
    tri01 tri_F_404 (.Y (F[404]), .A (nx5747), .E (nx5999)) ;
    inv01 ix5748 (.Y (nx5747), .A (D[404])) ;
    tri01 tri_F_405 (.Y (F[405]), .A (nx5750), .E (nx5999)) ;
    inv01 ix5751 (.Y (nx5750), .A (D[405])) ;
    tri01 tri_F_406 (.Y (F[406]), .A (nx5753), .E (nx6001)) ;
    inv01 ix5754 (.Y (nx5753), .A (D[406])) ;
    tri01 tri_F_407 (.Y (F[407]), .A (nx5756), .E (nx6001)) ;
    inv01 ix5757 (.Y (nx5756), .A (D[407])) ;
    tri01 tri_F_408 (.Y (F[408]), .A (nx5759), .E (nx6001)) ;
    inv01 ix5760 (.Y (nx5759), .A (D[408])) ;
    tri01 tri_F_409 (.Y (F[409]), .A (nx5762), .E (nx6001)) ;
    inv01 ix5763 (.Y (nx5762), .A (D[409])) ;
    tri01 tri_F_410 (.Y (F[410]), .A (nx5765), .E (nx6001)) ;
    inv01 ix5766 (.Y (nx5765), .A (D[410])) ;
    tri01 tri_F_411 (.Y (F[411]), .A (nx5768), .E (nx6001)) ;
    inv01 ix5769 (.Y (nx5768), .A (D[411])) ;
    tri01 tri_F_412 (.Y (F[412]), .A (nx5771), .E (nx6001)) ;
    inv01 ix5772 (.Y (nx5771), .A (D[412])) ;
    tri01 tri_F_413 (.Y (F[413]), .A (nx5774), .E (nx6003)) ;
    inv01 ix5775 (.Y (nx5774), .A (D[413])) ;
    tri01 tri_F_414 (.Y (F[414]), .A (nx5777), .E (nx6003)) ;
    inv01 ix5778 (.Y (nx5777), .A (D[414])) ;
    tri01 tri_F_415 (.Y (F[415]), .A (nx5780), .E (nx6003)) ;
    inv01 ix5781 (.Y (nx5780), .A (D[415])) ;
    tri01 tri_F_416 (.Y (F[416]), .A (nx5783), .E (nx6003)) ;
    inv01 ix5784 (.Y (nx5783), .A (D[416])) ;
    tri01 tri_F_417 (.Y (F[417]), .A (nx5786), .E (nx6003)) ;
    inv01 ix5787 (.Y (nx5786), .A (D[417])) ;
    tri01 tri_F_418 (.Y (F[418]), .A (nx5789), .E (nx6003)) ;
    inv01 ix5790 (.Y (nx5789), .A (D[418])) ;
    tri01 tri_F_419 (.Y (F[419]), .A (nx5792), .E (nx6003)) ;
    inv01 ix5793 (.Y (nx5792), .A (D[419])) ;
    tri01 tri_F_420 (.Y (F[420]), .A (nx5795), .E (nx6005)) ;
    inv01 ix5796 (.Y (nx5795), .A (D[420])) ;
    tri01 tri_F_421 (.Y (F[421]), .A (nx5798), .E (nx6005)) ;
    inv01 ix5799 (.Y (nx5798), .A (D[421])) ;
    tri01 tri_F_422 (.Y (F[422]), .A (nx5801), .E (nx6005)) ;
    inv01 ix5802 (.Y (nx5801), .A (D[422])) ;
    tri01 tri_F_423 (.Y (F[423]), .A (nx5804), .E (nx6005)) ;
    inv01 ix5805 (.Y (nx5804), .A (D[423])) ;
    tri01 tri_F_424 (.Y (F[424]), .A (nx5807), .E (nx6005)) ;
    inv01 ix5808 (.Y (nx5807), .A (D[424])) ;
    tri01 tri_F_425 (.Y (F[425]), .A (nx5810), .E (nx6005)) ;
    inv01 ix5811 (.Y (nx5810), .A (D[425])) ;
    tri01 tri_F_426 (.Y (F[426]), .A (nx5813), .E (nx6005)) ;
    inv01 ix5814 (.Y (nx5813), .A (D[426])) ;
    tri01 tri_F_427 (.Y (F[427]), .A (nx5816), .E (nx6007)) ;
    inv01 ix5817 (.Y (nx5816), .A (D[427])) ;
    tri01 tri_F_428 (.Y (F[428]), .A (nx5819), .E (nx6007)) ;
    inv01 ix5820 (.Y (nx5819), .A (D[428])) ;
    tri01 tri_F_429 (.Y (F[429]), .A (nx5822), .E (nx6007)) ;
    inv01 ix5823 (.Y (nx5822), .A (D[429])) ;
    tri01 tri_F_430 (.Y (F[430]), .A (nx5825), .E (nx6007)) ;
    inv01 ix5826 (.Y (nx5825), .A (D[430])) ;
    tri01 tri_F_431 (.Y (F[431]), .A (nx5828), .E (nx6007)) ;
    inv01 ix5829 (.Y (nx5828), .A (D[431])) ;
    tri01 tri_F_432 (.Y (F[432]), .A (nx5831), .E (nx6007)) ;
    inv01 ix5832 (.Y (nx5831), .A (D[432])) ;
    tri01 tri_F_433 (.Y (F[433]), .A (nx5834), .E (nx6007)) ;
    inv01 ix5835 (.Y (nx5834), .A (D[433])) ;
    tri01 tri_F_434 (.Y (F[434]), .A (nx5837), .E (nx6009)) ;
    inv01 ix5838 (.Y (nx5837), .A (D[434])) ;
    tri01 tri_F_435 (.Y (F[435]), .A (nx5840), .E (nx6009)) ;
    inv01 ix5841 (.Y (nx5840), .A (D[435])) ;
    tri01 tri_F_436 (.Y (F[436]), .A (nx5843), .E (nx6009)) ;
    inv01 ix5844 (.Y (nx5843), .A (D[436])) ;
    tri01 tri_F_437 (.Y (F[437]), .A (nx5846), .E (nx6009)) ;
    inv01 ix5847 (.Y (nx5846), .A (D[437])) ;
    tri01 tri_F_438 (.Y (F[438]), .A (nx5849), .E (nx6009)) ;
    inv01 ix5850 (.Y (nx5849), .A (D[438])) ;
    tri01 tri_F_439 (.Y (F[439]), .A (nx5852), .E (nx6009)) ;
    inv01 ix5853 (.Y (nx5852), .A (D[439])) ;
    tri01 tri_F_440 (.Y (F[440]), .A (nx5855), .E (nx6009)) ;
    inv01 ix5856 (.Y (nx5855), .A (D[440])) ;
    tri01 tri_F_441 (.Y (F[441]), .A (nx5858), .E (nx6011)) ;
    inv01 ix5859 (.Y (nx5858), .A (D[441])) ;
    tri01 tri_F_442 (.Y (F[442]), .A (nx5861), .E (nx6011)) ;
    inv01 ix5862 (.Y (nx5861), .A (D[442])) ;
    tri01 tri_F_443 (.Y (F[443]), .A (nx5864), .E (nx6011)) ;
    inv01 ix5865 (.Y (nx5864), .A (D[443])) ;
    tri01 tri_F_444 (.Y (F[444]), .A (nx5867), .E (nx6011)) ;
    inv01 ix5868 (.Y (nx5867), .A (D[444])) ;
    tri01 tri_F_445 (.Y (F[445]), .A (nx5870), .E (nx6011)) ;
    inv01 ix5871 (.Y (nx5870), .A (D[445])) ;
    tri01 tri_F_446 (.Y (F[446]), .A (nx5873), .E (nx6011)) ;
    inv01 ix5874 (.Y (nx5873), .A (D[446])) ;
    tri01 tri_F_447 (.Y (F[447]), .A (nx5876), .E (nx6011)) ;
    inv01 ix5877 (.Y (nx5876), .A (D[447])) ;
    inv01 ix5882 (.Y (nx5883), .A (EN)) ;
    inv01 ix5884 (.Y (nx5885), .A (nx6013)) ;
    inv01 ix5886 (.Y (nx5887), .A (nx6013)) ;
    inv01 ix5888 (.Y (nx5889), .A (nx6013)) ;
    inv01 ix5890 (.Y (nx5891), .A (nx6013)) ;
    inv01 ix5892 (.Y (nx5893), .A (nx6013)) ;
    inv01 ix5894 (.Y (nx5895), .A (nx6013)) ;
    inv01 ix5896 (.Y (nx5897), .A (nx6013)) ;
    inv01 ix5898 (.Y (nx5899), .A (nx6015)) ;
    inv01 ix5900 (.Y (nx5901), .A (nx6015)) ;
    inv01 ix5902 (.Y (nx5903), .A (nx6015)) ;
    inv01 ix5904 (.Y (nx5905), .A (nx6015)) ;
    inv01 ix5906 (.Y (nx5907), .A (nx6015)) ;
    inv01 ix5908 (.Y (nx5909), .A (nx6015)) ;
    inv01 ix5910 (.Y (nx5911), .A (nx6015)) ;
    inv01 ix5912 (.Y (nx5913), .A (nx6017)) ;
    inv01 ix5914 (.Y (nx5915), .A (nx6017)) ;
    inv01 ix5916 (.Y (nx5917), .A (nx6017)) ;
    inv01 ix5918 (.Y (nx5919), .A (nx6017)) ;
    inv01 ix5920 (.Y (nx5921), .A (nx6017)) ;
    inv01 ix5922 (.Y (nx5923), .A (nx6017)) ;
    inv01 ix5924 (.Y (nx5925), .A (nx6017)) ;
    inv01 ix5926 (.Y (nx5927), .A (nx6019)) ;
    inv01 ix5928 (.Y (nx5929), .A (nx6019)) ;
    inv01 ix5930 (.Y (nx5931), .A (nx6019)) ;
    inv01 ix5932 (.Y (nx5933), .A (nx6019)) ;
    inv01 ix5934 (.Y (nx5935), .A (nx6019)) ;
    inv01 ix5936 (.Y (nx5937), .A (nx6019)) ;
    inv01 ix5938 (.Y (nx5939), .A (nx6019)) ;
    inv01 ix5940 (.Y (nx5941), .A (nx6021)) ;
    inv01 ix5942 (.Y (nx5943), .A (nx6021)) ;
    inv01 ix5944 (.Y (nx5945), .A (nx6021)) ;
    inv01 ix5946 (.Y (nx5947), .A (nx6021)) ;
    inv01 ix5948 (.Y (nx5949), .A (nx6021)) ;
    inv01 ix5950 (.Y (nx5951), .A (nx6021)) ;
    inv01 ix5952 (.Y (nx5953), .A (nx6021)) ;
    inv01 ix5954 (.Y (nx5955), .A (nx6023)) ;
    inv01 ix5956 (.Y (nx5957), .A (nx6023)) ;
    inv01 ix5958 (.Y (nx5959), .A (nx6023)) ;
    inv01 ix5960 (.Y (nx5961), .A (nx6023)) ;
    inv01 ix5962 (.Y (nx5963), .A (nx6023)) ;
    inv01 ix5964 (.Y (nx5965), .A (nx6023)) ;
    inv01 ix5966 (.Y (nx5967), .A (nx6023)) ;
    inv01 ix5968 (.Y (nx5969), .A (nx6025)) ;
    inv01 ix5970 (.Y (nx5971), .A (nx6025)) ;
    inv01 ix5972 (.Y (nx5973), .A (nx6025)) ;
    inv01 ix5974 (.Y (nx5975), .A (nx6025)) ;
    inv01 ix5976 (.Y (nx5977), .A (nx6025)) ;
    inv01 ix5978 (.Y (nx5979), .A (nx6025)) ;
    inv01 ix5980 (.Y (nx5981), .A (nx6025)) ;
    inv01 ix5982 (.Y (nx5983), .A (nx6027)) ;
    inv01 ix5984 (.Y (nx5985), .A (nx6027)) ;
    inv01 ix5986 (.Y (nx5987), .A (nx6027)) ;
    inv01 ix5988 (.Y (nx5989), .A (nx6027)) ;
    inv01 ix5990 (.Y (nx5991), .A (nx6027)) ;
    inv01 ix5992 (.Y (nx5993), .A (nx6027)) ;
    inv01 ix5994 (.Y (nx5995), .A (nx6027)) ;
    inv01 ix5996 (.Y (nx5997), .A (nx6029)) ;
    inv01 ix5998 (.Y (nx5999), .A (nx6029)) ;
    inv01 ix6000 (.Y (nx6001), .A (nx6029)) ;
    inv01 ix6002 (.Y (nx6003), .A (nx6029)) ;
    inv01 ix6004 (.Y (nx6005), .A (nx6029)) ;
    inv01 ix6006 (.Y (nx6007), .A (nx6029)) ;
    inv01 ix6008 (.Y (nx6009), .A (nx6029)) ;
    inv01 ix6010 (.Y (nx6011), .A (nx5883)) ;
    inv01 ix6012 (.Y (nx6013), .A (nx6035)) ;
    inv01 ix6014 (.Y (nx6015), .A (nx6035)) ;
    inv01 ix6016 (.Y (nx6017), .A (nx6035)) ;
    inv01 ix6018 (.Y (nx6019), .A (nx6035)) ;
    inv01 ix6020 (.Y (nx6021), .A (nx6035)) ;
    inv01 ix6022 (.Y (nx6023), .A (nx6035)) ;
    inv01 ix6024 (.Y (nx6025), .A (nx6035)) ;
    inv01 ix6026 (.Y (nx6027), .A (nx6037)) ;
    inv01 ix6028 (.Y (nx6029), .A (nx6037)) ;
    inv01 ix6034 (.Y (nx6035), .A (nx5883)) ;
    inv01 ix6036 (.Y (nx6037), .A (nx5883)) ;
endmodule


module RAM_25 ( reset, CLK, W, R, address, dataIn, dataOut, MFC, counterOut ) ;

    input reset ;
    input CLK ;
    input W ;
    input R ;
    input [12:0]address ;
    input [15:0]dataIn ;
    output [399:0]dataOut ;
    output MFC ;
    output [3:0]counterOut ;

    wire nx12, nx30, nx34, nx42, nx46, nx52, nx98, nx104, nx114, nx116, nx118, 
         nx6151, nx6153, nx6156, nx6161, nx6168, nx6175, nx6177, nx6179, nx6181, 
         nx6183, nx6194, nx1, nx5;



    assign dataOut[399] = dataOut[0] ;
    assign dataOut[398] = dataOut[0] ;
    assign dataOut[397] = dataOut[0] ;
    assign dataOut[396] = dataOut[0] ;
    assign dataOut[395] = dataOut[0] ;
    assign dataOut[394] = dataOut[0] ;
    assign dataOut[393] = dataOut[0] ;
    assign dataOut[392] = dataOut[0] ;
    assign dataOut[391] = dataOut[0] ;
    assign dataOut[390] = dataOut[0] ;
    assign dataOut[389] = dataOut[0] ;
    assign dataOut[388] = dataOut[0] ;
    assign dataOut[387] = dataOut[0] ;
    assign dataOut[386] = dataOut[0] ;
    assign dataOut[385] = dataOut[0] ;
    assign dataOut[384] = dataOut[0] ;
    assign dataOut[383] = dataOut[0] ;
    assign dataOut[382] = dataOut[0] ;
    assign dataOut[381] = dataOut[0] ;
    assign dataOut[380] = dataOut[0] ;
    assign dataOut[379] = dataOut[0] ;
    assign dataOut[378] = dataOut[0] ;
    assign dataOut[377] = dataOut[0] ;
    assign dataOut[376] = dataOut[0] ;
    assign dataOut[375] = dataOut[0] ;
    assign dataOut[374] = dataOut[0] ;
    assign dataOut[373] = dataOut[0] ;
    assign dataOut[372] = dataOut[0] ;
    assign dataOut[371] = dataOut[0] ;
    assign dataOut[370] = dataOut[0] ;
    assign dataOut[369] = dataOut[0] ;
    assign dataOut[368] = dataOut[0] ;
    assign dataOut[367] = dataOut[0] ;
    assign dataOut[366] = dataOut[0] ;
    assign dataOut[365] = dataOut[0] ;
    assign dataOut[364] = dataOut[0] ;
    assign dataOut[363] = dataOut[0] ;
    assign dataOut[362] = dataOut[0] ;
    assign dataOut[361] = dataOut[0] ;
    assign dataOut[360] = dataOut[0] ;
    assign dataOut[359] = dataOut[0] ;
    assign dataOut[358] = dataOut[0] ;
    assign dataOut[357] = dataOut[0] ;
    assign dataOut[356] = dataOut[0] ;
    assign dataOut[355] = dataOut[0] ;
    assign dataOut[354] = dataOut[0] ;
    assign dataOut[353] = dataOut[0] ;
    assign dataOut[352] = dataOut[0] ;
    assign dataOut[351] = dataOut[0] ;
    assign dataOut[350] = dataOut[0] ;
    assign dataOut[349] = dataOut[0] ;
    assign dataOut[348] = dataOut[0] ;
    assign dataOut[347] = dataOut[0] ;
    assign dataOut[346] = dataOut[0] ;
    assign dataOut[345] = dataOut[0] ;
    assign dataOut[344] = dataOut[0] ;
    assign dataOut[343] = dataOut[0] ;
    assign dataOut[342] = dataOut[0] ;
    assign dataOut[341] = dataOut[0] ;
    assign dataOut[340] = dataOut[0] ;
    assign dataOut[339] = dataOut[0] ;
    assign dataOut[338] = dataOut[0] ;
    assign dataOut[337] = dataOut[0] ;
    assign dataOut[336] = dataOut[0] ;
    assign dataOut[335] = dataOut[0] ;
    assign dataOut[334] = dataOut[0] ;
    assign dataOut[333] = dataOut[0] ;
    assign dataOut[332] = dataOut[0] ;
    assign dataOut[331] = dataOut[0] ;
    assign dataOut[330] = dataOut[0] ;
    assign dataOut[329] = dataOut[0] ;
    assign dataOut[328] = dataOut[0] ;
    assign dataOut[327] = dataOut[0] ;
    assign dataOut[326] = dataOut[0] ;
    assign dataOut[325] = dataOut[0] ;
    assign dataOut[324] = dataOut[0] ;
    assign dataOut[323] = dataOut[0] ;
    assign dataOut[322] = dataOut[0] ;
    assign dataOut[321] = dataOut[0] ;
    assign dataOut[320] = dataOut[0] ;
    assign dataOut[319] = dataOut[0] ;
    assign dataOut[318] = dataOut[0] ;
    assign dataOut[317] = dataOut[0] ;
    assign dataOut[316] = dataOut[0] ;
    assign dataOut[315] = dataOut[0] ;
    assign dataOut[314] = dataOut[0] ;
    assign dataOut[313] = dataOut[0] ;
    assign dataOut[312] = dataOut[0] ;
    assign dataOut[311] = dataOut[0] ;
    assign dataOut[310] = dataOut[0] ;
    assign dataOut[309] = dataOut[0] ;
    assign dataOut[308] = dataOut[0] ;
    assign dataOut[307] = dataOut[0] ;
    assign dataOut[306] = dataOut[0] ;
    assign dataOut[305] = dataOut[0] ;
    assign dataOut[304] = dataOut[0] ;
    assign dataOut[303] = dataOut[0] ;
    assign dataOut[302] = dataOut[0] ;
    assign dataOut[301] = dataOut[0] ;
    assign dataOut[300] = dataOut[0] ;
    assign dataOut[299] = dataOut[0] ;
    assign dataOut[298] = dataOut[0] ;
    assign dataOut[297] = dataOut[0] ;
    assign dataOut[296] = dataOut[0] ;
    assign dataOut[295] = dataOut[0] ;
    assign dataOut[294] = dataOut[0] ;
    assign dataOut[293] = dataOut[0] ;
    assign dataOut[292] = dataOut[0] ;
    assign dataOut[291] = dataOut[0] ;
    assign dataOut[290] = dataOut[0] ;
    assign dataOut[289] = dataOut[0] ;
    assign dataOut[288] = dataOut[0] ;
    assign dataOut[287] = dataOut[0] ;
    assign dataOut[286] = dataOut[0] ;
    assign dataOut[285] = dataOut[0] ;
    assign dataOut[284] = dataOut[0] ;
    assign dataOut[283] = dataOut[0] ;
    assign dataOut[282] = dataOut[0] ;
    assign dataOut[281] = dataOut[0] ;
    assign dataOut[280] = dataOut[0] ;
    assign dataOut[279] = dataOut[0] ;
    assign dataOut[278] = dataOut[0] ;
    assign dataOut[277] = dataOut[0] ;
    assign dataOut[276] = dataOut[0] ;
    assign dataOut[275] = dataOut[0] ;
    assign dataOut[274] = dataOut[0] ;
    assign dataOut[273] = dataOut[0] ;
    assign dataOut[272] = dataOut[0] ;
    assign dataOut[271] = dataOut[0] ;
    assign dataOut[270] = dataOut[0] ;
    assign dataOut[269] = dataOut[0] ;
    assign dataOut[268] = dataOut[0] ;
    assign dataOut[267] = dataOut[0] ;
    assign dataOut[266] = dataOut[0] ;
    assign dataOut[265] = dataOut[0] ;
    assign dataOut[264] = dataOut[0] ;
    assign dataOut[263] = dataOut[0] ;
    assign dataOut[262] = dataOut[0] ;
    assign dataOut[261] = dataOut[0] ;
    assign dataOut[260] = dataOut[0] ;
    assign dataOut[259] = dataOut[0] ;
    assign dataOut[258] = dataOut[0] ;
    assign dataOut[257] = dataOut[0] ;
    assign dataOut[256] = dataOut[0] ;
    assign dataOut[255] = dataOut[0] ;
    assign dataOut[254] = dataOut[0] ;
    assign dataOut[253] = dataOut[0] ;
    assign dataOut[252] = dataOut[0] ;
    assign dataOut[251] = dataOut[0] ;
    assign dataOut[250] = dataOut[0] ;
    assign dataOut[249] = dataOut[0] ;
    assign dataOut[248] = dataOut[0] ;
    assign dataOut[247] = dataOut[0] ;
    assign dataOut[246] = dataOut[0] ;
    assign dataOut[245] = dataOut[0] ;
    assign dataOut[244] = dataOut[0] ;
    assign dataOut[243] = dataOut[0] ;
    assign dataOut[242] = dataOut[0] ;
    assign dataOut[241] = dataOut[0] ;
    assign dataOut[240] = dataOut[0] ;
    assign dataOut[239] = dataOut[0] ;
    assign dataOut[238] = dataOut[0] ;
    assign dataOut[237] = dataOut[0] ;
    assign dataOut[236] = dataOut[0] ;
    assign dataOut[235] = dataOut[0] ;
    assign dataOut[234] = dataOut[0] ;
    assign dataOut[233] = dataOut[0] ;
    assign dataOut[232] = dataOut[0] ;
    assign dataOut[231] = dataOut[0] ;
    assign dataOut[230] = dataOut[0] ;
    assign dataOut[229] = dataOut[0] ;
    assign dataOut[228] = dataOut[0] ;
    assign dataOut[227] = dataOut[0] ;
    assign dataOut[226] = dataOut[0] ;
    assign dataOut[225] = dataOut[0] ;
    assign dataOut[224] = dataOut[0] ;
    assign dataOut[223] = dataOut[0] ;
    assign dataOut[222] = dataOut[0] ;
    assign dataOut[221] = dataOut[0] ;
    assign dataOut[220] = dataOut[0] ;
    assign dataOut[219] = dataOut[0] ;
    assign dataOut[218] = dataOut[0] ;
    assign dataOut[217] = dataOut[0] ;
    assign dataOut[216] = dataOut[0] ;
    assign dataOut[215] = dataOut[0] ;
    assign dataOut[214] = dataOut[0] ;
    assign dataOut[213] = dataOut[0] ;
    assign dataOut[212] = dataOut[0] ;
    assign dataOut[211] = dataOut[0] ;
    assign dataOut[210] = dataOut[0] ;
    assign dataOut[209] = dataOut[0] ;
    assign dataOut[208] = dataOut[0] ;
    assign dataOut[207] = dataOut[0] ;
    assign dataOut[206] = dataOut[0] ;
    assign dataOut[205] = dataOut[0] ;
    assign dataOut[204] = dataOut[0] ;
    assign dataOut[203] = dataOut[0] ;
    assign dataOut[202] = dataOut[0] ;
    assign dataOut[201] = dataOut[0] ;
    assign dataOut[200] = dataOut[0] ;
    assign dataOut[199] = dataOut[0] ;
    assign dataOut[198] = dataOut[0] ;
    assign dataOut[197] = dataOut[0] ;
    assign dataOut[196] = dataOut[0] ;
    assign dataOut[195] = dataOut[0] ;
    assign dataOut[194] = dataOut[0] ;
    assign dataOut[193] = dataOut[0] ;
    assign dataOut[192] = dataOut[0] ;
    assign dataOut[191] = dataOut[0] ;
    assign dataOut[190] = dataOut[0] ;
    assign dataOut[189] = dataOut[0] ;
    assign dataOut[188] = dataOut[0] ;
    assign dataOut[187] = dataOut[0] ;
    assign dataOut[186] = dataOut[0] ;
    assign dataOut[185] = dataOut[0] ;
    assign dataOut[184] = dataOut[0] ;
    assign dataOut[183] = dataOut[0] ;
    assign dataOut[182] = dataOut[0] ;
    assign dataOut[181] = dataOut[0] ;
    assign dataOut[180] = dataOut[0] ;
    assign dataOut[179] = dataOut[0] ;
    assign dataOut[178] = dataOut[0] ;
    assign dataOut[177] = dataOut[0] ;
    assign dataOut[176] = dataOut[0] ;
    assign dataOut[175] = dataOut[0] ;
    assign dataOut[174] = dataOut[0] ;
    assign dataOut[173] = dataOut[0] ;
    assign dataOut[172] = dataOut[0] ;
    assign dataOut[171] = dataOut[0] ;
    assign dataOut[170] = dataOut[0] ;
    assign dataOut[169] = dataOut[0] ;
    assign dataOut[168] = dataOut[0] ;
    assign dataOut[167] = dataOut[0] ;
    assign dataOut[166] = dataOut[0] ;
    assign dataOut[165] = dataOut[0] ;
    assign dataOut[164] = dataOut[0] ;
    assign dataOut[163] = dataOut[0] ;
    assign dataOut[162] = dataOut[0] ;
    assign dataOut[161] = dataOut[0] ;
    assign dataOut[160] = dataOut[0] ;
    assign dataOut[159] = dataOut[0] ;
    assign dataOut[158] = dataOut[0] ;
    assign dataOut[157] = dataOut[0] ;
    assign dataOut[156] = dataOut[0] ;
    assign dataOut[155] = dataOut[0] ;
    assign dataOut[154] = dataOut[0] ;
    assign dataOut[153] = dataOut[0] ;
    assign dataOut[152] = dataOut[0] ;
    assign dataOut[151] = dataOut[0] ;
    assign dataOut[150] = dataOut[0] ;
    assign dataOut[149] = dataOut[0] ;
    assign dataOut[148] = dataOut[0] ;
    assign dataOut[147] = dataOut[0] ;
    assign dataOut[146] = dataOut[0] ;
    assign dataOut[145] = dataOut[0] ;
    assign dataOut[144] = dataOut[0] ;
    assign dataOut[143] = dataOut[0] ;
    assign dataOut[142] = dataOut[0] ;
    assign dataOut[141] = dataOut[0] ;
    assign dataOut[140] = dataOut[0] ;
    assign dataOut[139] = dataOut[0] ;
    assign dataOut[138] = dataOut[0] ;
    assign dataOut[137] = dataOut[0] ;
    assign dataOut[136] = dataOut[0] ;
    assign dataOut[135] = dataOut[0] ;
    assign dataOut[134] = dataOut[0] ;
    assign dataOut[133] = dataOut[0] ;
    assign dataOut[132] = dataOut[0] ;
    assign dataOut[131] = dataOut[0] ;
    assign dataOut[130] = dataOut[0] ;
    assign dataOut[129] = dataOut[0] ;
    assign dataOut[128] = dataOut[0] ;
    assign dataOut[127] = dataOut[0] ;
    assign dataOut[126] = dataOut[0] ;
    assign dataOut[125] = dataOut[0] ;
    assign dataOut[124] = dataOut[0] ;
    assign dataOut[123] = dataOut[0] ;
    assign dataOut[122] = dataOut[0] ;
    assign dataOut[121] = dataOut[0] ;
    assign dataOut[120] = dataOut[0] ;
    assign dataOut[119] = dataOut[0] ;
    assign dataOut[118] = dataOut[0] ;
    assign dataOut[117] = dataOut[0] ;
    assign dataOut[116] = dataOut[0] ;
    assign dataOut[115] = dataOut[0] ;
    assign dataOut[114] = dataOut[0] ;
    assign dataOut[113] = dataOut[0] ;
    assign dataOut[112] = dataOut[0] ;
    assign dataOut[111] = dataOut[0] ;
    assign dataOut[110] = dataOut[0] ;
    assign dataOut[109] = dataOut[0] ;
    assign dataOut[108] = dataOut[0] ;
    assign dataOut[107] = dataOut[0] ;
    assign dataOut[106] = dataOut[0] ;
    assign dataOut[105] = dataOut[0] ;
    assign dataOut[104] = dataOut[0] ;
    assign dataOut[103] = dataOut[0] ;
    assign dataOut[102] = dataOut[0] ;
    assign dataOut[101] = dataOut[0] ;
    assign dataOut[100] = dataOut[0] ;
    assign dataOut[99] = dataOut[0] ;
    assign dataOut[98] = dataOut[0] ;
    assign dataOut[97] = dataOut[0] ;
    assign dataOut[96] = dataOut[0] ;
    assign dataOut[95] = dataOut[0] ;
    assign dataOut[94] = dataOut[0] ;
    assign dataOut[93] = dataOut[0] ;
    assign dataOut[92] = dataOut[0] ;
    assign dataOut[91] = dataOut[0] ;
    assign dataOut[90] = dataOut[0] ;
    assign dataOut[89] = dataOut[0] ;
    assign dataOut[88] = dataOut[0] ;
    assign dataOut[87] = dataOut[0] ;
    assign dataOut[86] = dataOut[0] ;
    assign dataOut[85] = dataOut[0] ;
    assign dataOut[84] = dataOut[0] ;
    assign dataOut[83] = dataOut[0] ;
    assign dataOut[82] = dataOut[0] ;
    assign dataOut[81] = dataOut[0] ;
    assign dataOut[80] = dataOut[0] ;
    assign dataOut[79] = dataOut[0] ;
    assign dataOut[78] = dataOut[0] ;
    assign dataOut[77] = dataOut[0] ;
    assign dataOut[76] = dataOut[0] ;
    assign dataOut[75] = dataOut[0] ;
    assign dataOut[74] = dataOut[0] ;
    assign dataOut[73] = dataOut[0] ;
    assign dataOut[72] = dataOut[0] ;
    assign dataOut[71] = dataOut[0] ;
    assign dataOut[70] = dataOut[0] ;
    assign dataOut[69] = dataOut[0] ;
    assign dataOut[68] = dataOut[0] ;
    assign dataOut[67] = dataOut[0] ;
    assign dataOut[66] = dataOut[0] ;
    assign dataOut[65] = dataOut[0] ;
    assign dataOut[64] = dataOut[0] ;
    assign dataOut[63] = dataOut[0] ;
    assign dataOut[62] = dataOut[0] ;
    assign dataOut[61] = dataOut[0] ;
    assign dataOut[60] = dataOut[0] ;
    assign dataOut[59] = dataOut[0] ;
    assign dataOut[58] = dataOut[0] ;
    assign dataOut[57] = dataOut[0] ;
    assign dataOut[56] = dataOut[0] ;
    assign dataOut[55] = dataOut[0] ;
    assign dataOut[54] = dataOut[0] ;
    assign dataOut[53] = dataOut[0] ;
    assign dataOut[52] = dataOut[0] ;
    assign dataOut[51] = dataOut[0] ;
    assign dataOut[50] = dataOut[0] ;
    assign dataOut[49] = dataOut[0] ;
    assign dataOut[48] = dataOut[0] ;
    assign dataOut[47] = dataOut[0] ;
    assign dataOut[46] = dataOut[0] ;
    assign dataOut[45] = dataOut[0] ;
    assign dataOut[44] = dataOut[0] ;
    assign dataOut[43] = dataOut[0] ;
    assign dataOut[42] = dataOut[0] ;
    assign dataOut[41] = dataOut[0] ;
    assign dataOut[40] = dataOut[0] ;
    assign dataOut[39] = dataOut[0] ;
    assign dataOut[38] = dataOut[0] ;
    assign dataOut[37] = dataOut[0] ;
    assign dataOut[36] = dataOut[0] ;
    assign dataOut[35] = dataOut[0] ;
    assign dataOut[34] = dataOut[0] ;
    assign dataOut[33] = dataOut[0] ;
    assign dataOut[32] = dataOut[0] ;
    assign dataOut[31] = dataOut[0] ;
    assign dataOut[30] = dataOut[0] ;
    assign dataOut[29] = dataOut[0] ;
    assign dataOut[28] = dataOut[0] ;
    assign dataOut[27] = dataOut[0] ;
    assign dataOut[26] = dataOut[0] ;
    assign dataOut[25] = dataOut[0] ;
    assign dataOut[24] = dataOut[0] ;
    assign dataOut[23] = dataOut[0] ;
    assign dataOut[22] = dataOut[0] ;
    assign dataOut[21] = dataOut[0] ;
    assign dataOut[20] = dataOut[0] ;
    assign dataOut[19] = dataOut[0] ;
    assign dataOut[18] = dataOut[0] ;
    assign dataOut[17] = dataOut[0] ;
    assign dataOut[16] = dataOut[0] ;
    assign dataOut[15] = dataOut[0] ;
    assign dataOut[14] = dataOut[0] ;
    assign dataOut[13] = dataOut[0] ;
    assign dataOut[12] = dataOut[0] ;
    assign dataOut[11] = dataOut[0] ;
    assign dataOut[10] = dataOut[0] ;
    assign dataOut[9] = dataOut[0] ;
    assign dataOut[8] = dataOut[0] ;
    assign dataOut[7] = dataOut[0] ;
    assign dataOut[6] = dataOut[0] ;
    assign dataOut[5] = dataOut[0] ;
    assign dataOut[4] = dataOut[0] ;
    assign dataOut[3] = dataOut[0] ;
    assign dataOut[2] = dataOut[0] ;
    assign dataOut[1] = dataOut[0] ;
    fake_vcc ix117 (.Y (nx116)) ;
    ao21 ix61 (.Y (counterOut[1]), .A0 (dataIn[1]), .A1 (nx52), .B0 (nx46)) ;
    nor02_2x ix53 (.Y (nx52), .A0 (nx42), .A1 (nx46)) ;
    nor03_2x ix43 (.Y (nx42), .A0 (nx6151), .A1 (nx6153), .A2 (nx6156)) ;
    nand04 ix6152 (.Y (nx6151), .A0 (address[1]), .A1 (address[2]), .A2 (
           address[3]), .A3 (address[4])) ;
    nand03 ix6154 (.Y (nx6153), .A0 (address[5]), .A1 (address[6]), .A2 (nx12)
           ) ;
    nor02_2x ix13 (.Y (nx12), .A0 (address[12]), .A1 (address[11])) ;
    nand04 ix6157 (.Y (nx6156), .A0 (nx30), .A1 (nx34), .A2 (reset), .A3 (CLK)
           ) ;
    nor04 ix31 (.Y (nx30), .A0 (address[10]), .A1 (address[9]), .A2 (address[8])
          , .A3 (address[7])) ;
    nor02ii ix35 (.Y (nx34), .A0 (address[0]), .A1 (W)) ;
    inv01 ix6162 (.Y (nx6161), .A (R)) ;
    ao21 ix65 (.Y (counterOut[2]), .A0 (dataIn[2]), .A1 (nx52), .B0 (nx46)) ;
    ao21 ix57 (.Y (counterOut[0]), .A0 (dataIn[0]), .A1 (nx6168), .B0 (nx42)) ;
    and02 ix67 (.Y (counterOut[3]), .A0 (dataIn[3]), .A1 (nx52)) ;
    nor04 ix115 (.Y (nx114), .A0 (nx6175), .A1 (nx6177), .A2 (nx6179), .A3 (
          nx6183)) ;
    nand03 ix6176 (.Y (nx6175), .A0 (dataIn[7]), .A1 (dataIn[4]), .A2 (dataIn[5]
           )) ;
    nand02 ix6178 (.Y (nx6177), .A0 (dataIn[9]), .A1 (dataIn[12])) ;
    nand04 ix6180 (.Y (nx6179), .A0 (dataIn[0]), .A1 (dataIn[1]), .A2 (dataIn[2]
           ), .A3 (nx6181)) ;
    inv01 ix6182 (.Y (nx6181), .A (dataIn[15])) ;
    nand04 ix6184 (.Y (nx6183), .A0 (nx98), .A1 (nx104), .A2 (dataIn[3]), .A3 (
           nx6161)) ;
    nor04 ix99 (.Y (nx98), .A0 (dataIn[14]), .A1 (dataIn[13]), .A2 (dataIn[11])
          , .A3 (dataIn[10])) ;
    nor02_2x ix105 (.Y (nx104), .A0 (dataIn[8]), .A1 (dataIn[6])) ;
    and02 ix119 (.Y (nx118), .A0 (R), .A1 (CLK)) ;
    inv01 ix6169 (.Y (nx6168), .A (nx46)) ;
    nor02ii ix47 (.Y (nx46), .A0 (CLK), .A1 (R)) ;
    and03 ix129 (.Y (MFC), .A0 (reset), .A1 (R), .A2 (nx6194)) ;
    inv01 ix6193 (.Y (nx6194), .A (W)) ;
    latchr lat_dataOut_0__u1 (.QB (nx5), .D (nx116), .CLK (nx114), .R (nx118)) ;
    inv01 lat_dataOut_0__u2 (.Y (dataOut[0]), .A (nx5)) ;
    buf02 lat_dataOut_0__u3 (.Y (nx1), .A (nx5)) ;
endmodule


module nBitRegister_13 ( D, CLK, RST, EN, Q ) ;

    input [12:0]D ;
    input CLK ;
    input RST ;
    input EN ;
    output [12:0]Q ;

    wire nx194, nx204, nx214, nx224, nx234, nx244, nx254, nx264, nx274, nx284, 
         nx294, nx304, nx314, nx370, nx372, nx378, nx380, nx382, nx384;
    wire [12:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx194), .CLK (nx370), .R (
         nx378)) ;
    mux21_ni ix195 (.Y (nx194), .A0 (Q[0]), .A1 (D[0]), .S0 (nx382)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx204), .CLK (nx370), .R (
         nx378)) ;
    mux21_ni ix205 (.Y (nx204), .A0 (Q[1]), .A1 (D[1]), .S0 (nx382)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx214), .CLK (nx370), .R (
         nx378)) ;
    mux21_ni ix215 (.Y (nx214), .A0 (Q[2]), .A1 (D[2]), .S0 (nx382)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx224), .CLK (nx370), .R (
         nx378)) ;
    mux21_ni ix225 (.Y (nx224), .A0 (Q[3]), .A1 (D[3]), .S0 (nx382)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx234), .CLK (nx370), .R (
         nx378)) ;
    mux21_ni ix235 (.Y (nx234), .A0 (Q[4]), .A1 (D[4]), .S0 (nx382)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx244), .CLK (nx370), .R (
         nx378)) ;
    mux21_ni ix245 (.Y (nx244), .A0 (Q[5]), .A1 (D[5]), .S0 (nx382)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx254), .CLK (nx370), .R (
         nx378)) ;
    mux21_ni ix255 (.Y (nx254), .A0 (Q[6]), .A1 (D[6]), .S0 (nx382)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx264), .CLK (nx372), .R (
         nx380)) ;
    mux21_ni ix265 (.Y (nx264), .A0 (Q[7]), .A1 (D[7]), .S0 (nx384)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx274), .CLK (nx372), .R (
         nx380)) ;
    mux21_ni ix275 (.Y (nx274), .A0 (Q[8]), .A1 (D[8]), .S0 (nx384)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx284), .CLK (nx372), .R (
         nx380)) ;
    mux21_ni ix285 (.Y (nx284), .A0 (Q[9]), .A1 (D[9]), .S0 (nx384)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx294), .CLK (nx372), .R (
         nx380)) ;
    mux21_ni ix295 (.Y (nx294), .A0 (Q[10]), .A1 (D[10]), .S0 (nx384)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx304), .CLK (nx372), .R (
         nx380)) ;
    mux21_ni ix305 (.Y (nx304), .A0 (Q[11]), .A1 (D[11]), .S0 (nx384)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx314), .CLK (nx372), .R (
         nx380)) ;
    mux21_ni ix315 (.Y (nx314), .A0 (Q[12]), .A1 (D[12]), .S0 (nx384)) ;
    inv02 ix369 (.Y (nx370), .A (CLK)) ;
    inv02 ix371 (.Y (nx372), .A (CLK)) ;
    buf02 ix377 (.Y (nx378), .A (RST)) ;
    buf02 ix379 (.Y (nx380), .A (RST)) ;
    buf02 ix381 (.Y (nx382), .A (EN)) ;
    buf02 ix383 (.Y (nx384), .A (EN)) ;
endmodule


module triStateBuffer_13 ( D, EN, F ) ;

    input [12:0]D ;
    input EN ;
    output [12:0]F ;

    wire nx185, nx188, nx191, nx194, nx197, nx200, nx203, nx206, nx209, nx212, 
         nx215, nx218, nx221, nx228, nx230;



    tri01 tri_F_0 (.Y (F[0]), .A (nx185), .E (nx228)) ;
    inv01 ix186 (.Y (nx185), .A (D[0])) ;
    tri01 tri_F_1 (.Y (F[1]), .A (nx188), .E (nx228)) ;
    inv01 ix189 (.Y (nx188), .A (D[1])) ;
    tri01 tri_F_2 (.Y (F[2]), .A (nx191), .E (nx228)) ;
    inv01 ix192 (.Y (nx191), .A (D[2])) ;
    tri01 tri_F_3 (.Y (F[3]), .A (nx194), .E (nx228)) ;
    inv01 ix195 (.Y (nx194), .A (D[3])) ;
    tri01 tri_F_4 (.Y (F[4]), .A (nx197), .E (nx228)) ;
    inv01 ix198 (.Y (nx197), .A (D[4])) ;
    tri01 tri_F_5 (.Y (F[5]), .A (nx200), .E (nx228)) ;
    inv01 ix201 (.Y (nx200), .A (D[5])) ;
    tri01 tri_F_6 (.Y (F[6]), .A (nx203), .E (nx228)) ;
    inv01 ix204 (.Y (nx203), .A (D[6])) ;
    tri01 tri_F_7 (.Y (F[7]), .A (nx206), .E (nx230)) ;
    inv01 ix207 (.Y (nx206), .A (D[7])) ;
    tri01 tri_F_8 (.Y (F[8]), .A (nx209), .E (nx230)) ;
    inv01 ix210 (.Y (nx209), .A (D[8])) ;
    tri01 tri_F_9 (.Y (F[9]), .A (nx212), .E (nx230)) ;
    inv01 ix213 (.Y (nx212), .A (D[9])) ;
    tri01 tri_F_10 (.Y (F[10]), .A (nx215), .E (nx230)) ;
    inv01 ix216 (.Y (nx215), .A (D[10])) ;
    tri01 tri_F_11 (.Y (F[11]), .A (nx218), .E (nx230)) ;
    inv01 ix219 (.Y (nx218), .A (D[11])) ;
    tri01 tri_F_12 (.Y (F[12]), .A (nx221), .E (nx230)) ;
    inv01 ix222 (.Y (nx221), .A (D[12])) ;
    buf02 ix227 (.Y (nx228), .A (EN)) ;
    buf02 ix229 (.Y (nx230), .A (EN)) ;
endmodule


module nBitRegister_1 ( D, CLK, RST, EN, Q ) ;

    input [0:0]D ;
    input CLK ;
    input RST ;
    input EN ;
    output [0:0]Q ;

    wire NOT_CLK, nx50;
    wire [0:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx50), .CLK (NOT_CLK), .R (
         RST)) ;
    mux21_ni ix51 (.Y (nx50), .A0 (Q[0]), .A1 (D[0]), .S0 (EN)) ;
    inv01 ix63 (.Y (NOT_CLK), .A (CLK)) ;
endmodule

