package constants is 

type state is (RI ,RL); 

end constants;